
module LZSS_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2XL U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVXL U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module LZSS ( clk, reset, data, data_valid, drop_done, busy, codeword, enc_num,
        out_valid, finish );
  input [31:0] data;
  output [10:0] codeword;
  output [11:0] enc_num;
  input clk, reset, data_valid, drop_done;
  output busy, out_valid, finish;
  wire   n51439, n51440, n51441, n51442, n51443, n51444, n51445, n51446,
         n51447, N23551, N23552, N23553, N23554, N23555, N23556, N23557,
         N23558, N23559, N23560, N23561, N23562, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9689, n9690, n9693, n9695, n9696,
         n9697, n9698, n9699, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9712, n9714, n9715, n9716, n9719, n9721, n9724, n9726, n9727, n9728,
         n9729, n9730, n9732, n9733, n9734, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9747, n9748, n9750, n9751, n9754, n9756, n9757,
         n9759, n9760, n9763, n9764, n9768, n9770, n9771, n9772, n9773, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9787, n9788, n9789,
         n9790, n9791, n9792, n9794, n9795, n9797, n9798, n9799, n9802, n9804,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9815, n9816,
         n9817, n9819, n9820, n9821, n9824, n9825, n9826, n9828, n9829, n9830,
         n9832, n9836, n9837, n9838, n9839, n9840, n9841, n9843, n9844, n9845,
         n9846, n9847, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9862, n9863, n9864, n9865, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9888, n9892, n9893, n9894, n9895, n9896, n9898, n9899,
         n9900, n9901, n9902, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9917, n9918, n9919, n9921, n9922, n9923, n9924,
         n9927, n9928, n9930, n9931, n9933, n9934, n9935, n9937, n9938, n9939,
         n9942, n9943, n9944, n9945, n9946, n9948, n9949, n9950, n9951, n9952,
         n9954, n9956, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9966,
         n9967, n9968, n9969, n9970, n9971, n9973, n9974, n9977, n9978, n9979,
         n9982, n9983, n9986, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9996, n9998, n9999, n10000, n10001, n10002, n10004, n10005, n10006,
         n10007, n10010, n10011, n10012, n10013, n10015, n10016, n10017,
         n10018, n10019, n10020, n10022, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10032, n10033, n10034, n10036, n10037,
         n10040, n10044, n10045, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10097,
         n10098, n10099, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10126, n10128, n10129, n10130, n10131, n10134, n10135, n10136,
         n10137, n10138, n10140, n10141, n10142, n10143, n10144, n10147,
         n10148, n10149, n10150, n10152, n10153, n10155, n10156, n10157,
         n10158, n10161, n10162, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10182, n10184, n10196, n10197, n10198, n10199,
         n10200, n10203, n10204, n10205, n10206, n10208, n10210, n10212,
         n10215, n10216, n10217, n10218, n10219, n10220, n10222, n10223,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10251, n10252, n10253, n10254, n10255, n10257, n10272, n10273,
         n10274, n10292, n10293, n10295, n10301, n10302, n10303, n10306,
         n10311, n10319, n10331, n10334, n10336, n10338, n10339, n10340,
         n10341, n10355, n10357, n10362, n10367, n10368, n10369, n10376,
         n10377, n10378, n10381, n10382, n10383, n10384, n10385, n10387,
         n10393, n10394, n10395, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10446, n10447,
         n10448, n10456, n10463, n10464, n10469, n10470, n10471, n10480,
         n10481, n10483, n10484, n10485, n10487, n10492, n10493, n10498,
         n10501, n10502, n10503, n10504, n10505, n10506, n10509, n10512,
         n10518, n10519, n10520, n10522, n10525, n10526, n10527, n10529,
         n10530, n10532, n10542, n10543, n10544, n10548, n10553, n10554,
         n10555, n10556, n10559, n10564, n10565, n10566, n10567, n10570,
         n10572, n10573, n10577, n10585, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10619, n10621, n10622,
         n10624, n10625, n10626, n10629, n10630, n10631, n10632, n10635,
         n10638, n10639, n10641, n10644, n10646, n10651, n10657, n10658,
         n10659, n10661, n10662, n10669, n10671, n10672, n10677, n10679,
         n10683, n10686, n10689, n10699, n10700, n10702, n10705, n10706,
         n10708, n10709, n10710, n10715, n10719, n10724, n10725, n10726,
         n10727, n10729, n10730, n10732, n10733, n10734, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10771, n10772, n10775, n10776, n10779,
         n10793, n10798, n10801, n10806, n10807, n10808, n10810, n10814,
         n10815, n10819, n10820, n10821, n10827, n10829, n10837, n10839,
         n10842, n10843, n10845, n10846, n10847, n10848, n10852, n10853,
         n10854, n10855, n10861, n10863, n10865, n10869, n10870, n10872,
         n10875, n10877, n10879, n10902, n10903, n10904, n10905, n10906,
         n10923, n10926, n10927, n10928, n10938, n10939, n10940, n10941,
         n10942, n10946, n10947, n10957, n10958, n10959, n10960, n10965,
         n10966, n10968, n10969, n10973, n10974, n10976, n10982, n10983,
         n10990, n10991, n10992, n10993, n10994, n10996, n10997, n10998,
         n11000, n11001, n11002, n11003, n11006, n11007, n11008, n11009,
         n11010, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11057, n11058,
         n11059, n11061, n11064, n11065, n11066, n11067, n11068, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11100,
         n11101, n11102, n11103, n11106, n11107, n11108, n11109, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11122,
         n11124, n11125, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11145, n11146, n11147, n11148, n11149, n11200, n11201, n11204,
         n11205, n11208, n11209, n11210, n11211, n11217, n11218, n11228,
         n11241, n11242, n11262, n11263, n11264, n11265, n11272, n11273,
         n11274, n11280, n11281, n11282, n11283, n11291, n11299, n11300,
         n11301, n11308, n11309, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11332, n11333, n11334, n11335, n11336,
         n11339, n11342, n11343, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11404, n11405, n11406, n11407, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11422, n11423, n11424, n11425, n11426, n11429, n11430,
         n11431, n11432, n11435, n11436, n11437, n11438, n11441, n11442,
         n11443, n11509, n11510, n11511, n11512, n11515, n11516, n11519,
         n11520, n11521, n11524, n11525, n11537, n11538, n11541, n11542,
         n11543, n11544, n11549, n11550, n11551, n11555, n11556, n11558,
         n11565, n11566, n11567, n11568, n11575, n11576, n11578, n11584,
         n11585, n11586, n11594, n11595, n11600, n11601, n11605, n11606,
         n11607, n11613, n11614, n11620, n11621, n11622, n11625, n11626,
         n11627, n11628, n11631, n11632, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11667, n11668, n11669,
         n11670, n11672, n11673, n11674, n11675, n11679, n11680, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11725, n11726, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11750, n11751, n11752, n11753,
         n11756, n11757, n11758, n11760, n11761, n11762, n11763, n11764,
         n11765, n11768, n11769, n11770, n11771, n11772, n11775, n11776,
         n11777, n11778, n11848, n11849, n11850, n11869, n11870, n11874,
         n11883, n11884, n11885, n11886, n11893, n11894, n11895, n11896,
         n11897, n11901, n11902, n11904, n11906, n11907, n11915, n11916,
         n11917, n11924, n11925, n11932, n11933, n11934, n11935, n11942,
         n11943, n11954, n11955, n11958, n11959, n11960, n11961, n11967,
         n11968, n11969, n11970, n11972, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11993, n11994, n11995, n11996,
         n11998, n11999, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12040, n12041, n12042, n12043, n12046, n12047, n12048,
         n12049, n12050, n12051, n12054, n12055, n12056, n12057, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12081, n12083, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12144, n12145, n12146, n12147, n12150, n12151,
         n12152, n12153, n12154, n12156, n12157, n12165, n12166, n12167,
         n12168, n12169, n12170, n12183, n12186, n12188, n12190, n12194,
         n12196, n12207, n12210, n12212, n12213, n12219, n12221, n12228,
         n12230, n12238, n12246, n12251, n12252, n12255, n12260, n12262,
         n12264, n12270, n12274, n12278, n12280, n12287, n12292, n12297,
         n12303, n12306, n12311, n12316, n12318, n12322, n12323, n12324,
         n12326, n12329, n12333, n12342, n12344, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12395, n12403,
         n12408, n12415, n12417, n12424, n12427, n12433, n12445, n12449,
         n12452, n12453, n12455, n12457, n12459, n12461, n12466, n12474,
         n12476, n12479, n12482, n12485, n12486, n12488, n12490, n12493,
         n12501, n12506, n12518, n12530, n12535, n12538, n12539, n12542,
         n12549, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12594, n12596, n12597, n12602,
         n12604, n12611, n12614, n12618, n12624, n12629, n12634, n12639,
         n12640, n12643, n12648, n12651, n12665, n12668, n12671, n12672,
         n12675, n12686, n12692, n12702, n12703, n12706, n12708, n12711,
         n12715, n12717, n12723, n12726, n12731, n12736, n12741, n12742,
         n12744, n12746, n12747, n12749, n12751, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12806, n12807, n12808, n12811, n12813, n12821, n12824,
         n12826, n12831, n12834, n12838, n12840, n12847, n12848, n12851,
         n12855, n12856, n12858, n12867, n12872, n12873, n12876, n12878,
         n12887, n12892, n12893, n12896, n12901, n12904, n12906, n12907,
         n12909, n12915, n12918, n12922, n12929, n12931, n12940, n12942,
         n12951, n12954, n12957, n12959, n12960, n12962, n12967, n12970,
         n12976, n13014, n13015, n13016, n13017, n13018, n13019, n13021,
         n13022, n13023, n13024, n13025, n13026, n13028, n13030, n13031,
         n13033, n13034, n13036, n13037, n13039, n13040, n13042, n13043,
         n13045, n13046, n13048, n13049, n13051, n13052, n13056, n13060,
         n13062, n13063, n13068, n13072, n13076, n13078, n13079, n13084,
         n13087, n13090, n13092, n13093, n13096, n13099, n13102, n13104,
         n13105, n13108, n13109, n13111, n13112, n13114, n13116, n13117,
         n13118, n13120, n13121, n13123, n13124, n13126, n13128, n13129,
         n13130, n13132, n13133, n13135, n13136, n13138, n13140, n13141,
         n13142, n13144, n13145, n13147, n13148, n13150, n13152, n13153,
         n13154, n13156, n13157, n13159, n13160, n13162, n13164, n13165,
         n13166, n13168, n13169, n13171, n13172, n13174, n13176, n13177,
         n13178, n13180, n13181, n13183, n13184, n13186, n13188, n13189,
         n13190, n13192, n13193, n13195, n13196, n13198, n13200, n13201,
         n13202, n13204, n13205, n13207, n13208, n13210, n13212, n13213,
         n13214, n13216, n13217, n13219, n13220, n13222, n13224, n13225,
         n13226, n13228, n13229, n13231, n13232, n13234, n13236, n13237,
         n13238, n13240, n13241, n13243, n13244, n13246, n13248, n13249,
         n13250, n13252, n13253, n13255, n13256, n13258, n13260, n13261,
         n13262, n13264, n13265, n13267, n13268, n13270, n13272, n13273,
         n13274, n13276, n13277, n13279, n13280, n13282, n13284, n13285,
         n13286, n13288, n13289, n13291, n13292, n13294, n13296, n13297,
         n13298, n13300, n13301, n13303, n13304, n13306, n13308, n13309,
         n13310, n13312, n13313, n13315, n13316, n13318, n13320, n13321,
         n13322, n13324, n13325, n13327, n13328, n13330, n13332, n13333,
         n13334, n13336, n13337, n13339, n13340, n13342, n13344, n13345,
         n13346, n13348, n13349, n13351, n13352, n13354, n13356, n13357,
         n13358, n13360, n13361, n13363, n13364, n13366, n13368, n13369,
         n13370, n13372, n13373, n13375, n13376, n13378, n13380, n13381,
         n13382, n13384, n13385, n13387, n13388, n13390, n13392, n13393,
         n13394, n13396, n13397, n13399, n13400, n13402, n13404, n13405,
         n13406, n13408, n13409, n13411, n13412, n13414, n13416, n13417,
         n13418, n13420, n13421, n13423, n13424, n13426, n13428, n13429,
         n13430, n13432, n13433, n13435, n13436, n13438, n13440, n13441,
         n13442, n13444, n13445, n13447, n13448, n13450, n13452, n13453,
         n13454, n13456, n13457, n13459, n13460, n13462, n13464, n13465,
         n13466, n13468, n13469, n13471, n13472, n13474, n13476, n13477,
         n13478, n13480, n13481, n13483, n13484, n13486, n13488, n13489,
         n13490, n13492, n13493, n13495, n13496, n13498, n13500, n13501,
         n13502, n13504, n13505, n13507, n13508, n13510, n13512, n13513,
         n13514, n13516, n13517, n13519, n13520, n13522, n13524, n13525,
         n13526, n13528, n13529, n13531, n13532, n13534, n13536, n13537,
         n13538, n13540, n13541, n13543, n13544, n13546, n13548, n13549,
         n13550, n13552, n13553, n13555, n13556, n13558, n13560, n13561,
         n13562, n13564, n13565, n13567, n13568, n13570, n13572, n13573,
         n13574, n13576, n13577, n13579, n13580, n13582, n13584, n13585,
         n13586, n13588, n13589, n13591, n13592, n13594, n13596, n13597,
         n13598, n13600, n13601, n13603, n13604, n13606, n13608, n13609,
         n13610, n13612, n13613, n13615, n13616, n13618, n13620, n13621,
         n13622, n13624, n13625, n13627, n13628, n13630, n13632, n13633,
         n13634, n13636, n13637, n13639, n13640, n13642, n13644, n13645,
         n13646, n13648, n13649, n13651, n13652, n13654, n13656, n13657,
         n13658, n13660, n13661, n13663, n13664, n13666, n13668, n13669,
         n13670, n13672, n13673, n13675, n13676, n13678, n13680, n13681,
         n13682, n13684, n13685, n13687, n13688, n13690, n13692, n13693,
         n13694, n13696, n13697, n13699, n13700, n13702, n13704, n13705,
         n13706, n13708, n13709, n13711, n13712, n13714, n13716, n13717,
         n13718, n13720, n13721, n13723, n13724, n13726, n13728, n13729,
         n13730, n13732, n13733, n13735, n13736, n13738, n13740, n13741,
         n13742, n13744, n13745, n13747, n13748, n13750, n13752, n13753,
         n13754, n13756, n13757, n13759, n13760, n13762, n13764, n13765,
         n13766, n13768, n13769, n13771, n13772, n13774, n13776, n13777,
         n13778, n13780, n13781, n13783, n13784, n13786, n13788, n13789,
         n13790, n13792, n13793, n13795, n13796, n13798, n13800, n13801,
         n13802, n13804, n13805, n13807, n13808, n13810, n13812, n13813,
         n13814, n13816, n13817, n13819, n13820, n13822, n13824, n13825,
         n13826, n13828, n13829, n13831, n13832, n13834, n13836, n13837,
         n13838, n13840, n13841, n13843, n13844, n13846, n13848, n13849,
         n13850, n13852, n13853, n13855, n13856, n13858, n13860, n13861,
         n13862, n13864, n13865, n13867, n13868, n13870, n13872, n13873,
         n13874, n13876, n13877, n13879, n13880, n13882, n13884, n13885,
         n13886, n13888, n13889, n13891, n13892, n13894, n13896, n13897,
         n13898, n13900, n13901, n13903, n13904, n13906, n13908, n13909,
         n13910, n13912, n13913, n13915, n13916, n13918, n13920, n13921,
         n13922, n13924, n13925, n13927, n13928, n13930, n13932, n13933,
         n13934, n13936, n13937, n13939, n13940, n13942, n13944, n13945,
         n13946, n13948, n13949, n13951, n13952, n13954, n13956, n13957,
         n13958, n13960, n13961, n13963, n13964, n13966, n13968, n13969,
         n13970, n13972, n13973, n13975, n13976, n13978, n13980, n13981,
         n13982, n13984, n13985, n13987, n13988, n13990, n13992, n13993,
         n13994, n13996, n13997, n13999, n14000, n14002, n14004, n14005,
         n14006, n14008, n14009, n14011, n14012, n14014, n14016, n14017,
         n14018, n14020, n14021, n14023, n14024, n14026, n14028, n14029,
         n14030, n14032, n14033, n14035, n14036, n14038, n14040, n14041,
         n14042, n14044, n14045, n14047, n14048, n14050, n14052, n14053,
         n14054, n14056, n14057, n14059, n14060, n14062, n14064, n14065,
         n14066, n14068, n14069, n14071, n14072, n14074, n14076, n14077,
         n14078, n14080, n14081, n14083, n14084, n14086, n14088, n14089,
         n14090, n14092, n14093, n14095, n14096, n14098, n14100, n14101,
         n14102, n14104, n14105, n14107, n14108, n14110, n14112, n14113,
         n14114, n14116, n14117, n14119, n14120, n14122, n14124, n14125,
         n14126, n14128, n14129, n14131, n14132, n14134, n14136, n14137,
         n14138, n14140, n14141, n14143, n14144, n14146, n14148, n14149,
         n14150, n14152, n14153, n14155, n14156, n14158, n14160, n14161,
         n14162, n14164, n14165, n14167, n14168, n14170, n14172, n14173,
         n14174, n14176, n14177, n14179, n14180, n14182, n14184, n14185,
         n14186, n14188, n14189, n14191, n14192, n14194, n14196, n14197,
         n14198, n14200, n14201, n14203, n14204, n14206, n14208, n14209,
         n14210, n14212, n14213, n14215, n14216, n14218, n14220, n14221,
         n14222, n14224, n14225, n14227, n14228, n14230, n14232, n14233,
         n14234, n14236, n14237, n14239, n14240, n14242, n14244, n14245,
         n14246, n14248, n14249, n14251, n14252, n14254, n14256, n14257,
         n14258, n14260, n14261, n14263, n14264, n14266, n14268, n14269,
         n14270, n14272, n14273, n14275, n14276, n14278, n14280, n14281,
         n14282, n14284, n14285, n14287, n14288, n14290, n14292, n14293,
         n14294, n14296, n14297, n14299, n14300, n14302, n14304, n14305,
         n14306, n14308, n14309, n14311, n14312, n14314, n14316, n14317,
         n14318, n14320, n14321, n14323, n14324, n14326, n14328, n14329,
         n14330, n14332, n14333, n14335, n14336, n14338, n14340, n14341,
         n14342, n14344, n14345, n14347, n14348, n14350, n14352, n14353,
         n14354, n14356, n14357, n14359, n14360, n14362, n14364, n14365,
         n14366, n14368, n14369, n14371, n14372, n14374, n14376, n14377,
         n14378, n14380, n14381, n14383, n14384, n14386, n14388, n14389,
         n14390, n14392, n14393, n14395, n14396, n14398, n14400, n14401,
         n14402, n14404, n14405, n14407, n14408, n14410, n14412, n14413,
         n14414, n14416, n14417, n14419, n14420, n14422, n14424, n14425,
         n14426, n14428, n14429, n14431, n14432, n14434, n14436, n14437,
         n14438, n14440, n14441, n14443, n14444, n14446, n14448, n14449,
         n14450, n14452, n14453, n14455, n14456, n14458, n14460, n14461,
         n14462, n14464, n14465, n14467, n14468, n14470, n14472, n14473,
         n14474, n14476, n14477, n14479, n14480, n14482, n14484, n14485,
         n14486, n14488, n14489, n14491, n14492, n14494, n14496, n14497,
         n14498, n14500, n14501, n14503, n14504, n14506, n14508, n14509,
         n14510, n14512, n14513, n14515, n14516, n14518, n14520, n14521,
         n14522, n14524, n14525, n14527, n14528, n14530, n14532, n14533,
         n14534, n14536, n14537, n14539, n14540, n14542, n14544, n14545,
         n14546, n14548, n14549, n14551, n14552, n14554, n14556, n14557,
         n14558, n14560, n14561, n14563, n14564, n14566, n14568, n14569,
         n14570, n14572, n14573, n14575, n14576, n14578, n14580, n14581,
         n14582, n14584, n14585, n14587, n14588, n14590, n14592, n14593,
         n14594, n14596, n14597, n14599, n14600, n14602, n14604, n14605,
         n14606, n14608, n14609, n14611, n14612, n14614, n14616, n14617,
         n14618, n14620, n14621, n14623, n14624, n14626, n14628, n14629,
         n14630, n14632, n14633, n14635, n14636, n14638, n14640, n14641,
         n14642, n14644, n14645, n14647, n14648, n14650, n14652, n14653,
         n14654, n14656, n14657, n14659, n14660, n14662, n14664, n14665,
         n14666, n14668, n14669, n14671, n14672, n14674, n14676, n14677,
         n14678, n14680, n14681, n14683, n14684, n14686, n14688, n14689,
         n14690, n14692, n14693, n14695, n14696, n14698, n14700, n14701,
         n14702, n14704, n14705, n14707, n14708, n14710, n14712, n14713,
         n14714, n14716, n14717, n14719, n14720, n14722, n14724, n14725,
         n14726, n14728, n14729, n14731, n14732, n14734, n14736, n14737,
         n14738, n14740, n14741, n14743, n14744, n14746, n14748, n14749,
         n14750, n14752, n14753, n14755, n14756, n14758, n14760, n14761,
         n14762, n14764, n14765, n14767, n14768, n14770, n14772, n14773,
         n14774, n14776, n14777, n14779, n14780, n14782, n14784, n14785,
         n14786, n14788, n14789, n14791, n14792, n14794, n14796, n14797,
         n14798, n14800, n14801, n14803, n14804, n14806, n14808, n14809,
         n14810, n14812, n14813, n14815, n14816, n14818, n14820, n14821,
         n14822, n14824, n14825, n14827, n14828, n14830, n14832, n14833,
         n14834, n14836, n14837, n14839, n14840, n14842, n14844, n14845,
         n14846, n14848, n14849, n14851, n14852, n14854, n14856, n14857,
         n14858, n14860, n14861, n14863, n14864, n14866, n14868, n14869,
         n14870, n14872, n14873, n14875, n14876, n14878, n14880, n14881,
         n14882, n14884, n14885, n14887, n14888, n14890, n14892, n14893,
         n14894, n14896, n14897, n14899, n14900, n14902, n14904, n14905,
         n14906, n14908, n14909, n14911, n14912, n14914, n14916, n14917,
         n14918, n14920, n14921, n14923, n14924, n14926, n14928, n14929,
         n14930, n14932, n14933, n14935, n14936, n14938, n14940, n14941,
         n14942, n14944, n14945, n14947, n14948, n14950, n14952, n14953,
         n14954, n14956, n14957, n14959, n14960, n14962, n14964, n14965,
         n14966, n14968, n14969, n14971, n14972, n14974, n14976, n14977,
         n14978, n14980, n14981, n14983, n14984, n14986, n14988, n14989,
         n14990, n14992, n14993, n14995, n14996, n14998, n15000, n15001,
         n15002, n15004, n15005, n15007, n15008, n15010, n15012, n15013,
         n15014, n15016, n15017, n15019, n15020, n15022, n15024, n15025,
         n15026, n15028, n15029, n15031, n15032, n15034, n15036, n15037,
         n15038, n15040, n15041, n15043, n15044, n15046, n15048, n15049,
         n15050, n15052, n15053, n15055, n15056, n15058, n15060, n15061,
         n15062, n15064, n15065, n15067, n15068, n15070, n15072, n15073,
         n15074, n15076, n15077, n15079, n15080, n15082, n15084, n15085,
         n15086, n15088, n15089, n15091, n15092, n15094, n15096, n15097,
         n15098, n15100, n15101, n15103, n15104, n15106, n15108, n15109,
         n15110, n15112, n15113, n15115, n15116, n15118, n15120, n15121,
         n15122, n15124, n15125, n15127, n15128, n15130, n15132, n15133,
         n15134, n15136, n15137, n15139, n15140, n15142, n15144, n15145,
         n15146, n15148, n15149, n15151, n15152, n15154, n15156, n15157,
         n15158, n15160, n15161, n15163, n15164, n15166, n15168, n15169,
         n15170, n15172, n15173, n15175, n15176, n15178, n15180, n15181,
         n15182, n15184, n15185, n15187, n15188, n15190, n15192, n15193,
         n15194, n15196, n15197, n15199, n15200, n15202, n15204, n15205,
         n15206, n15208, n15209, n15211, n15212, n15214, n15216, n15217,
         n15218, n15220, n15221, n15223, n15224, n15226, n15228, n15229,
         n15230, n15232, n15233, n15235, n15236, n15238, n15240, n15241,
         n15242, n15244, n15245, n15247, n15248, n15250, n15252, n15253,
         n15254, n15256, n15257, n15259, n15260, n15262, n15264, n15265,
         n15266, n15268, n15269, n15271, n15272, n15274, n15276, n15277,
         n15278, n15280, n15281, n15283, n15284, n15286, n15288, n15289,
         n15290, n15292, n15293, n15295, n15296, n15298, n15300, n15301,
         n15302, n15304, n15305, n15307, n15308, n15310, n15312, n15313,
         n15314, n15316, n15317, n15319, n15320, n15322, n15324, n15325,
         n15326, n15328, n15329, n15331, n15332, n15334, n15336, n15337,
         n15338, n15340, n15341, n15343, n15344, n15346, n15348, n15349,
         n15350, n15352, n15353, n15355, n15356, n15358, n15360, n15361,
         n15362, n15364, n15365, n15367, n15368, n15370, n15372, n15373,
         n15374, n15376, n15377, n15379, n15380, n15382, n15384, n15385,
         n15386, n15388, n15389, n15391, n15392, n15394, n15396, n15397,
         n15398, n15400, n15401, n15403, n15404, n15406, n15408, n15409,
         n15410, n15412, n15413, n15415, n15416, n15418, n15420, n15421,
         n15422, n15424, n15425, n15427, n15428, n15430, n15432, n15433,
         n15434, n15436, n15437, n15439, n15440, n15442, n15444, n15445,
         n15446, n15448, n15449, n15451, n15452, n15454, n15456, n15457,
         n15458, n15460, n15461, n15463, n15464, n15466, n15468, n15469,
         n15470, n15472, n15473, n15475, n15476, n15478, n15480, n15481,
         n15482, n15484, n15485, n15487, n15488, n15490, n15492, n15493,
         n15494, n15496, n15497, n15499, n15500, n15502, n15504, n15505,
         n15506, n15508, n15509, n15511, n15512, n15514, n15516, n15517,
         n15518, n15520, n15521, n15523, n15524, n15526, n15528, n15529,
         n15530, n15532, n15533, n15535, n15536, n15538, n15540, n15541,
         n15542, n15544, n15545, n15547, n15548, n15550, n15552, n15553,
         n15554, n15556, n15557, n15559, n15560, n15562, n15564, n15565,
         n15566, n15568, n15569, n15571, n15572, n15574, n15576, n15577,
         n15578, n15580, n15581, n15583, n15584, n15586, n15588, n15589,
         n15590, n15592, n15593, n15595, n15596, n15598, n15600, n15601,
         n15602, n15604, n15605, n15607, n15608, n15610, n15612, n15613,
         n15614, n15616, n15617, n15619, n15620, n15622, n15624, n15625,
         n15626, n15628, n15629, n15631, n15632, n15634, n15636, n15637,
         n15638, n15640, n15641, n15643, n15644, n15646, n15648, n15649,
         n15650, n15652, n15653, n15655, n15656, n15658, n15660, n15661,
         n15662, n15664, n15665, n15667, n15668, n15670, n15672, n15673,
         n15674, n15676, n15677, n15679, n15680, n15682, n15684, n15685,
         n15686, n15688, n15689, n15691, n15692, n15694, n15696, n15697,
         n15698, n15700, n15701, n15703, n15704, n15706, n15708, n15709,
         n15710, n15712, n15713, n15715, n15716, n15718, n15720, n15721,
         n15722, n15724, n15725, n15727, n15728, n15730, n15732, n15733,
         n15734, n15736, n15737, n15739, n15740, n15742, n15744, n15745,
         n15746, n15748, n15749, n15751, n15752, n15754, n15756, n15757,
         n15758, n15760, n15761, n15763, n15764, n15766, n15768, n15769,
         n15770, n15772, n15773, n15775, n15776, n15778, n15780, n15781,
         n15782, n15784, n15785, n15787, n15788, n15790, n15792, n15793,
         n15794, n15796, n15797, n15799, n15800, n15802, n15804, n15805,
         n15806, n15808, n15809, n15811, n15812, n15814, n15816, n15817,
         n15818, n15820, n15821, n15823, n15824, n15826, n15828, n15829,
         n15830, n15832, n15833, n15835, n15836, n15838, n15840, n15841,
         n15842, n15844, n15845, n15847, n15848, n15850, n15852, n15853,
         n15854, n15856, n15857, n15859, n15860, n15862, n15864, n15865,
         n15866, n15868, n15869, n15871, n15872, n15874, n15876, n15877,
         n15878, n15880, n15881, n15883, n15884, n15886, n15888, n15889,
         n15890, n15892, n15893, n15895, n15896, n15898, n15900, n15901,
         n15902, n15904, n15905, n15907, n15908, n15910, n15912, n15913,
         n15914, n15916, n15917, n15919, n15920, n15922, n15924, n15925,
         n15926, n15928, n15929, n15931, n15932, n15934, n15936, n15937,
         n15938, n15940, n15941, n15943, n15944, n15946, n15948, n15949,
         n15950, n15952, n15953, n15955, n15956, n15958, n15960, n15961,
         n15962, n15964, n15965, n15967, n15968, n15970, n15972, n15973,
         n15974, n15976, n15977, n15979, n15980, n15982, n15984, n15985,
         n15986, n15988, n15989, n15991, n15992, n15994, n15996, n15997,
         n15998, n16000, n16001, n16003, n16004, n16006, n16008, n16009,
         n16010, n16012, n16013, n16015, n16016, n16018, n16020, n16021,
         n16022, n16024, n16025, n16027, n16028, n16030, n16032, n16033,
         n16034, n16036, n16037, n16039, n16040, n16042, n16044, n16045,
         n16046, n16048, n16049, n16051, n16052, n16054, n16056, n16057,
         n16058, n16060, n16061, n16063, n16064, n16066, n16068, n16069,
         n16070, n16072, n16073, n16075, n16076, n16078, n16080, n16081,
         n16082, n16084, n16085, n16087, n16088, n16090, n16092, n16093,
         n16094, n16096, n16097, n16099, n16100, n16102, n16104, n16105,
         n16106, n16108, n16109, n16111, n16112, n16114, n16116, n16117,
         n16118, n16120, n16121, n16123, n16124, n16126, n16128, n16129,
         n16130, n16132, n16133, n16135, n16136, n16138, n16140, n16141,
         n16142, n16144, n16145, n16147, n16148, n16150, n16152, n16153,
         n16154, n16156, n16157, n16159, n16160, n16162, n16164, n16165,
         n16166, n16168, n16169, n16171, n16172, n16174, n16176, n16177,
         n16178, n16180, n16181, n16183, n16184, n16186, n16188, n16189,
         n16190, n16192, n16193, n16195, n16196, n16198, n16200, n16201,
         n16202, n16204, n16205, n16207, n16208, n16210, n16212, n16213,
         n16214, n16216, n16217, n16219, n16220, n16222, n16224, n16225,
         n16226, n16228, n16229, n16231, n16232, n16234, n16236, n16237,
         n16238, n16240, n16241, n16243, n16244, n16246, n16248, n16249,
         n16250, n16252, n16253, n16255, n16256, n16258, n16260, n16261,
         n16262, n16264, n16265, n16267, n16268, n16270, n16272, n16273,
         n16274, n16276, n16277, n16279, n16280, n16282, n16284, n16285,
         n16286, n16288, n16289, n16291, n16292, n16294, n16296, n16297,
         n16298, n16300, n16301, n16303, n16304, n16306, n16308, n16309,
         n16310, n16312, n16313, n16315, n16316, n16318, n16320, n16321,
         n16322, n16324, n16325, n16327, n16328, n16330, n16332, n16333,
         n16334, n16336, n16337, n16339, n16340, n16342, n16344, n16345,
         n16346, n16348, n16349, n16351, n16352, n16354, n16356, n16357,
         n16358, n16360, n16361, n16363, n16364, n16366, n16368, n16369,
         n16370, n16372, n16373, n16375, n16376, n16378, n16380, n16381,
         n16382, n16384, n16385, n16387, n16388, n16390, n16392, n16393,
         n16394, n16396, n16397, n16399, n16400, n16402, n16404, n16405,
         n16406, n16408, n16409, n16411, n16412, n16414, n16416, n16417,
         n16418, n16420, n16421, n16423, n16424, n16426, n16428, n16429,
         n16430, n16432, n16433, n16435, n16436, n16438, n16440, n16441,
         n16442, n16444, n16445, n16447, n16448, n16450, n16452, n16453,
         n16454, n16456, n16457, n16459, n16460, n16462, n16464, n16465,
         n16466, n16468, n16469, n16471, n16472, n16474, n16476, n16477,
         n16478, n16480, n16481, n16483, n16484, n16486, n16488, n16489,
         n16490, n16492, n16493, n16495, n16496, n16498, n16500, n16501,
         n16502, n16504, n16505, n16507, n16508, n16510, n16512, n16513,
         n16514, n16516, n16517, n16519, n16520, n16522, n16524, n16525,
         n16526, n16528, n16529, n16531, n16532, n16534, n16536, n16537,
         n16538, n16540, n16541, n16543, n16544, n16546, n16548, n16549,
         n16550, n16552, n16553, n16555, n16556, n16558, n16560, n16561,
         n16562, n16564, n16565, n16567, n16568, n16570, n16572, n16573,
         n16574, n16576, n16577, n16579, n16580, n16582, n16584, n16585,
         n16586, n16588, n16589, n16591, n16592, n16594, n16596, n16597,
         n16598, n16600, n16601, n16603, n16604, n16606, n16608, n16609,
         n16610, n16612, n16613, n16615, n16616, n16618, n16620, n16621,
         n16622, n16624, n16625, n16627, n16628, n16630, n16632, n16633,
         n16634, n16636, n16637, n16639, n16640, n16642, n16644, n16645,
         n16646, n16648, n16649, n16651, n16652, n16654, n16656, n16657,
         n16658, n16660, n16661, n16663, n16664, n16666, n16668, n16669,
         n16670, n16672, n16673, n16675, n16676, n16678, n16680, n16681,
         n16682, n16684, n16685, n16687, n16688, n16690, n16692, n16693,
         n16694, n16696, n16697, n16699, n16700, n16702, n16704, n16705,
         n16706, n16708, n16709, n16711, n16712, n16714, n16716, n16717,
         n16718, n16720, n16721, n16723, n16724, n16726, n16728, n16729,
         n16730, n16732, n16733, n16735, n16736, n16738, n16740, n16741,
         n16742, n16744, n16745, n16747, n16748, n16750, n16752, n16753,
         n16754, n16756, n16757, n16759, n16760, n16762, n16764, n16765,
         n16766, n16768, n16769, n16771, n16772, n16774, n16776, n16777,
         n16778, n16780, n16781, n16783, n16784, n16786, n16788, n16789,
         n16790, n16792, n16793, n16795, n16796, n16798, n16800, n16801,
         n16802, n16804, n16805, n16807, n16808, n16810, n16812, n16813,
         n16814, n16816, n16817, n16819, n16820, n16822, n16824, n16825,
         n16826, n16828, n16829, n16831, n16832, n16834, n16836, n16837,
         n16838, n16840, n16841, n16843, n16844, n16846, n16848, n16849,
         n16850, n16852, n16853, n16855, n16856, n16858, n16860, n16861,
         n16862, n16864, n16865, n16867, n16868, n16870, n16872, n16873,
         n16874, n16876, n16877, n16879, n16880, n16882, n16884, n16885,
         n16886, n16888, n16889, n16891, n16892, n16894, n16896, n16897,
         n16898, n16900, n16901, n16903, n16904, n16906, n16908, n16909,
         n16910, n16912, n16913, n16915, n16916, n16918, n16920, n16921,
         n16922, n16924, n16925, n16927, n16928, n16930, n16932, n16933,
         n16934, n16936, n16937, n16939, n16940, n16942, n16944, n16945,
         n16946, n16948, n16949, n16951, n16952, n16954, n16956, n16957,
         n16958, n16960, n16961, n16963, n16964, n16966, n16968, n16969,
         n16970, n16972, n16973, n16975, n16976, n16978, n16980, n16981,
         n16982, n16984, n16985, n16987, n16988, n16990, n16992, n16993,
         n16994, n16996, n16997, n16999, n17000, n17002, n17004, n17005,
         n17006, n17008, n17009, n17011, n17012, n17014, n17016, n17017,
         n17018, n17020, n17021, n17023, n17024, n17026, n17028, n17029,
         n17030, n17032, n17033, n17035, n17036, n17038, n17040, n17041,
         n17042, n17044, n17045, n17047, n17048, n17050, n17052, n17053,
         n17054, n17056, n17057, n17059, n17060, n17062, n17064, n17065,
         n17066, n17068, n17069, n17071, n17072, n17074, n17076, n17077,
         n17078, n17080, n17081, n17083, n17084, n17086, n17088, n17089,
         n17090, n17092, n17093, n17095, n17096, n17098, n17100, n17101,
         n17102, n17104, n17105, n17107, n17108, n17110, n17112, n17113,
         n17114, n17116, n17117, n17119, n17120, n17122, n17124, n17125,
         n17126, n17128, n17129, n17131, n17132, n17134, n17136, n17137,
         n17138, n17140, n17141, n17143, n17144, n17146, n17148, n17149,
         n17150, n17152, n17153, n17155, n17156, n17158, n17160, n17161,
         n17162, n17164, n17165, n17167, n17168, n17170, n17172, n17173,
         n17174, n17176, n17177, n17179, n17180, n17182, n17184, n17185,
         n17186, n17188, n17189, n17191, n17192, n17194, n17196, n17197,
         n17198, n17200, n17201, n17203, n17204, n17206, n17208, n17209,
         n17210, n17212, n17213, n17215, n17216, n17218, n17220, n17221,
         n17222, n17224, n17225, n17227, n17228, n17230, n17232, n17233,
         n17234, n17236, n17237, n17239, n17240, n17242, n17244, n17245,
         n17246, n17248, n17249, n17251, n17252, n17254, n17256, n17257,
         n17258, n17260, n17261, n17263, n17264, n17266, n17268, n17269,
         n17270, n17272, n17273, n17275, n17276, n17278, n17280, n17281,
         n17282, n17284, n17285, n17287, n17288, n17290, n17292, n17293,
         n17294, n17296, n17297, n17299, n17300, n17302, n17304, n17305,
         n17306, n17308, n17309, n17311, n17312, n17314, n17316, n17317,
         n17318, n17320, n17321, n17323, n17324, n17326, n17328, n17329,
         n17330, n17332, n17333, n17335, n17336, n17338, n17340, n17341,
         n17342, n17344, n17345, n17347, n17348, n17350, n17352, n17353,
         n17354, n17356, n17357, n17359, n17360, n17362, n17364, n17365,
         n17366, n17368, n17369, n17371, n17372, n17374, n17376, n17377,
         n17378, n17380, n17381, n17383, n17384, n17386, n17388, n17389,
         n17390, n17392, n17393, n17395, n17396, n17398, n17400, n17401,
         n17402, n17404, n17405, n17407, n17408, n17410, n17412, n17413,
         n17414, n17416, n17417, n17419, n17420, n17422, n17424, n17425,
         n17426, n17428, n17429, n17431, n17432, n17434, n17436, n17437,
         n17438, n17440, n17441, n17443, n17444, n17446, n17448, n17449,
         n17450, n17452, n17453, n17455, n17456, n17458, n17460, n17461,
         n17462, n17464, n17465, n17467, n17468, n17470, n17472, n17473,
         n17474, n17476, n17477, n17479, n17480, n17482, n17484, n17485,
         n17486, n17488, n17489, n17491, n17492, n17494, n17496, n17497,
         n17498, n17500, n17501, n17503, n17504, n17506, n17508, n17509,
         n17510, n17512, n17513, n17515, n17516, n17518, n17520, n17521,
         n17522, n17524, n17525, n17527, n17528, n17530, n17532, n17533,
         n17534, n17536, n17537, n17539, n17540, n17542, n17544, n17545,
         n17546, n17548, n17549, n17551, n17552, n17554, n17556, n17557,
         n17558, n17560, n17561, n17563, n17564, n17566, n17568, n17569,
         n17570, n17572, n17573, n17575, n17576, n17578, n17580, n17581,
         n17582, n17584, n17585, n17587, n17588, n17590, n17592, n17593,
         n17594, n17596, n17597, n17599, n17600, n17602, n17604, n17605,
         n17606, n17608, n17609, n17611, n17612, n17614, n17616, n17617,
         n17618, n17620, n17621, n17623, n17624, n17626, n17628, n17629,
         n17630, n17632, n17633, n17635, n17636, n17638, n17640, n17641,
         n17642, n17644, n17645, n17647, n17648, n17650, n17652, n17653,
         n17654, n17656, n17657, n17659, n17660, n17662, n17664, n17665,
         n17666, n17668, n17669, n17671, n17672, n17674, n17676, n17677,
         n17678, n17680, n17681, n17683, n17684, n17686, n17688, n17689,
         n17690, n17692, n17693, n17695, n17696, n17698, n17700, n17701,
         n17702, n17704, n17705, n17707, n17708, n17710, n17712, n17713,
         n17714, n17716, n17717, n17719, n17720, n17722, n17724, n17725,
         n17726, n17728, n17729, n17731, n17732, n17734, n17736, n17737,
         n17738, n17740, n17741, n17743, n17744, n17746, n17748, n17749,
         n17750, n17752, n17753, n17755, n17756, n17758, n17760, n17761,
         n17762, n17764, n17765, n17767, n17768, n17770, n17772, n17773,
         n17774, n17776, n17777, n17779, n17780, n17782, n17784, n17785,
         n17786, n17788, n17789, n17791, n17792, n17794, n17796, n17797,
         n17798, n17800, n17801, n17803, n17804, n17806, n17808, n17809,
         n17810, n17812, n17813, n17815, n17816, n17818, n17820, n17821,
         n17822, n17824, n17825, n17827, n17828, n17830, n17832, n17833,
         n17834, n17836, n17837, n17839, n17840, n17842, n17844, n17845,
         n17846, n17848, n17849, n17851, n17852, n17854, n17856, n17857,
         n17858, n17860, n17861, n17863, n17864, n17866, n17868, n17869,
         n17870, n17872, n17873, n17875, n17876, n17878, n17880, n17881,
         n17882, n17884, n17885, n17887, n17888, n17890, n17892, n17893,
         n17894, n17896, n17897, n17899, n17900, n17902, n17904, n17905,
         n17906, n17908, n17909, n17911, n17912, n17914, n17916, n17917,
         n17918, n17920, n17921, n17923, n17924, n17926, n17928, n17929,
         n17930, n17932, n17933, n17935, n17936, n17938, n17940, n17941,
         n17942, n17944, n17945, n17947, n17948, n17950, n17952, n17953,
         n17954, n17956, n17957, n17959, n17960, n17962, n17964, n17965,
         n17966, n17968, n17969, n17971, n17972, n17974, n17976, n17977,
         n17978, n17980, n17981, n17983, n17984, n17986, n17988, n17989,
         n17990, n17992, n17993, n17995, n17996, n17998, n18000, n18001,
         n18002, n18004, n18005, n18007, n18008, n18010, n18012, n18013,
         n18014, n18016, n18017, n18019, n18020, n18022, n18024, n18025,
         n18026, n18028, n18029, n18031, n18032, n18034, n18036, n18037,
         n18038, n18040, n18041, n18043, n18044, n18046, n18048, n18049,
         n18050, n18052, n18053, n18055, n18056, n18058, n18060, n18061,
         n18062, n18064, n18065, n18067, n18068, n18070, n18072, n18073,
         n18074, n18076, n18077, n18079, n18080, n18082, n18084, n18085,
         n18086, n18088, n18089, n18091, n18092, n18094, n18096, n18097,
         n18098, n18100, n18101, n18103, n18104, n18106, n18108, n18109,
         n18110, n18112, n18113, n18115, n18116, n18118, n18120, n18121,
         n18122, n18124, n18125, n18127, n18128, n18130, n18132, n18133,
         n18134, n18136, n18137, n18139, n18140, n18142, n18144, n18145,
         n18146, n18148, n18149, n18151, n18152, n18154, n18156, n18157,
         n18158, n18160, n18161, n18163, n18164, n18166, n18168, n18169,
         n18170, n18172, n18173, n18175, n18176, n18178, n18180, n18181,
         n18182, n18184, n18185, n18187, n18188, n18190, n18192, n18193,
         n18194, n18196, n18197, n18199, n18200, n18202, n18204, n18205,
         n18206, n18208, n18209, n18211, n18212, n18214, n18216, n18217,
         n18218, n18220, n18221, n18223, n18224, n18226, n18228, n18229,
         n18232, n18235, n18236, n18238, n18240, n18241, n18244, n18247,
         n18250, n18252, n18253, n18256, n18259, n18262, n18264, n18265,
         n18268, n18271, n18274, n18276, n18277, n18280, n18283, n18286,
         n18288, n18289, n18292, n18295, n18298, n18300, n18301, n18304,
         n18307, n18310, n18312, n18313, n18316, n18319, n18322, n18324,
         n18325, n18328, n18331, n18334, n18336, n18337, n18340, n18343,
         n18346, n18348, n18349, n18352, n18355, n18358, n18360, n18361,
         n18364, n18367, n18370, n18372, n18373, n18376, n18379, n18382,
         n18384, n18385, n18388, n18391, n18394, n18396, n18397, n18400,
         n18403, n18406, n18408, n18409, n18412, n18415, n18418, n18420,
         n18421, n18424, n18427, n18430, n18432, n18433, n18436, n18439,
         n18442, n18444, n18445, n18448, n18451, n18454, n18456, n18457,
         n18460, n18463, n18466, n18468, n18469, n18472, n18475, n18478,
         n18480, n18481, n18484, n18487, n18490, n18492, n18493, n18496,
         n18499, n18502, n18504, n18505, n18508, n18511, n18514, n18516,
         n18517, n18520, n18523, n18526, n18528, n18529, n18532, n18535,
         n18538, n18540, n18541, n18544, n18547, n18550, n18552, n18553,
         n18556, n18559, n18562, n18564, n18565, n18568, n18571, n18574,
         n18576, n18577, n18580, n18583, n18586, n18588, n18589, n18592,
         n18595, n18598, n18600, n18601, n18604, n18607, n18610, n18612,
         n18613, n18616, n18619, n18622, n18624, n18625, n18628, n18631,
         n18634, n18636, n18637, n18640, n18643, n18646, n18648, n18649,
         n18652, n18655, n18658, n18660, n18661, n18664, n18667, n18670,
         n18672, n18673, n18676, n18679, n18682, n18684, n18685, n18688,
         n18691, n18694, n18696, n18697, n18700, n18703, n18706, n18708,
         n18709, n18712, n18715, n18718, n18720, n18721, n18724, n18727,
         n18730, n18732, n18733, n18736, n18739, n18742, n18744, n18745,
         n18748, n18751, n18754, n18756, n18757, n18760, n18763, n18766,
         n18768, n18769, n18772, n18775, n18778, n18780, n18781, n18784,
         n18787, n18790, n18792, n18793, n18796, n18799, n18802, n18804,
         n18805, n18808, n18811, n18814, n18816, n18817, n18820, n18823,
         n18826, n18828, n18829, n18832, n18835, n18838, n18840, n18841,
         n18844, n18847, n18850, n18852, n18853, n18856, n18859, n18862,
         n18864, n18865, n18868, n18871, n18874, n18876, n18877, n18880,
         n18883, n18886, n18888, n18889, n18892, n18895, n18898, n18900,
         n18901, n18904, n18907, n18910, n18912, n18913, n18916, n18919,
         n18922, n18924, n18925, n18928, n18931, n18934, n18936, n18937,
         n18940, n18943, n18946, n18948, n18949, n18952, n18955, n18958,
         n18960, n18961, n18964, n18967, n18970, n18972, n18973, n18976,
         n18979, n18982, n18984, n18985, n18988, n18991, n18994, n18996,
         n18997, n19000, n19003, n19006, n19008, n19009, n19012, n19015,
         n19018, n19020, n19021, n19024, n19027, n19030, n19032, n19033,
         n19036, n19039, n19042, n19044, n19045, n19048, n19051, n19054,
         n19056, n19057, n19060, n19063, n19066, n19068, n19069, n19072,
         n19075, n19078, n19080, n19081, n19084, n19087, n19090, n19092,
         n19093, n19096, n19099, n19102, n19104, n19105, n19108, n19111,
         n19114, n19116, n19117, n19120, n19123, n19126, n19128, n19129,
         n19132, n19135, n19138, n19140, n19141, n19144, n19147, n19150,
         n19152, n19153, n19156, n19158, n19159, n19161, n19162, n19164,
         n19165, n19167, n19168, n19170, n19171, n19173, n19174, n19176,
         n19177, n19179, n19180, n19181, n19182, n19184, n19185, n19186,
         n19187, n19189, n19191, n19193, n19195, n19197, n19199, n19202,
         n19203, n19207, n19208, n19210, n19211, n19214, n19215, n19218,
         n19219, n19222, n19223, n19226, n19227, n19230, n19231, n19234,
         n19235, n19238, n19239, n19240, n19241, n19243, n19247, n19249,
         n19251, n19252, n19253, n19255, n19256, n19257, n19259, n19260,
         n19261, n19263, n19264, n19265, n19267, n19268, n19269, n19271,
         n19272, n19273, n19275, n19276, n19277, n19278, n19281, n19283,
         n19284, n19285, n19286, n19287, n19290, n19292, n19293, n19294,
         n19295, n19296, n19299, n19300, n19301, n19302, n19305, n19306,
         n19307, n19308, n19311, n19312, n19313, n19314, n19317, n19318,
         n19319, n19320, n19323, n19324, n19325, n19326, n19329, n19330,
         n19331, n19332, n19334, n19335, n19336, n19338, n19339, n19340,
         n19341, n19343, n19344, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19528, n19533, n19534, n19535, n19536, n19537,
         n19538, n19543, n19544, n19545, n19546, n19547, n19548, n19553,
         n19554, n19555, n19556, n19557, n19558, n19563, n19564, n19565,
         n19566, n19567, n19568, n19573, n19574, n19575, n19576, n19577,
         n19578, n19583, n19584, n19585, n19586, n19587, n19588, n19593,
         n19594, n19595, n19596, n19597, n19598, n19603, n19604, n19605,
         n19606, n19607, n19608, n19613, n19614, n19615, n19616, n19617,
         n19618, n19623, n19624, n19625, n19626, n19627, n19628, n19633,
         n19634, n19635, n19636, n19637, n19638, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19654, n19655, n19656, n19657,
         n19658, n19660, n19665, n19666, n19667, n19668, n19669, n19670,
         n19675, n19676, n19677, n19678, n19679, n19680, n19685, n19686,
         n19687, n19688, n19689, n19690, n19695, n19696, n19697, n19698,
         n19699, n19700, n19705, n19706, n19707, n19708, n19709, n19710,
         n19715, n19716, n19717, n19718, n19719, n19720, n19725, n19726,
         n19727, n19728, n19729, n19731, n19736, n19737, n19738, n19739,
         n19740, n19741, n19746, n19747, n19748, n19749, n19750, n19751,
         n19756, n19757, n19758, n19759, n19760, n19761, n19766, n19767,
         n19768, n19769, n19770, n19771, n19776, n19777, n19778, n19779,
         n19780, n19781, n19786, n19787, n19788, n19789, n19790, n19791,
         n19796, n19797, n19798, n19799, n19800, n19801, n19806, n19807,
         n19808, n19810, n19811, n19816, n19817, n19818, n19819, n19820,
         n19821, n19826, n19827, n19828, n19829, n19830, n19831, n19836,
         n19837, n19838, n19839, n19840, n19841, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19857, n19858, n19859, n19860,
         n19861, n19862, n19867, n19868, n19869, n19870, n19871, n19872,
         n19877, n19878, n19879, n19880, n19881, n19882, n19887, n19888,
         n19889, n19890, n19891, n19892, n19897, n19898, n19899, n19900,
         n19901, n19902, n19907, n19908, n19909, n19910, n19911, n19912,
         n19917, n19918, n19919, n19920, n19921, n19922, n19927, n19928,
         n19929, n19930, n19931, n19932, n19937, n19938, n19939, n19940,
         n19941, n19942, n19947, n19948, n19949, n19950, n19951, n19952,
         n19957, n19958, n19959, n19960, n19961, n19962, n19967, n19968,
         n19969, n19970, n19971, n19972, n19977, n19978, n19979, n19980,
         n19981, n19982, n19987, n19988, n19989, n19990, n19991, n19993,
         n19998, n19999, n20000, n20001, n20002, n20003, n20008, n20009,
         n20010, n20011, n20012, n20014, n20015, n20020, n20021, n20022,
         n20023, n20024, n20025, n20030, n20031, n20032, n20033, n20034,
         n20035, n20040, n20041, n20042, n20043, n20044, n20045, n20050,
         n20051, n20052, n20053, n20054, n20055, n20060, n20061, n20062,
         n20063, n20064, n20065, n20070, n20071, n20072, n20073, n20074,
         n20075, n20080, n20081, n20082, n20083, n20084, n20085, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20101, n20102,
         n20103, n20104, n20105, n20106, n20111, n20112, n20113, n20114,
         n20115, n20117, n20122, n20123, n20124, n20125, n20126, n20127,
         n20132, n20133, n20134, n20135, n20136, n20137, n20142, n20143,
         n20144, n20145, n20146, n20147, n20152, n20153, n20154, n20155,
         n20156, n20157, n20162, n20163, n20164, n20165, n20166, n20167,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20183,
         n20184, n20185, n20186, n20187, n20189, n20194, n20195, n20196,
         n20197, n20198, n20199, n20204, n20205, n20206, n20207, n20208,
         n20209, n20214, n20215, n20216, n20217, n20218, n20219, n20224,
         n20225, n20226, n20227, n20228, n20229, n20234, n20235, n20236,
         n20237, n20238, n20239, n20244, n20245, n20246, n20247, n20248,
         n20249, n20254, n20255, n20256, n20257, n20258, n20260, n20266,
         n20267, n20268, n20269, n20270, n20271, n20276, n20277, n20278,
         n20279, n20280, n20281, n20286, n20287, n20288, n20289, n20290,
         n20291, n20296, n20297, n20298, n20299, n20300, n20301, n20381,
         n20382, n20388, n20389, n20390, n20391, n20392, n20393, n20398,
         n20399, n20400, n20401, n20402, n20403, n20408, n20409, n20410,
         n20411, n20412, n20413, n20424, n20429, n20430, n20431, n20432,
         n20433, n20434, n20439, n20440, n20441, n20442, n20443, n20444,
         n20449, n20450, n20451, n20452, n20453, n20455, n20460, n20461,
         n20462, n20463, n20464, n20466, n20471, n20472, n20473, n20474,
         n20475, n20476, n20481, n20482, n20483, n20484, n20485, n20486,
         n20491, n20492, n20493, n20494, n20495, n20496, n20501, n20502,
         n20503, n20504, n20505, n20506, n20792, n20797, n20798, n20799,
         n20800, n20801, n20802, n20807, n20808, n20809, n20810, n20811,
         n20813, n20818, n20819, n20820, n20821, n20822, n20823, n20828,
         n20829, n20830, n20831, n20832, n20834, n20839, n20840, n20841,
         n20842, n20843, n20845, n20850, n20851, n20852, n20853, n20854,
         n20855, n20860, n20861, n20862, n20863, n20864, n20865, n20870,
         n20871, n20872, n20873, n20874, n20876, n20877, n20882, n20883,
         n20884, n20885, n20886, n20887, n20892, n20893, n20894, n20895,
         n20896, n20897, n20902, n20903, n20904, n20905, n20906, n20908,
         n20913, n20914, n20915, n20916, n20917, n20918, n20923, n20924,
         n20925, n20926, n20927, n20929, n20934, n20935, n20936, n20937,
         n20938, n20939, n20944, n20945, n20946, n20947, n20948, n20949,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20965,
         n20966, n20967, n20968, n20969, n20970, n20975, n20976, n20977,
         n20978, n20979, n20981, n20986, n20987, n20988, n20989, n20990,
         n20991, n20996, n20997, n20998, n20999, n21000, n21001, n21006,
         n21007, n21008, n21009, n21010, n21011, n21016, n21017, n21018,
         n21019, n21020, n21021, n21026, n21027, n21028, n21029, n21030,
         n21032, n21037, n21038, n21039, n21040, n21041, n21042, n21047,
         n21048, n21049, n21050, n21051, n21052, n21057, n21058, n21059,
         n21060, n21061, n21062, n21067, n21068, n21069, n21070, n21071,
         n21072, n21077, n21078, n21079, n21080, n21081, n21082, n21087,
         n21088, n21089, n21090, n21091, n21092, n21097, n21098, n21099,
         n21100, n21101, n21102, n21107, n21108, n21109, n21110, n21111,
         n21112, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21128, n21129, n21130, n21131, n21132, n21133, n21138, n21139,
         n21140, n21141, n21142, n21143, n21148, n21149, n21150, n21151,
         n21152, n21153, n21158, n21159, n21160, n21161, n21162, n21163,
         n21168, n21169, n21170, n21171, n21172, n21173, n21178, n21179,
         n21180, n21181, n21182, n21183, n21188, n21189, n21190, n21191,
         n21192, n21193, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21209, n21210, n21211, n21212, n21213, n21214, n21219,
         n21220, n21221, n21222, n21223, n21224, n21229, n21230, n21231,
         n21232, n21233, n21234, n21239, n21240, n21241, n21242, n21243,
         n21244, n21249, n21250, n21251, n21252, n21253, n21254, n21259,
         n21260, n21261, n21262, n21263, n21264, n21269, n21270, n21271,
         n21272, n21273, n21274, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21290, n21291, n21292, n21293, n21294, n21295,
         n21300, n21301, n21302, n21303, n21304, n21305, n21310, n21311,
         n21312, n21313, n21314, n21315, n21320, n21321, n21322, n21323,
         n21324, n21325, n21330, n21331, n21332, n21333, n21334, n21335,
         n21340, n21341, n21342, n21343, n21344, n21345, n21350, n21351,
         n21352, n21353, n21354, n21355, n21360, n21361, n21362, n21363,
         n21364, n21365, n21370, n21371, n21372, n21373, n21374, n21375,
         n21380, n21381, n21382, n21383, n21384, n21385, n21390, n21391,
         n21392, n21393, n21394, n21395, n21400, n21401, n21402, n21403,
         n21404, n21405, n21410, n21411, n21412, n21413, n21414, n21415,
         n21420, n21421, n21422, n21423, n21424, n21425, n21430, n21431,
         n21432, n21433, n21434, n21435, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21451, n21452, n21453, n21454, n21455,
         n21456, n21461, n21462, n21463, n21464, n21465, n21466, n21471,
         n21472, n21473, n21474, n21475, n21476, n21481, n21482, n21483,
         n21484, n21485, n21486, n21491, n21492, n21493, n21494, n21495,
         n21496, n21501, n21502, n21503, n21504, n21505, n21506, n21511,
         n21512, n21513, n21514, n21515, n21516, n21521, n21522, n21523,
         n21524, n21525, n21526, n21531, n21532, n21533, n21534, n21535,
         n21536, n21541, n21542, n21543, n21544, n21545, n21546, n21551,
         n21552, n21553, n21554, n21555, n21556, n21561, n21562, n21563,
         n21564, n21565, n21566, n21571, n21572, n21573, n21574, n21575,
         n21576, n21581, n21582, n21583, n21584, n21585, n21586, n21591,
         n21592, n21593, n21594, n21595, n21596, n21601, n21602, n21603,
         n21604, n21605, n21607, n21608, n21613, n21614, n21615, n21616,
         n21617, n21618, n21623, n21624, n21625, n21626, n21627, n21628,
         n21633, n21634, n21635, n21636, n21637, n21638, n21643, n21644,
         n21645, n21646, n21647, n21648, n21653, n21654, n21655, n21656,
         n21657, n21658, n21663, n21664, n21665, n21666, n21667, n21668,
         n21673, n21674, n21675, n21676, n21677, n21678, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21694, n21695, n21696,
         n21697, n21698, n21699, n21704, n21705, n21706, n21707, n21708,
         n21709, n21714, n21715, n21716, n21717, n21718, n21719, n21724,
         n21725, n21726, n21727, n21728, n21729, n21734, n21735, n21736,
         n21737, n21738, n21739, n21744, n21745, n21746, n21747, n21748,
         n21749, n21754, n21755, n21756, n21757, n21758, n21759, n21764,
         n21765, n21766, n21767, n21768, n21769, n21774, n21775, n21776,
         n21777, n21778, n21779, n21784, n21785, n21786, n21787, n21788,
         n21790, n21795, n21796, n21797, n21798, n21799, n21801, n21806,
         n21807, n21808, n21809, n21810, n21811, n21816, n21817, n21818,
         n21819, n21820, n21821, n21826, n21827, n21828, n21829, n21830,
         n21831, n21836, n21837, n21838, n21839, n21840, n21841, n21846,
         n21847, n21848, n21849, n21850, n21851, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21867, n21868, n21869, n21870,
         n21871, n21872, n21877, n21878, n21879, n21880, n21881, n21882,
         n21887, n21888, n21889, n21890, n21891, n21892, n21897, n21898,
         n21899, n21900, n21901, n21902, n21907, n21908, n21909, n21910,
         n21911, n21913, n21918, n21919, n21920, n21921, n21922, n21923,
         n21928, n21929, n21930, n21931, n21932, n21933, n21938, n21939,
         n21940, n21941, n21942, n21943, n21948, n21949, n21950, n21951,
         n21952, n21953, n21958, n21959, n21960, n21961, n21962, n21963,
         n21968, n21969, n21970, n21971, n21972, n21973, n21978, n21979,
         n21980, n21981, n21982, n21983, n21988, n21989, n21990, n21991,
         n21992, n21993, n21998, n21999, n22000, n22001, n22002, n22003,
         n22008, n22009, n22010, n22011, n22012, n22013, n22018, n22019,
         n22020, n22021, n22022, n22023, n22028, n22029, n22030, n22031,
         n22032, n22033, n22038, n22039, n22040, n22041, n22042, n22043,
         n22048, n22049, n22050, n22051, n22052, n22053, n22058, n22059,
         n22060, n22061, n22062, n22063, n22068, n22069, n22070, n22071,
         n22072, n22073, n22078, n22079, n22080, n22081, n22082, n22084,
         n22089, n22090, n22091, n22092, n22093, n22094, n22098, n22316,
         n22317, n22318, n22319, n22320, n22321, n22326, n22327, n22328,
         n22329, n22330, n22331, n22336, n22337, n22338, n22339, n22340,
         n22341, n22346, n22347, n22348, n22349, n22350, n22351, n22356,
         n22357, n22358, n22359, n22360, n22361, n22366, n22367, n22368,
         n22369, n22370, n22371, n22376, n22377, n22378, n22379, n22380,
         n22381, n22386, n22387, n22388, n22389, n22390, n22391, n22396,
         n22397, n22398, n22399, n22400, n22401, n22406, n22407, n22408,
         n22409, n22410, n22411, n22416, n22417, n22418, n22419, n22420,
         n22421, n22426, n22427, n22428, n22429, n22430, n22431, n22436,
         n22437, n22438, n22439, n22440, n22441, n22446, n22447, n22448,
         n22449, n22450, n22451, n22456, n22457, n22458, n22459, n22460,
         n22461, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22478, n22479, n22480, n22481, n22482, n22483, n22488,
         n22489, n22490, n22491, n22492, n22493, n22498, n22499, n22500,
         n22501, n22502, n22503, n22508, n22509, n22510, n22511, n22512,
         n22513, n22518, n22519, n22520, n22521, n22522, n22523, n22528,
         n22529, n22530, n22531, n22532, n22533, n22538, n22539, n22540,
         n22541, n22542, n22543, n22548, n22549, n22550, n22551, n22552,
         n22553, n22554, n22559, n22560, n22561, n22562, n22563, n22564,
         n22569, n22570, n22571, n22572, n22573, n22574, n22579, n22580,
         n22581, n22582, n22583, n22584, n22589, n22590, n22591, n22592,
         n22593, n22594, n22599, n22600, n22601, n22602, n22603, n22604,
         n22609, n22610, n22611, n22612, n22613, n22614, n22619, n22620,
         n22621, n22622, n22623, n22624, n22629, n22630, n22631, n22632,
         n22633, n22634, n22635, n22640, n22641, n22642, n22643, n22644,
         n22645, n22650, n22651, n22652, n22653, n22654, n22655, n22660,
         n22661, n22662, n22663, n22664, n22665, n22670, n22671, n22672,
         n22673, n22674, n22675, n22680, n22681, n22682, n22683, n22684,
         n22685, n22690, n22691, n22692, n22693, n22694, n22695, n22700,
         n22701, n22702, n22703, n22704, n22705, n22710, n22711, n22712,
         n22713, n22714, n22715, n22720, n22721, n22722, n22723, n22724,
         n22725, n22730, n22731, n22732, n22733, n22734, n22735, n22740,
         n22741, n22742, n22743, n22744, n22745, n22750, n22751, n22752,
         n22753, n22754, n22755, n22760, n22761, n22762, n22763, n22764,
         n22765, n22770, n22771, n22772, n22773, n22774, n22775, n22780,
         n22781, n22782, n22783, n22784, n22785, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22801, n22802, n22803, n22804,
         n22805, n22806, n22811, n22812, n22813, n22814, n22815, n22816,
         n22821, n22822, n22823, n22824, n22825, n22826, n22831, n22832,
         n22833, n22834, n22835, n22836, n22841, n22842, n22843, n22844,
         n22845, n22846, n22851, n22852, n22853, n22854, n22855, n22857,
         n22862, n22863, n22864, n22865, n22866, n22867, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22882,
         n22883, n22884, n22885, n22886, n22887, n22893, n22894, n22895,
         n22896, n22897, n22898, n22903, n22904, n22905, n22906, n22907,
         n22908, n22913, n22914, n22915, n22916, n22917, n22918, n22923,
         n22924, n22925, n22926, n22927, n22928, n22933, n22934, n22935,
         n22936, n22937, n22938, n22943, n22944, n22945, n22946, n22947,
         n22948, n22953, n22954, n22955, n22956, n22957, n22958, n22963,
         n22964, n22965, n22966, n22967, n22968, n22973, n22974, n22975,
         n22976, n22977, n22978, n22983, n22984, n22985, n22986, n22987,
         n22988, n22993, n22994, n22995, n22996, n22997, n22998, n23003,
         n23004, n23005, n23006, n23007, n23008, n23013, n23014, n23015,
         n23016, n23017, n23018, n23023, n23024, n23025, n23026, n23027,
         n23028, n23033, n23034, n23035, n23036, n23037, n23038, n23043,
         n23044, n23045, n23046, n23047, n23048, n23053, n23054, n23055,
         n23056, n23057, n23058, n23063, n23064, n23065, n23066, n23067,
         n23068, n23073, n23074, n23075, n23076, n23077, n23078, n23083,
         n23084, n23085, n23086, n23087, n23088, n23093, n23094, n23095,
         n23096, n23097, n23098, n23103, n23104, n23105, n23106, n23107,
         n23108, n23113, n23114, n23115, n23116, n23117, n23118, n23123,
         n23124, n23125, n23126, n23127, n23128, n23133, n23134, n23135,
         n23136, n23137, n23138, n23143, n23144, n23145, n23146, n23147,
         n23148, n23153, n23154, n23155, n23156, n23157, n23158, n23163,
         n23164, n23165, n23166, n23167, n23168, n23173, n23174, n23175,
         n23176, n23177, n23178, n23183, n23184, n23185, n23186, n23187,
         n23188, n23193, n23194, n23195, n23196, n23197, n23198, n23203,
         n23204, n23205, n23206, n23207, n23208, n23213, n23214, n23215,
         n23216, n23217, n23218, n23223, n23224, n23225, n23226, n23227,
         n23228, n23233, n23234, n23235, n23236, n23237, n23238, n23243,
         n23244, n23245, n23246, n23247, n23248, n23253, n23254, n23255,
         n23256, n23257, n23258, n23263, n23264, n23265, n23266, n23267,
         n23269, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
         n23285, n23286, n23287, n23288, n23289, n23290, n23295, n23296,
         n23297, n23298, n23299, n23300, n23305, n23306, n23307, n23308,
         n23309, n23311, n23316, n23317, n23318, n23319, n23320, n23321,
         n23326, n23327, n23328, n23329, n23330, n23331, n23336, n23337,
         n23338, n23339, n23340, n23342, n23347, n23348, n23349, n23350,
         n23351, n23352, n23357, n23358, n23359, n23360, n23361, n23362,
         n23448, n23449, n23450, n23451, n23452, n23453, n23458, n23459,
         n23460, n23461, n23462, n23463, n23468, n23469, n23470, n23471,
         n23472, n23473, n23478, n23479, n23480, n23481, n23482, n23483,
         n23488, n23489, n23490, n23491, n23492, n23493, n23498, n23499,
         n23500, n23501, n23502, n23503, n23508, n23509, n23510, n23511,
         n23512, n23513, n23518, n23519, n23520, n23521, n23522, n23523,
         n23528, n23529, n23530, n23531, n23532, n23533, n23538, n23539,
         n23540, n23541, n23542, n23543, n23548, n23549, n23550, n235510,
         n235520, n235530, n235580, n235590, n235600, n235610, n235620, n23563,
         n23568, n23569, n23570, n23571, n23572, n23574, n23579, n23580,
         n23581, n23582, n23583, n23585, n23590, n23591, n23592, n23593,
         n23594, n23595, n23600, n23601, n23602, n23603, n23604, n23605,
         n23606, n23611, n23612, n23613, n23614, n23615, n23616, n23621,
         n23622, n23623, n23624, n23625, n23626, n23631, n23632, n23633,
         n23634, n23635, n23636, n23641, n23642, n23643, n23644, n23645,
         n23646, n23651, n23652, n23653, n23654, n23655, n23656, n23661,
         n23662, n23663, n23664, n23665, n23666, n23671, n23672, n23673,
         n23674, n23675, n23676, n23681, n23682, n23683, n23684, n23685,
         n23686, n23687, n23688, n23693, n23694, n23695, n23696, n23697,
         n23698, n23703, n23704, n23705, n23706, n23707, n23708, n23713,
         n23714, n23715, n23716, n23717, n23718, n23723, n23724, n23725,
         n23726, n23727, n23728, n23733, n23734, n23735, n23736, n23737,
         n23738, n23743, n23744, n23745, n23746, n23747, n23748, n23753,
         n23754, n23755, n23756, n23757, n23758, n23763, n23764, n23765,
         n23766, n23767, n23768, n23774, n23775, n23776, n23777, n23778,
         n23779, n23784, n23785, n23786, n23787, n23788, n23789, n23804,
         n23805, n23806, n23807, n23808, n23809, n23814, n23815, n23816,
         n23817, n23818, n23819, n23834, n23835, n23836, n23837, n23838,
         n23839, n23844, n23845, n23846, n23847, n23848, n23849, n23854,
         n23855, n23856, n23857, n23858, n23859, n23934, n23935, n23936,
         n23937, n23938, n23939, n23944, n23945, n23946, n23947, n23948,
         n23949, n23954, n23955, n23956, n23957, n23958, n23959, n23964,
         n23965, n23966, n23967, n23968, n23969, n23974, n23975, n23976,
         n23977, n23978, n23979, n23984, n23985, n23986, n23987, n23988,
         n23989, n23994, n23995, n23996, n23997, n23998, n23999, n24004,
         n24005, n24006, n24007, n24008, n24009, n24010, n24015, n24016,
         n24017, n24018, n24019, n24020, n24025, n24026, n24027, n24028,
         n24029, n24030, n24035, n24036, n24037, n24038, n24039, n24040,
         n24045, n24046, n24047, n24048, n24049, n24050, n24055, n24056,
         n24057, n24058, n24059, n24060, n24065, n24066, n24067, n24068,
         n24069, n24070, n24075, n24076, n24077, n24078, n24079, n24080,
         n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24096,
         n24097, n24098, n24099, n24100, n24101, n24106, n24107, n24108,
         n24109, n24110, n24111, n24116, n24117, n24118, n24119, n24120,
         n24121, n24126, n24127, n24128, n24129, n24130, n24131, n24136,
         n24137, n24138, n24139, n24140, n24142, n24147, n24148, n24149,
         n24150, n24151, n24152, n24157, n24158, n24159, n24160, n24161,
         n24162, n24167, n24168, n24169, n24170, n24171, n24173, n24174,
         n24175, n24180, n24181, n24182, n24183, n24184, n24185, n24190,
         n24191, n24192, n24193, n24194, n24195, n24200, n24201, n24202,
         n24203, n24204, n24205, n24210, n24211, n24212, n24213, n24214,
         n24215, n24220, n24221, n24222, n24223, n24224, n24225, n24230,
         n24231, n24232, n24233, n24234, n24235, n24240, n24241, n24242,
         n24243, n24244, n24245, n24250, n24251, n24252, n24253, n24254,
         n24255, n24260, n24261, n24262, n24263, n24264, n24265, n24270,
         n24271, n24272, n24273, n24274, n24275, n24280, n24281, n24282,
         n24283, n24284, n24285, n24290, n24291, n24292, n24293, n24294,
         n24295, n24300, n24301, n24302, n24303, n24304, n24305, n24310,
         n24311, n24312, n24313, n24314, n24315, n24320, n24321, n24322,
         n24323, n24324, n24325, n24330, n24331, n24332, n24333, n24334,
         n24335, n24340, n24341, n24342, n24343, n24344, n24345, n24350,
         n24351, n24352, n24353, n24354, n24355, n24360, n24361, n24362,
         n24363, n24364, n24365, n24370, n24371, n24372, n24373, n24374,
         n24375, n24376, n24377, n24382, n24383, n24384, n24385, n24386,
         n24387, n24392, n24393, n24394, n24395, n24396, n24397, n24402,
         n24403, n24404, n24405, n24406, n24407, n24412, n24413, n24414,
         n24415, n24416, n24417, n24422, n24423, n24424, n24425, n24426,
         n24427, n24432, n24433, n24434, n24435, n24436, n24437, n24442,
         n24443, n24444, n24445, n24446, n24447, n24452, n24453, n24454,
         n24455, n24456, n24457, n24462, n24463, n24464, n24465, n24466,
         n24467, n24472, n24473, n24474, n24475, n24476, n24477, n24482,
         n24483, n24484, n24485, n24486, n24487, n24492, n24493, n24494,
         n24495, n24496, n24497, n24502, n24503, n24504, n24505, n24506,
         n24507, n24512, n24513, n24514, n24515, n24516, n24517, n24522,
         n24523, n24524, n24525, n24526, n24527, n24532, n24533, n24534,
         n24535, n24536, n24537, n24542, n24543, n24544, n24545, n24546,
         n24548, n24553, n24554, n24555, n24556, n24557, n24559, n24564,
         n24565, n24566, n24567, n24568, n24569, n24574, n24575, n24576,
         n24577, n24578, n24579, n24584, n24585, n24586, n24587, n24588,
         n24589, n24594, n24595, n24596, n24597, n24598, n24599, n24604,
         n24605, n24606, n24607, n24608, n24609, n24614, n24615, n24616,
         n24617, n24618, n24619, n24624, n24625, n24626, n24627, n24628,
         n24629, n24634, n24635, n24636, n24637, n24638, n24640, n24645,
         n24646, n24647, n24648, n24649, n24651, n24656, n24657, n24658,
         n24659, n24660, n24661, n24665, n24667, n24670, n24671, n24672,
         n24675, n24678, n24680, n24683, n24684, n24685, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24711, n24712,
         n24717, n24718, n24722, n24732, n24733, n24734, n24735, n24736,
         n24737, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
         n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756,
         n24757, n24762, n24763, n24764, n24765, n24766, n24767, n24772,
         n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780,
         n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24792,
         n24793, n24794, n24795, n24796, n24797, n24802, n24803, n24804,
         n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812,
         n24813, n24814, n24815, n24816, n24817, n24822, n24823, n24824,
         n24825, n24826, n24827, n24832, n24833, n24834, n24835, n24836,
         n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
         n24845, n24846, n24847, n24852, n24853, n24854, n24855, n24856,
         n24857, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
         n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
         n24877, n24882, n24883, n24884, n24885, n24886, n24887, n24892,
         n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900,
         n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24912,
         n24913, n24914, n24915, n24916, n24917, n24922, n24923, n24924,
         n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932,
         n24933, n24934, n24935, n24936, n24937, n24942, n24943, n24944,
         n24945, n24946, n24947, n24952, n24953, n24954, n24955, n24956,
         n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
         n24965, n24966, n24967, n24972, n24973, n24974, n24977, n24982,
         n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990,
         n24991, n24992, n24993, n24994, n24995, n24996, n24997, n25002,
         n25003, n25004, n25005, n25006, n25007, n25012, n25013, n25014,
         n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022,
         n25023, n25024, n25025, n25026, n25027, n25032, n25033, n25034,
         n25035, n25036, n25037, n25042, n25043, n25044, n25045, n25046,
         n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054,
         n25055, n25056, n25057, n25062, n25063, n25064, n25065, n25066,
         n25067, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
         n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086,
         n25087, n25092, n25093, n25094, n25095, n25096, n25097, n25102,
         n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110,
         n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25122,
         n25123, n25124, n25125, n25126, n25127, n25132, n25133, n25134,
         n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142,
         n25143, n25144, n25145, n25146, n25147, n25152, n25153, n25154,
         n25155, n25156, n25157, n25162, n25163, n25164, n25165, n25166,
         n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174,
         n25175, n25176, n25177, n25182, n25183, n25184, n25185, n25186,
         n25187, n25192, n25193, n25194, n25195, n25196, n25197, n25198,
         n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206,
         n25207, n25693, n25694, n25695, n25696, n25697, n25698, n25703,
         n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711,
         n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25723,
         n25724, n25725, n25726, n25727, n25728, n25733, n25734, n25735,
         n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
         n25744, n25745, n25746, n25747, n25748, n25753, n25754, n25755,
         n25756, n25757, n25758, n25763, n25764, n25765, n25766, n25767,
         n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
         n25776, n25777, n25778, n25783, n25784, n25785, n25786, n25787,
         n25788, n25793, n25794, n25795, n25796, n25797, n25798, n25799,
         n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807,
         n25808, n25813, n25814, n25815, n25816, n25817, n25818, n25823,
         n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831,
         n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25843,
         n25844, n25845, n25846, n25847, n25848, n25853, n25854, n25855,
         n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
         n25864, n25865, n25866, n25867, n25868, n25873, n25874, n25875,
         n25876, n25877, n25878, n25883, n25884, n25885, n25886, n25887,
         n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895,
         n25896, n25897, n25898, n25903, n25904, n25905, n25906, n25907,
         n25908, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
         n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927,
         n25928, n25933, n25934, n25935, n25936, n25937, n25938, n25943,
         n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
         n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25963,
         n25964, n25965, n25966, n25967, n25968, n25973, n25974, n25975,
         n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983,
         n25984, n25985, n25986, n25987, n25988, n25993, n25994, n25995,
         n25996, n25997, n25998, n26003, n26004, n26005, n26006, n26007,
         n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015,
         n26016, n26017, n26018, n26023, n26024, n26025, n26026, n26027,
         n26028, n26033, n26034, n26035, n26036, n26037, n26038, n26039,
         n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047,
         n26048, n26053, n26054, n26055, n26056, n26057, n26058, n26063,
         n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
         n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26083,
         n26084, n26085, n26086, n26087, n26088, n26093, n26094, n26095,
         n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
         n26104, n26105, n26106, n26107, n26108, n26113, n26114, n26115,
         n26116, n26117, n26118, n26123, n26124, n26125, n26126, n26127,
         n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
         n26136, n26137, n26138, n26143, n26144, n26145, n26146, n26147,
         n26148, n26153, n26154, n26155, n26156, n26157, n26158, n26159,
         n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
         n26168, n26173, n26174, n26175, n26176, n26177, n26178, n26183,
         n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191,
         n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26203,
         n26204, n26205, n26206, n26207, n26208, n26213, n26214, n26215,
         n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223,
         n26224, n26225, n26226, n26227, n26228, n26233, n26234, n26235,
         n26236, n26237, n26238, n26243, n26244, n26245, n26246, n26247,
         n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255,
         n26256, n26257, n26258, n26263, n26264, n26265, n26266, n26267,
         n26268, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
         n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287,
         n26288, n26293, n26294, n26295, n26296, n26297, n26298, n26303,
         n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311,
         n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26323,
         n26324, n26325, n26326, n26327, n26328, n26333, n26334, n26335,
         n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
         n26344, n26345, n26346, n26347, n26348, n26353, n26354, n26355,
         n26356, n26357, n26358, n26363, n26364, n26365, n26366, n26367,
         n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
         n26376, n26377, n26378, n26383, n26384, n26385, n26386, n26387,
         n26388, n26393, n26394, n26395, n26396, n26397, n26398, n26399,
         n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
         n26408, n26409, n26414, n26415, n26416, n26417, n26418, n26419,
         n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
         n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439,
         n26444, n26445, n26446, n26447, n26448, n26449, n26454, n26455,
         n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
         n26464, n26465, n26466, n26467, n26468, n26469, n26474, n26475,
         n26476, n26477, n26478, n26479, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26504, n26505, n26506, n26507,
         n26508, n26509, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26534, n26535, n26536, n26537, n26538, n26539,
         n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
         n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
         n26564, n26565, n26566, n26567, n26568, n26569, n26574, n26575,
         n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583,
         n26584, n26585, n26586, n26587, n26588, n26589, n26594, n26595,
         n26596, n26597, n26598, n26599, n26604, n26605, n26606, n26607,
         n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
         n26616, n26617, n26618, n26619, n26624, n26625, n26626, n26627,
         n26628, n26629, n26634, n26635, n26636, n26637, n26638, n26639,
         n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
         n26648, n26649, n26650, n26655, n26656, n26657, n26658, n26659,
         n26660, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
         n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
         n26680, n26685, n26686, n26687, n26688, n26689, n26690, n26695,
         n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703,
         n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26715,
         n26716, n26717, n26718, n26719, n26720, n26725, n26726, n26727,
         n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735,
         n26736, n26737, n26738, n26739, n26740, n26745, n26746, n26747,
         n26749, n26750, n26755, n26756, n26757, n26758, n26759, n26760,
         n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,
         n26769, n26770, n26775, n26776, n26777, n26778, n26779, n26780,
         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
         n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,
         n26805, n26806, n26807, n26808, n26809, n26810, n26815, n26816,
         n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
         n26825, n26826, n26827, n26828, n26829, n26830, n26835, n26836,
         n26837, n26838, n26839, n26840, n26845, n26846, n26847, n26848,
         n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
         n26857, n26858, n26859, n26860, n26865, n26866, n26867, n26868,
         n26869, n26870, n26875, n26876, n26877, n26878, n26879, n26880,
         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
         n26889, n26890, n26891, n26896, n26897, n26898, n26899, n26900,
         n26901, n26906, n26907, n26908, n26909, n26910, n26911, n26912,
         n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
         n26921, n26926, n26927, n26928, n26929, n26930, n26931, n26936,
         n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,
         n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26956,
         n26957, n26958, n26959, n26960, n26961, n26966, n26967, n26968,
         n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976,
         n26977, n26978, n26979, n26980, n26981, n26986, n26987, n26988,
         n26989, n26990, n26991, n26996, n26997, n26998, n26999, n27000,
         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
         n27009, n27010, n27011, n27016, n27017, n27018, n27019, n27020,
         n27021, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
         n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
         n27041, n27046, n27047, n27048, n27049, n27050, n27051, n27056,
         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
         n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27076,
         n27077, n27078, n27079, n27080, n27081, n27086, n27087, n27088,
         n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,
         n27097, n27098, n27099, n27100, n27101, n27106, n27107, n27108,
         n27109, n27110, n27111, n27116, n27117, n27118, n27119, n27120,
         n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
         n27129, n27130, n27131, n27132, n27137, n27138, n27139, n27140,
         n27141, n27142, n27147, n27148, n27149, n27150, n27151, n27152,
         n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
         n27161, n27162, n27167, n27168, n27169, n27170, n27171, n27172,
         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
         n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192,
         n27197, n27198, n27199, n27200, n27201, n27202, n27207, n27208,
         n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,
         n27217, n27218, n27219, n27220, n27221, n27222, n27227, n27228,
         n27229, n27230, n27231, n27232, n27237, n27238, n27239, n27240,
         n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
         n27249, n27250, n27251, n27252, n27257, n27258, n27259, n27260,
         n27261, n27262, n27267, n27268, n27269, n27270, n27271, n27272,
         n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,
         n27281, n27282, n27287, n27288, n27289, n27290, n27291, n27292,
         n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
         n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,
         n27317, n27318, n27319, n27320, n27321, n27322, n27327, n27328,
         n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,
         n27337, n27338, n27339, n27340, n27341, n27342, n27347, n27348,
         n27349, n27350, n27351, n27352, n27357, n27358, n27359, n27360,
         n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
         n27369, n27370, n27371, n27372, n27373, n27378, n27379, n27380,
         n27381, n27382, n27383, n27388, n27389, n27390, n27391, n27392,
         n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,
         n27401, n27402, n27403, n27408, n27409, n27410, n27411, n27412,
         n27413, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
         n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
         n27433, n27438, n27439, n27440, n27443, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27468, n27469, n27470,
         n27473, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
         n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492,
         n27493, n27498, n27499, n27500, n27501, n27502, n27503, n27508,
         n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516,
         n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27528,
         n27529, n27530, n27531, n27532, n27533, n27538, n27539, n27540,
         n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548,
         n27549, n27550, n27551, n27552, n27553, n27558, n27559, n27560,
         n27561, n27562, n27563, n27568, n27569, n27570, n27571, n27572,
         n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580,
         n27581, n27582, n27583, n27588, n27589, n27590, n27591, n27592,
         n27593, n27598, n27599, n27600, n27601, n27602, n27603, n27604,
         n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612,
         n27613, n27614, n27679, n27680, n27681, n27682, n27683, n27684,
         n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696,
         n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704,
         n27709, n27710, n27711, n27712, n27713, n27714, n27719, n27720,
         n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27730,
         n27731, n27732, n27734, n27979, n27980, n27981, n27982, n27983,
         n27984, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28009, n28010, n28011, n28012, n28013, n28014, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28039,
         n28040, n28041, n28042, n28043, n28044, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28069, n28070, n28071,
         n28072, n28073, n28074, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28100, n28101, n28102, n28103,
         n28104, n28105, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28130, n28131, n28132, n28133, n28134, n28135,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28160, n28161, n28162, n28163, n28164, n28165, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28190, n28191,
         n28192, n28193, n28194, n28195, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28220, n28221, n28222, n28223,
         n28224, n28225, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28250, n28251, n28252, n28253, n28254, n28255,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28280, n28281, n28282, n28283, n28284, n28285, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28310, n28311,
         n28312, n28313, n28314, n28315, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28340, n28341, n28342, n28343,
         n28344, n28345, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28370, n28371, n28372, n28373, n28374, n28375,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28400, n28401, n28402, n28403, n28404, n28405, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28430, n28431,
         n28432, n28433, n28434, n28435, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28460, n28461, n28462, n28463,
         n28464, n28465, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28490, n28491, n28492, n28493, n28494, n28495,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28520, n28521, n28522, n28523, n28524, n28525, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28550, n28551,
         n28552, n28553, n28554, n28555, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n29001, n29002, n29003, n29004,
         n29005, n29006, n29011, n29012, n29013, n29014, n29015, n29016,
         n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024,
         n29025, n29026, n29031, n29032, n29033, n29034, n29035, n29036,
         n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048,
         n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056,
         n29061, n29062, n29063, n29064, n29065, n29066, n29071, n29072,
         n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
         n29081, n29082, n29083, n29084, n29085, n29086, n29091, n29092,
         n29093, n29094, n29095, n29096, n29101, n29102, n29103, n29104,
         n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112,
         n29113, n29114, n29115, n29116, n29117, n29122, n29123, n29124,
         n29126, n29127, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29152, n29153, n29154, n29156, n29157, n29162,
         n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
         n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29182,
         n29183, n29184, n29185, n29186, n29187, n29192, n29193, n29194,
         n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202,
         n29203, n29204, n29205, n29206, n29207, n29212, n29213, n29214,
         n29215, n29216, n29217, n29222, n29223, n29224, n29225, n29226,
         n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234,
         n29235, n29236, n29237, n29242, n29243, n29244, n29245, n29246,
         n29247, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
         n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266,
         n29267, n29272, n29273, n29274, n29275, n29276, n29277, n29282,
         n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290,
         n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29302,
         n29303, n29304, n29305, n29306, n29307, n29312, n29313, n29314,
         n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322,
         n29323, n29324, n29325, n29326, n29327, n29332, n29333, n29334,
         n29335, n29336, n29337, n29342, n29343, n29344, n29345, n29346,
         n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354,
         n29355, n29356, n29357, n29362, n29363, n29364, n29365, n29366,
         n29367, n29372, n29373, n29374, n29375, n29376, n29377, n29378,
         n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
         n29387, n29392, n29393, n29394, n29395, n29396, n29397, n29402,
         n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29422,
         n29423, n29424, n29425, n29426, n29427, n29432, n29433, n29434,
         n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442,
         n29443, n29444, n29445, n29446, n29447, n29452, n29453, n29454,
         n29455, n29456, n29457, n29462, n29463, n29464, n29465, n29466,
         n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
         n29475, n29476, n29477, n29478, n29483, n29484, n29485, n29486,
         n29487, n29488, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29507, n29508, n29513, n29514, n29515, n29516, n29517, n29518,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538,
         n29543, n29544, n29545, n29546, n29547, n29548, n29553, n29554,
         n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562,
         n29563, n29564, n29565, n29566, n29567, n29568, n29573, n29574,
         n29575, n29576, n29577, n29578, n29583, n29584, n29585, n29586,
         n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594,
         n29595, n29596, n29597, n29598, n29603, n29604, n29605, n29606,
         n29607, n29608, n29613, n29614, n29615, n29616, n29617, n29618,
         n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
         n29627, n29628, n29633, n29634, n29635, n29636, n29637, n29638,
         n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
         n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
         n29663, n29664, n29665, n29666, n29667, n29668, n29673, n29674,
         n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682,
         n29683, n29684, n29685, n29686, n29687, n29688, n29693, n29694,
         n29695, n29696, n29697, n29698, n29703, n29704, n29705, n29706,
         n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
         n29715, n29716, n29717, n29718, n29719, n29724, n29725, n29726,
         n29727, n29728, n29729, n29734, n29735, n29736, n29737, n29738,
         n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
         n29747, n29748, n29749, n29754, n29755, n29756, n29757, n29758,
         n29759, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
         n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778,
         n29779, n29784, n29785, n29786, n29787, n29788, n29789, n29794,
         n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802,
         n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29814,
         n29815, n29816, n29817, n29818, n29819, n29824, n29825, n29826,
         n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
         n29835, n29836, n29837, n29838, n29839, n29844, n29845, n29846,
         n29847, n29848, n29849, n29854, n29855, n29856, n29857, n29858,
         n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866,
         n29867, n29868, n29869, n29874, n29875, n29876, n29877, n29878,
         n29879, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
         n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898,
         n29899, n29904, n29905, n29906, n29907, n29908, n29909, n29914,
         n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922,
         n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29934,
         n29935, n29936, n29937, n29938, n29939, n29944, n29945, n29946,
         n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954,
         n29955, n29956, n29957, n29958, n29959, n29964, n29965, n29966,
         n29967, n29968, n29969, n29974, n29975, n29976, n29977, n29978,
         n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986,
         n29987, n29988, n29989, n29994, n29995, n29996, n29997, n29998,
         n29999, n30004, n30005, n30006, n30007, n30008, n30009, n30010,
         n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018,
         n30019, n30024, n30025, n30026, n30027, n30028, n30029, n30034,
         n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042,
         n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30054,
         n30055, n30056, n30057, n30058, n30059, n30064, n30065, n30066,
         n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074,
         n30075, n30076, n30077, n30078, n30079, n30084, n30085, n30086,
         n30087, n30088, n30089, n30094, n30095, n30096, n30097, n30098,
         n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
         n30107, n30108, n30109, n30114, n30115, n30116, n30117, n30118,
         n30119, n30124, n30125, n30126, n30127, n30128, n30129, n30130,
         n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138,
         n30139, n30144, n30145, n30146, n30147, n30148, n30149, n30154,
         n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162,
         n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30174,
         n30175, n30176, n30177, n30178, n30179, n30184, n30185, n30186,
         n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194,
         n30195, n30196, n30197, n30198, n30199, n30200, n30205, n30206,
         n30207, n30208, n30209, n30210, n30215, n30216, n30217, n30218,
         n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226,
         n30227, n30228, n30229, n30230, n30235, n30236, n30237, n30238,
         n30239, n30240, n30245, n30246, n30247, n30248, n30249, n30250,
         n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258,
         n30259, n30260, n30265, n30266, n30267, n30268, n30269, n30270,
         n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282,
         n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290,
         n30295, n30296, n30297, n30298, n30299, n30300, n30305, n30306,
         n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314,
         n30315, n30316, n30317, n30318, n30319, n30320, n30325, n30326,
         n30327, n30328, n30329, n30330, n30335, n30336, n30337, n30338,
         n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346,
         n30347, n30348, n30349, n30350, n30355, n30356, n30357, n30358,
         n30359, n30360, n30365, n30366, n30367, n30368, n30369, n30370,
         n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378,
         n30379, n30380, n30385, n30386, n30387, n30388, n30389, n30390,
         n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402,
         n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410,
         n30415, n30416, n30417, n30418, n30419, n30420, n30425, n30426,
         n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434,
         n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442,
         n30447, n30448, n30449, n30450, n30451, n30452, n30457, n30458,
         n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466,
         n30467, n30468, n30469, n30470, n30471, n30472, n30477, n30478,
         n30479, n30480, n30481, n30482, n30487, n30488, n30489, n30490,
         n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498,
         n30499, n30500, n30501, n30502, n30507, n30508, n30509, n30510,
         n30511, n30512, n30517, n30518, n30519, n30520, n30521, n30522,
         n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530,
         n30531, n30532, n30537, n30538, n30539, n30540, n30541, n30542,
         n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554,
         n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562,
         n30567, n30568, n30569, n30570, n30571, n30572, n30577, n30578,
         n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586,
         n30587, n30588, n30589, n30590, n30591, n30592, n30597, n30598,
         n30599, n30600, n30601, n30602, n30607, n30608, n30609, n30610,
         n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618,
         n30619, n30620, n30621, n30622, n30627, n30628, n30629, n30630,
         n30631, n30632, n30637, n30638, n30639, n30640, n30641, n30642,
         n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650,
         n30651, n30652, n30657, n30658, n30659, n30660, n30661, n30662,
         n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674,
         n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
         n30683, n30688, n30689, n30690, n30691, n30692, n30693, n30698,
         n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706,
         n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30718,
         n30719, n30720, n30721, n30722, n30723, n30728, n30729, n30730,
         n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738,
         n30739, n30740, n30741, n30742, n30743, n30748, n30749, n30750,
         n30751, n30752, n30753, n30758, n30759, n30760, n30761, n30762,
         n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
         n30771, n30772, n30773, n30778, n30779, n30780, n30781, n30782,
         n30783, n30788, n30789, n30790, n30791, n30792, n30793, n30794,
         n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802,
         n30803, n30808, n30809, n30810, n30811, n30812, n30813, n30818,
         n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826,
         n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30838,
         n30839, n30840, n30841, n30842, n30843, n30848, n30849, n30850,
         n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858,
         n30859, n30860, n30861, n30862, n30863, n30868, n30869, n30870,
         n30871, n30872, n30873, n30878, n30879, n30880, n30881, n30882,
         n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890,
         n30891, n30892, n30893, n30898, n30899, n30900, n30901, n30902,
         n30903, n30908, n30909, n30910, n30911, n30912, n30913, n30914,
         n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922,
         n30923, n30928, n30929, n30930, n30931, n30932, n30933, n30938,
         n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946,
         n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30958,
         n30959, n30960, n30961, n30962, n30963, n30968, n30969, n30970,
         n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978,
         n30979, n30980, n30981, n30982, n30983, n30988, n30989, n30990,
         n30991, n30992, n30993, n30998, n30999, n31000, n31001, n31002,
         n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010,
         n31011, n31012, n31013, n31018, n31019, n31020, n31021, n31022,
         n31023, n31028, n31029, n31030, n31031, n31032, n31033, n31034,
         n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042,
         n31043, n31048, n31049, n31050, n31051, n31052, n31053, n31058,
         n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066,
         n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31078,
         n31079, n31080, n31081, n31082, n31083, n31088, n31089, n31090,
         n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098,
         n31099, n31100, n31101, n31102, n31103, n31108, n31109, n31110,
         n31111, n31112, n31113, n31118, n31119, n31120, n31121, n31122,
         n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130,
         n31131, n31132, n31133, n31138, n31139, n31140, n31141, n31142,
         n31143, n31148, n31149, n31150, n31151, n31152, n31153, n31154,
         n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162,
         n31163, n31164, n31169, n31170, n31171, n31172, n31173, n31174,
         n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186,
         n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194,
         n31199, n31200, n31201, n31202, n31203, n31204, n31209, n31210,
         n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218,
         n31219, n31220, n31221, n31222, n31223, n31224, n31229, n31230,
         n31231, n31232, n31233, n31234, n31239, n31240, n31241, n31242,
         n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250,
         n31251, n31252, n31253, n31254, n31259, n31260, n31261, n31262,
         n31263, n31264, n31269, n31270, n31271, n31272, n31273, n31274,
         n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282,
         n31283, n31284, n31289, n31290, n31291, n31292, n31293, n31294,
         n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306,
         n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314,
         n31319, n31320, n31321, n31322, n31323, n31324, n31329, n31330,
         n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338,
         n31339, n31340, n31341, n31342, n31343, n31344, n31349, n31350,
         n31351, n31352, n31353, n31354, n31359, n31360, n31361, n31362,
         n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370,
         n31371, n31372, n31373, n31374, n31379, n31380, n31381, n31382,
         n31383, n31384, n31389, n31390, n31391, n31392, n31393, n31394,
         n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402,
         n31403, n31404, n31409, n31410, n31411, n31412, n31413, n31414,
         n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426,
         n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434,
         n31439, n31440, n31441, n31442, n31443, n31444, n31449, n31450,
         n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458,
         n31459, n31460, n31461, n31462, n31463, n31464, n31469, n31470,
         n31471, n31472, n31473, n31474, n31479, n31480, n31481, n31482,
         n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
         n31491, n31492, n31493, n31494, n31499, n31500, n31501, n31502,
         n31503, n31504, n31509, n31510, n31511, n31512, n31513, n31514,
         n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522,
         n31523, n31524, n31529, n31530, n31531, n31532, n31533, n31534,
         n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546,
         n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554,
         n31559, n31560, n31561, n31562, n31563, n31564, n31569, n31570,
         n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578,
         n31579, n31580, n31581, n31582, n31583, n31584, n31589, n31590,
         n31591, n31592, n31593, n31594, n31599, n31600, n31601, n31602,
         n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610,
         n31611, n31612, n31613, n31614, n31619, n31620, n31621, n31622,
         n31623, n31624, n31629, n31630, n31631, n31632, n31633, n31634,
         n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642,
         n31643, n31644, n31645, n31650, n31651, n31652, n31653, n31654,
         n31655, n31660, n31661, n31662, n31663, n31664, n31665, n31666,
         n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674,
         n31675, n31680, n31681, n31682, n31683, n31684, n31685, n31690,
         n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698,
         n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31710,
         n31711, n31712, n31713, n31714, n31715, n31720, n31721, n31722,
         n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730,
         n31731, n31732, n31733, n31734, n31735, n31740, n31741, n31742,
         n31743, n31744, n31745, n31750, n31751, n31752, n31753, n31754,
         n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762,
         n31763, n31764, n31765, n31770, n31771, n31772, n31773, n31774,
         n31775, n31780, n31781, n31782, n31783, n31784, n31785, n31786,
         n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794,
         n31795, n31800, n31801, n31802, n31803, n31804, n31805, n31810,
         n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818,
         n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31830,
         n31831, n31832, n31833, n31834, n31835, n31840, n31841, n31842,
         n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850,
         n31851, n31852, n31853, n31854, n31855, n31860, n31861, n31862,
         n31863, n31864, n31865, n31870, n31871, n31872, n31873, n31874,
         n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882,
         n31883, n31884, n31885, n31886, n31891, n31892, n31893, n31894,
         n31895, n31896, n31901, n31902, n31903, n31904, n31905, n31906,
         n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914,
         n31915, n31916, n31921, n31922, n31923, n31924, n31925, n31926,
         n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938,
         n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946,
         n31951, n31952, n31953, n31954, n31955, n31956, n31961, n31962,
         n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970,
         n31971, n31972, n31973, n31974, n31975, n31976, n31981, n31982,
         n31983, n31984, n31985, n31986, n31991, n31992, n31993, n31994,
         n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002,
         n32003, n32004, n32005, n32006, n32011, n32012, n32013, n32014,
         n32015, n32016, n32021, n32022, n32023, n32024, n32025, n32026,
         n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034,
         n32035, n32036, n32041, n32042, n32043, n32044, n32045, n32046,
         n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058,
         n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066,
         n32071, n32072, n32073, n32074, n32075, n32076, n32081, n32082,
         n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090,
         n32091, n32092, n32093, n32094, n32095, n32096, n32101, n32102,
         n32103, n32104, n32105, n32106, n32111, n32112, n32113, n32114,
         n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
         n32123, n32124, n32125, n32126, n32131, n32132, n32133, n32134,
         n32135, n32136, n32141, n32142, n32143, n32144, n32145, n32146,
         n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154,
         n32155, n32156, n32161, n32162, n32163, n32164, n32165, n32166,
         n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178,
         n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186,
         n32191, n32192, n32193, n32194, n32195, n32196, n32201, n32202,
         n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
         n32211, n32212, n32213, n32214, n32215, n32216, n32221, n32222,
         n32223, n32224, n32225, n32226, n32231, n32232, n32233, n32234,
         n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242,
         n32243, n32244, n32245, n32246, n32251, n32252, n32253, n32254,
         n32255, n32256, n32261, n32262, n32263, n32264, n32265, n32266,
         n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274,
         n32275, n32276, n32281, n32282, n32283, n32284, n32285, n32286,
         n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298,
         n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306,
         n32311, n32312, n32313, n32314, n32315, n32316, n32321, n32322,
         n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330,
         n32331, n32332, n32333, n32334, n32335, n32336, n32341, n32342,
         n32343, n32344, n32345, n32346, n32351, n32352, n32353, n32354,
         n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
         n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370,
         n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391,
         n32392, n32393, n32394, n32395, n32397, n32398, n32399, n32400,
         n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408,
         n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416,
         n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424,
         n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432,
         n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440,
         n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448,
         n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456,
         n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464,
         n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472,
         n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480,
         n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488,
         n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496,
         n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504,
         n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512,
         n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520,
         n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528,
         n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536,
         n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544,
         n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552,
         n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560,
         n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568,
         n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576,
         n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584,
         n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592,
         n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600,
         n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608,
         n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616,
         n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624,
         n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632,
         n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640,
         n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648,
         n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656,
         n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664,
         n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672,
         n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680,
         n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688,
         n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696,
         n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704,
         n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712,
         n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720,
         n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728,
         n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736,
         n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744,
         n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752,
         n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760,
         n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768,
         n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776,
         n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784,
         n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792,
         n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800,
         n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808,
         n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816,
         n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824,
         n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832,
         n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840,
         n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848,
         n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856,
         n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864,
         n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872,
         n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880,
         n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888,
         n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896,
         n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904,
         n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912,
         n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920,
         n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928,
         n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936,
         n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944,
         n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952,
         n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960,
         n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968,
         n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976,
         n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984,
         n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992,
         n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000,
         n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008,
         n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016,
         n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024,
         n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032,
         n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040,
         n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048,
         n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056,
         n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064,
         n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072,
         n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080,
         n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088,
         n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096,
         n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104,
         n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112,
         n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120,
         n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128,
         n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136,
         n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144,
         n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152,
         n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160,
         n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168,
         n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176,
         n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184,
         n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192,
         n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200,
         n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208,
         n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216,
         n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224,
         n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232,
         n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240,
         n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248,
         n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
         n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264,
         n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272,
         n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280,
         n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288,
         n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296,
         n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304,
         n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312,
         n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320,
         n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328,
         n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336,
         n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344,
         n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352,
         n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360,
         n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368,
         n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376,
         n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384,
         n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392,
         n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400,
         n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408,
         n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416,
         n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424,
         n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432,
         n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440,
         n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448,
         n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456,
         n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464,
         n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472,
         n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480,
         n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488,
         n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496,
         n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504,
         n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512,
         n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520,
         n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528,
         n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536,
         n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544,
         n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552,
         n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560,
         n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568,
         n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576,
         n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584,
         n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592,
         n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600,
         n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608,
         n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616,
         n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624,
         n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632,
         n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640,
         n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648,
         n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656,
         n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664,
         n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672,
         n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680,
         n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688,
         n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696,
         n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704,
         n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712,
         n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720,
         n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728,
         n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736,
         n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744,
         n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752,
         n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760,
         n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768,
         n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776,
         n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784,
         n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792,
         n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800,
         n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808,
         n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816,
         n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824,
         n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832,
         n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840,
         n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848,
         n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856,
         n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864,
         n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872,
         n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880,
         n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888,
         n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896,
         n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904,
         n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912,
         n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920,
         n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928,
         n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936,
         n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944,
         n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952,
         n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960,
         n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968,
         n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976,
         n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984,
         n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992,
         n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000,
         n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008,
         n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016,
         n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024,
         n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032,
         n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040,
         n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048,
         n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056,
         n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064,
         n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072,
         n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080,
         n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088,
         n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096,
         n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104,
         n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112,
         n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120,
         n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128,
         n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136,
         n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144,
         n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152,
         n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160,
         n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168,
         n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176,
         n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184,
         n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192,
         n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200,
         n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208,
         n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216,
         n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224,
         n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232,
         n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240,
         n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248,
         n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256,
         n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264,
         n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272,
         n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280,
         n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288,
         n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296,
         n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304,
         n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312,
         n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320,
         n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328,
         n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336,
         n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344,
         n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352,
         n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360,
         n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368,
         n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376,
         n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384,
         n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392,
         n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400,
         n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408,
         n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416,
         n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424,
         n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432,
         n34435, n34436, n34437, n34438, n34439, n34441, n34442, n34443,
         n34444, n34445, n34447, n34448, n34449, n34450, n34451, n34452,
         n34453, n34454, n34455, n34456, n34457, n34458, n34460, n34461,
         n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472,
         n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480,
         n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488,
         n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496,
         n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504,
         n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512,
         n34513, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, net151225, net151243, net151246,
         net151248, net151249, net151251, net151253, net151258, net151261,
         net151263, net151264, net151265, net151266, net151270, net151271,
         net151275, net151279, net151283, net151299, net151304, net151308,
         net151325, net151327, net151330, net151333, net151340, net151347,
         net151348, net151349, net151356, net151373, net151374, net151380,
         net151394, net151401, net151404, net151420, net151426, net151430,
         net151431, net151435, net151440, net151443, net151444, net151445,
         net151448, net151451, net151452, net151453, net151456, net151458,
         net151462, net151465, net151467, net151473, net151477, net151479,
         net151481, net151491, net151494, net151495, net151503, net151504,
         net151509, net151514, net151530, net151532, net151536, net151539,
         net151541, net151542, net151550, net151554, net151555, net151557,
         net151558, net151562, net151566, net151571, net151584, net151586,
         net151587, net151593, net151594, net151599, net151600, net151601,
         net151612, net151644, net151652, net151653, net151662, net151666,
         net151670, net151672, net151673, net151705, net151708, net151711,
         net151712, net151720, net151721, net151723, net151726, net151728,
         net151733, net151737, net151738, net151741, net151744, net151746,
         net151750, net151751, net151753, net151757, net151758, net151766,
         net151767, net151769, net151772, net151773, net151775, net151779,
         net151785, net151786, net151788, net151789, net151790, net151793,
         net151806, net151809, net151812, net151819, net151847, net151848,
         net151857, net151860, net152412, net168842, net168843, net168846,
         net168848, net168849, net168850, net168852, net171098, net171099,
         net171101, net171103, net171104, net171105, net171108, net171111,
         net171113, net171114, net171117, net171119, net171122, net171124,
         net171125, net171126, net171127, net171129, net171132, net171134,
         net171136, net171139, net171140, net171142, net171143, net171145,
         net171146, net171148, net171151, net171152, net171153, net171156,
         net171158, net171160, net171168, net171169, net171175, net171178,
         net171180, net171182, net171183, net171185, net171188, net171189,
         net171191, net171192, net171196, net171198, net171199, net171200,
         net171201, net171205, net171207, net171210, net171211, net171214,
         net171218, net171222, net171231, net171233, net171234, net171236,
         net171237, net171238, net171240, net171242, net171245, net171247,
         net171248, net171249, net171252, net171255, net171257, net171259,
         net171262, net171264, net171270, net171272, net171274, net171278,
         net171280, net171283, net171288, net171290, net171294, net171297,
         net171300, net171301, net171304, net171305, net171307, net171309,
         net171313, net171314, net171315, net171318, net171319, net171321,
         net171327, net171328, net171349, net171380, net171386, net171388,
         net171390, net171392, net171394, net171396, net171398, net171401,
         net171403, net171406, net171408, net171412, net171414, net171416,
         net171417, net171418, net171421, net171423, net171425, net171427,
         net171430, net171433, net171435, net171437, net171439, net171440,
         net171441, net171443, net171445, net171447, net171448, net171449,
         net171453, net171456, net171458, net171459, net171460, net171461,
         net171462, net171467, net171469, net171470, net171471, net171472,
         net171474, net171476, net171477, net171478, net171480, net171482,
         net171483, net171486, net171489, net171490, net171491, net171523,
         net171524, net171525, net171528, net171530, net171532, net171533,
         net171534, net171535, net171537, net171538, net171540, net171542,
         net171544, net171545, net171546, net171547, net171548, net171550,
         net171551, net171554, net171555, net172112, net207642, net207653,
         net208565, net209087, net209099, net209101, net209103, net209111,
         net209124, net209136, net209142, net209144, net209145, net209151,
         net209155, net209158, net209161, net209165, net209171, net209172,
         net209175, net209176, net209179, net209182, net209185, net209197,
         net209202, net209203, net209210, net209211, net209225, net209228,
         net209231, net209234, net209242, net209249, net209250, net209253,
         net209254, net209255, net209258, net209259, net209267, net209268,
         net209277, net209280, net209283, net209284, net209287, net209288,
         net209289, net209290, net209291, net209296, net209298, net209300,
         net209301, net209302, net209303, net209307, net209308, net209310,
         net209311, net209312, net209313, net209314, net209315, net209316,
         net209317, net209320, net209323, net209325, net209333, net209335,
         net209341, net209342, net209343, net209344, net209347, net209350,
         net209355, net209362, net209367, net209372, net209395, net209402,
         net209441, net209446, net209455, net209463, net209466, net209469,
         net209476, net209479, net209482, net209483, net209486, net209503,
         net209504, net209507, net209509, net209513, net209516, net209517,
         net209519, net209520, net209528, net209529, net209537, net209543,
         net209546, net209547, net209549, net209557, net209565, net209570,
         net209572, net209582, net209583, net209584, net209589, net209591,
         net209592, net209595, net209602, net209603, net209604, net209605,
         net209606, net209615, net209617, net209620, net209622, net209623,
         net209624, net209627, net209628, net209629, net209631, net209633,
         net209634, net209635, net209636, net209638, net209642, net209659,
         net209661, net209663, net209664, net209669, net209675, net209676,
         net209689, net209697, net209701, net209732, net209733, net209736,
         net209739, net209746, net209749, net209750, net209753, net209760,
         net209763, net209764, net209767, net209768, net209769, net209772,
         net209773, net209778, net209781, net209784, net209787, net209791,
         net209800, net209814, net209817, net209821, net209840, net209844,
         net209846, net209862, net209868, net209873, net209884, net209885,
         net209893, net209894, net209898, net209899, net209900, net209901,
         net209902, net209903, net209919, net209923, net209924, net209926,
         net209927, net209930, net209944, net209953, net209956, net209958,
         net209960, net209964, net209969, net209971, net209974, net209976,
         net209977, net209992, net209996, net210007, net210034, net210043,
         net210047, net210057, net210058, net210067, net210075, net210078,
         net210081, net210089, net210091, net210099, net210100, net210109,
         net210132, net210140, net210142, net210148, net210205, net210207,
         net210209, net210210, net210211, net210213, net210216, net210221,
         net210222, net210233, net210234, net210238, net210239, net210242,
         net210251, net210254, net210255, net210258, net210259, net210348,
         net210350, net210353, net210356, net210363, net210366, net210368,
         net210371, net210390, net210392, net210416, net210417, net210424,
         net210426, net210434, net210435, net210441, net210442, net210443,
         net210444, net210445, net210460, net210462, net210469, net210473,
         net210475, net210476, net210477, net210479, net210481, net210490,
         net210492, net210494, net210497, net210499, net210507, net210510,
         net210512, net210516, net210517, net210520, net210522, net210523,
         net210524, net210525, net210526, net210528, net210531, net210536,
         net210537, net210539, net210543, net210544, net210548, net210550,
         net210552, net210553, net210554, net210555, net210556, net210557,
         net210559, net210561, net210567, net210579, net210580, net210581,
         net210582, net210583, net210584, net210585, net210587, net210596,
         net210597, net210598, net210599, net210601, net210615, net210616,
         net210617, net210618, net210620, net210621, net210623, net210635,
         net210639, net210641, net210643, net210646, net210650, net210659,
         net210660, net210665, net210667, net210668, net210669, net210670,
         net210673, net210675, net210677, net210680, net210682, net210688,
         net210690, net210695, net210698, net210699, net210702, net210704,
         net210705, net210749, net210770, net210771, net210772, net210848,
         net210919, net211102, net211147, net211150, net211152, net211155,
         net211167, net211170, net211182, net211184, net211187, net211188,
         net211189, net211190, net211197, net211246, net211247, net211248,
         net211249, net211251, net211252, net211253, net211254, net211256,
         net211257, net211258, net211259, net211261, net211262, net211263,
         net211264, net211271, net211348, net211351, net211433, net211435,
         net211438, net211439, net211440, net211441, net211443, net211444,
         net211445, net211446, net211448, net211450, net211453, net211456,
         net211458, net211461, net211463, net211466, net211468, net211469,
         net211470, net211471, net211473, net211474, net211475, net211476,
         net211478, net211479, net211480, net211481, net211483, net211485,
         net211488, net211489, net211490, net211491, net211508, net211511,
         net211513, net211516, net211518, net211521, net211523, net211526,
         net211558, net211559, net211560, net211561, net211563, net211565,
         net211568, net211574, net211576, net211579, net211580, net211581,
         net211582, net211584, net211585, net211588, net211590, net211591,
         net211594, net211597, net211600, net211602, net211603, net211606,
         net211608, net211611, net211613, net211614, net211615, net211616,
         net211618, net211619, net211620, net211621, net211623, net211626,
         net211629, net211630, net211631, net211635, net211637, net211640,
         net211641, net211642, net211643, net211644, net211651, net211652,
         net211653, net211654, net211656, net211657, net211658, net211659,
         net211660, net211667, net211768, net211770, net211773, net211775,
         net211778, net211780, net211783, net211785, net211788, net211790,
         net211793, net211794, net211795, net211796, net211957, net211959,
         net211962, net211965, net211967, net211968, net211969, net211970,
         net211972, net211973, net211974, net211975, net211982, net211984,
         net211987, net211990, net211992, net211993, net211994, net211995,
         net211997, net212000, net212002, net212005, net212017, net212020,
         net212022, net212023, net212024, net212025, net212027, net212030,
         net212037, net212038, net212041, net212043, net212044, net212045,
         net212046, net212048, net212049, net212050, net212051, net212053,
         net212055, net212058, net212059, net212060, net212061, net212063,
         net212065, net212068, net212069, net212070, net212071, net212073,
         net212074, net212075, net212076, net212078, net212079, net212080,
         net212081, net212088, net212089, net212090, net212091, net212092,
         net212094, net212096, net212099, net212101, net212104, net212105,
         net212106, net212107, net212114, net212115, net212116, net212117,
         net212119, net212120, net212121, net212122, net212124, net212125,
         net212126, net212129, net212130, net212131, net212132, net212134,
         net212135, net212136, net212137, net212144, net212145, net212146,
         net212147, net212154, net212155, net212156, net212157, net212159,
         net212160, net212161, net212162, net212164, net212165, net212166,
         net212169, net212170, net212171, net212172, net212174, net212175,
         net212176, net212177, net212184, net212185, net212186, net212187,
         net212189, net212190, net212192, net212194, net212195, net212196,
         net212212, net212213, net212214, net212238, net212262, net212374,
         net212377, net212385, net212386, net212387, net212388, net212463,
         net212466, net212474, net212475, net212476, net212552, net212553,
         net212554, net212555, net212557, net212558, net212559, net212560,
         net212562, net212565, net212567, net212569, net212570, net212642,
         net212643, net212664, net212691, net212694, net212711, net212714,
         net212716, net212719, net212726, net212729, net212731, net212734,
         net212736, net212739, net212741, net212744, net212826, net212829,
         net212831, net212834, net212836, net212839, net212846, net212849,
         net212851, net212854, net212856, net212859, net212861, net212864,
         net212866, net212869, net212871, net212874, net212896, net212899,
         net212901, net212904, net212906, net212909, net212911, net212912,
         net212913, net212981, net212982, net212983, net212984, net213016,
         net213017, net213021, net213022, net213023, net213115, net213116,
         net213125, net213126, net213190, net213191, net213192, net213193,
         net213195, net213196, net213197, net213198, net213200, net213201,
         net213202, net213203, net213205, net213206, net213207, net213208,
         net213210, net213211, net213212, net213213, net213215, net213216,
         net213217, net213218, net213220, net213221, net213222, net213223,
         net213225, net213226, net213227, net213228, net213230, net213231,
         net213232, net213233, net213234, net213236, net213239, net213312,
         net213315, net213317, net213320, net213342, net213345, net213347,
         net213350, net213352, net213353, net213354, net213355, net213357,
         net213360, net213362, net213363, net213364, net213365, net213402,
         net213405, net213422, net213423, net213447, net213450, net213462,
         net213464, net213467, net213469, net213472, net213473, net213474,
         net213475, net213477, net213480, net213487, net213490, net213497,
         net213500, net213502, net213505, net213507, net213510, net213512,
         net213515, net213517, net213520, net213522, net213525, net213527,
         net213530, net213532, net213535, net213537, net213540, net213542,
         net213545, net213552, net213555, net213557, net213560, net213562,
         net213565, net213567, net213570, net213572, net213575, net213582,
         net213585, net213587, net213590, net213592, net213595, net213597,
         net213598, net213599, net213602, net213603, net213606, net213608,
         net213611, net213613, net213616, net213618, net213621, net213623,
         net213626, net213633, net213636, net213653, net213659, net213660,
         net213661, net213666, net213675, net213678, net213679, net213680,
         net213687, net213700, net213701, net213702, net213703, net213731,
         net213732, net213733, net213734, net213824, net213901, net213902,
         net213950, net214016, net214154, net214265, net214389, net214390,
         net214391, net214392, net214433, net214435, net214515, net214641,
         net214643, net214644, net214646, net214649, net214662, net214663,
         net214669, net214672, net214673, net214674, net214675, net214677,
         net214678, net214680, net214681, net214683, net214685, net214686,
         net214688, net214690, net214691, net214724, net214729, net214730,
         net214735, net214736, net214737, net214738, net214739, net214740,
         net214744, net214746, net214748, net214750, net214752, net214754,
         net214755, net214756, net214757, net214758, net214759, net214762,
         net214763, net214766, net214767, net214774, net214777, net214778,
         net214781, net214782, net214783, net214786, net214787, net214879,
         net214882, net214952, net214955, net214958, net214960, net214961,
         net214962, net214963, net214964, net214970, net214973, net214979,
         net214981, net214982, net214984, net214985, net214988, net214989,
         net214990, net214991, net214997, net214998, net214999, net215000,
         net215004, net215005, net215013, net215014, net215015, net215016,
         net215017, net215018, net215020, net215021, net215022, net215023,
         net215040, net215041, net215042, net215043, net215044, net215045,
         net215049, net215050, net215051, net215052, net215053, net215054,
         net215057, net215059, net215060, net215061, net215062, net215063,
         net215069, net215070, net215071, net215072, net215078, net215079,
         net215080, net215081, net215093, net215095, net215096, net215097,
         net215098, net215099, net215102, net215104, net215114, net215116,
         net215117, net215119, net215120, net215121, net215122, net215123,
         net215124, net215125, net215126, net215129, net215131, net215132,
         net215134, net215135, net215141, net215143, net215144, net215146,
         net215147, net215148, net215149, net215155, net215156, net215158,
         net215164, net215165, net215166, net215167, net215182, net215183,
         net215186, net215189, net215192, net215194, net215200, net215201,
         net215202, net215203, net215204, net215207, net215209, net215210,
         net215213, net215216, net215222, net215225, net215227, net215228,
         net215231, net215232, net215233, net215271, net215274, net215276,
         net215277, net215279, net215289, net215292, net215294, net215295,
         net215298, net215301, net215304, net215305, net215306, net215312,
         net215313, net215315, net215348, net215349, net215352, net215353,
         net215361, net215362, net215366, net215367, net215369, net215370,
         net215373, net215375, net215376, net215377, net215378, net215385,
         net215386, net215387, net215395, net215396, net215402, net215403,
         net215404, net215405, net215420, net215421, net215429, net215430,
         net215432, net215433, net215434, net215438, net215439, net215465,
         net215466, net215467, net215468, net215818, net215819, net215821,
         net215822, net215825, net215827, net215828, net215831, net215834,
         net215903, net215904, net215905, net215906, net215912, net215915,
         net216020, net216023, net216025, net216026, net216043, net216044,
         net216045, net216046, net216047, net216050, net216137, net216138,
         net216158, net216166, net216167, net216175, net216176, net216180,
         net216183, net216184, net216185, net216189, net216191, net216198,
         net216199, net216201, net216202, net216203, net216207, net216210,
         net216211, net216212, net216216, net216217, net216225, net216226,
         net216229, net216230, net216238, net216239, net216243, net216246,
         net216247, net216248, net216249, net216250, net216253, net216254,
         net216256, net216257, net216258, net216259, net216263, net216264,
         net216265, net216266, net216267, net216268, net216272, net216273,
         net216274, net216275, net216276, net216277, net216283, net216284,
         net216285, net216286, net216290, net216291, net216299, net216300,
         net216301, net216302, net216303, net216304, net216308, net216309,
         net216310, net216311, net216312, net216313, net216319, net216320,
         net216326, net216327, net216328, net216329, net216333, net216334,
         net216336, net216337, net216338, net216344, net216345, net216346,
         net216347, net216348, net216355, net216358, net216360, net216361,
         net216363, net216364, net216365, net216366, net216367, net216394,
         net216396, net216397, net216400, net216403, net216407, net216408,
         net216425, net216426, net216427, net216428, net216434, net216435,
         net216443, net216444, net216461, net216462, net216470, net216471,
         net216488, net216489, net216490, net216491, net216492, net216497,
         net216498, net216499, net216502, net216506, net216507, net216508,
         net216511, net216515, net216516, net216517, net216520, net216594,
         net216595, net216597, net216749, net216750, net216758, net216759,
         net216805, net216808, net216814, net216817, net216868, net216871,
         net216877, net216878, net216879, net216880, net216904, net216907,
         net216913, net216914, net216915, net216916, net217276, net217274,
         net217272, net217270, net217268, net217266, net217264, net217262,
         net217260, net217258, net217256, net217254, net217252, net217250,
         net217248, net217246, net217244, net217242, net217240, net217238,
         net217236, net217234, net217232, net217230, net217228, net217226,
         net217224, net217222, net217220, net217218, net217216, net217214,
         net217212, net217210, net217206, net217202, net217196, net217190,
         net217188, net217186, net217184, net217182, net217180, net217178,
         net217176, net217174, net217172, net217170, net217168, net217166,
         net217164, net217162, net217160, net217158, net217156, net217154,
         net217152, net217150, net217148, net217146, net217144, net217142,
         net217140, net217138, net217136, net217134, net217132, net217128,
         net217126, net217124, net217122, net217120, net217118, net217116,
         net217114, net217112, net217108, net217106, net217104, net217102,
         net217100, net217098, net217096, net217094, net217092, net217088,
         net217086, net217084, net217082, net217080, net217078, net217076,
         net217074, net217072, net217070, net217068, net217066, net217064,
         net217062, net217060, net217058, net217056, net217054, net217052,
         net217050, net217048, net217046, net217044, net217042, net217038,
         net217036, net217034, net217032, net217030, net217028, net217026,
         net217024, net217022, net217020, net217018, net217016, net217012,
         net217010, net217008, net217004, net217002, net217000, net216998,
         net216996, net216994, net216992, net216990, net216988, net216986,
         net216984, net216982, net216980, net216978, net216976, net216974,
         net216972, net216970, net216968, net216966, net216964, net216962,
         net217288, net217286, net217284, net217282, net217280, net217278,
         net218278, net218276, net218274, net218272, net218270, net218268,
         net218266, net218264, net218262, net218260, net218258, net218256,
         net218254, net218252, net218250, net218248, net218246, net218244,
         net218242, net218240, net218238, net218236, net218234, net218232,
         net218230, net218228, net218226, net218224, net218222, net218220,
         net218218, net218216, net218214, net218212, net218210, net218208,
         net218206, net218204, net218202, net218200, net218198, net218196,
         net218194, net218192, net218190, net218188, net218186, net218184,
         net218182, net218180, net218178, net218176, net218174, net218172,
         net218170, net218168, net218166, net218164, net218162, net218160,
         net218158, net218156, net218154, net218152, net218150, net218148,
         net218146, net218144, net218138, net218136, net218132, net218130,
         net218128, net218126, net218124, net218122, net218120, net218118,
         net218116, net218114, net218112, net218110, net218108, net218106,
         net218104, net218102, net218100, net218098, net218096, net218094,
         net218092, net218090, net218088, net218086, net218084, net218082,
         net218080, net218078, net218076, net218074, net218072, net218070,
         net218068, net218066, net218064, net218062, net218060, net218058,
         net218056, net218054, net218052, net218050, net218048, net218046,
         net218044, net218042, net218040, net218038, net218036, net218034,
         net218030, net218028, net218026, net218024, net218022, net218020,
         net218018, net218016, net218014, net218012, net218010, net218008,
         net218006, net218004, net218002, net218000, net217998, net217996,
         net217994, net217992, net217990, net217988, net217986, net217984,
         net217982, net217980, net217978, net217976, net217974, net217972,
         net217970, net217968, net217964, net217962, net217960, net217956,
         net217954, net217952, net217950, net217946, net217944, net217942,
         net217940, net217938, net217936, net217934, net217932, net217930,
         net218292, net218286, net218284, net218282, net218598, net218596,
         net218594, net218592, net218590, net218588, net218586, net218584,
         net218582, net218580, net218578, net218576, net218574, net218572,
         net218570, net218568, net218566, net218564, net218562, net218560,
         net218558, net218556, net218554, net218552, net218550, net218548,
         net218546, net218544, net218542, net218540, net218538, net218536,
         net218534, net218532, net218530, net218528, net218526, net218524,
         net218520, net218518, net218516, net218512, net218510, net218508,
         net218506, net218504, net218502, net218500, net218496, net218494,
         net218490, net218488, net218486, net218484, net218482, net218480,
         net218478, net218476, net218474, net218472, net218468, net218464,
         net218462, net218458, net218456, net218454, net218452, net218450,
         net218446, net218442, net218440, net218438, net218434, net218432,
         net218430, net218428, net218426, net218424, net218422, net218420,
         net218418, net218416, net218414, net218412, net218410, net218408,
         net218406, net218404, net218402, net218400, net218398, net218396,
         net218394, net218392, net218388, net218386, net218384, net218380,
         net218378, net218376, net218374, net218372, net218370, net218368,
         net218366, net218364, net218360, net218358, net218356, net218354,
         net218352, net218350, net218348, net218346, net218344, net218342,
         net218340, net218338, net218336, net218334, net218332, net218330,
         net218328, net218326, net218324, net218322, net218320, net218316,
         net218314, net218312, net218310, net218308, net218304, net218302,
         net218300, net218298, net218296, net218294, net218606, net218604,
         net218602, net218954, net218952, net218950, net218948, net218946,
         net218944, net218942, net218940, net218938, net218936, net218934,
         net218932, net218930, net218928, net218926, net218924, net218922,
         net218920, net218918, net218916, net218914, net218912, net218910,
         net218908, net218906, net218904, net218902, net218900, net218898,
         net218896, net218894, net218892, net218890, net218888, net218886,
         net218884, net218882, net218880, net218878, net218876, net218874,
         net218872, net218870, net218868, net218866, net218864, net218862,
         net218860, net218856, net218854, net218852, net218850, net218848,
         net218846, net218844, net218842, net218840, net218838, net218836,
         net218834, net218832, net218830, net218828, net218824, net218822,
         net218820, net218818, net218816, net218814, net218812, net218810,
         net218808, net218806, net218804, net218802, net218800, net218798,
         net218796, net218794, net218792, net218790, net218788, net218786,
         net218782, net218780, net218778, net218776, net218774, net218772,
         net218770, net218768, net218766, net218764, net218762, net218760,
         net218758, net218756, net218754, net218752, net218750, net218748,
         net218746, net218744, net218742, net218740, net218738, net218736,
         net218732, net218730, net218728, net218724, net218722, net218720,
         net218716, net218712, net218710, net218708, net218704, net218702,
         net218700, net218698, net218696, net218694, net218688, net218684,
         net218680, net218678, net218676, net218674, net218672, net218670,
         net218668, net218666, net218664, net218660, net218658, net218656,
         net218654, net218652, net218650, net218648, net218646, net218644,
         net218642, net218640, net218636, net218634, net218632, net218628,
         net218626, net218624, net218622, net218620, net218618, net218616,
         net218614, net218612, net218610, net218966, net218964, net218962,
         net218960, net218958, net218956, net219356, net219346, net219336,
         net219330, net219324, net219322, net219314, net219310, net219308,
         net219492, net219484, net219480, net219478, net219472, net219468,
         net219466, net219460, net219450, net219444, net219442, net219434,
         net219494, net221988, net221986, net221984, net221982, net221980,
         net221978, net221976, net221974, net221972, net221970, net221968,
         net221966, net221964, net221962, net221960, net221956, net221954,
         net221952, net221950, net221948, net221946, net221944, net221942,
         net221940, net221938, net221936, net221934, net221932, net221930,
         net221928, net221926, net221924, net221922, net221920, net221918,
         net221916, net221914, net221912, net221910, net221908, net221906,
         net221904, net221902, net221900, net221894, net221892, net221890,
         net221888, net221886, net221884, net221882, net221880, net221878,
         net221874, net221872, net221870, net221868, net221866, net221864,
         net221862, net221860, net221858, net221856, net221854, net221852,
         net221850, net221848, net221846, net221844, net221840, net221838,
         net221836, net221834, net221832, net221830, net221828, net221826,
         net221824, net221822, net221820, net221818, net221816, net221814,
         net221812, net221810, net221808, net221806, net221804, net221802,
         net221800, net221798, net221796, net221794, net221792, net221790,
         net221788, net221786, net221784, net221780, net221778, net221776,
         net221774, net221772, net221770, net221768, net221766, net221764,
         net221762, net221760, net221758, net221756, net221754, net221752,
         net221744, net221740, net221736, net221734, net221732, net221730,
         net221726, net221724, net221722, net221720, net221718, net221716,
         net221992, net221990, net234007, net234488, net234521, net234523,
         net234527, net234529, net234760, net234762, net234998, net235251,
         net236115, net238789, net238790, net238801, net238868, net238947,
         net256309, net258199, net258207, net258262, net258261, net258320,
         net258903, net258961, net259019, net259031, net259034, net259626,
         net259641, net259645, net259649, net259653, net259661, net259665,
         net259677, net259747, net259841, net259873, net260247, net260251,
         net260277, net260295, net260299, net260302, net260332, net260346,
         net260352, net260355, net260367, net260376, net260384, net260394,
         net260403, net260412, net260427, net260431, net260449, net260461,
         net260470, net260474, net260488, net260492, net260494, net260527,
         net260830, net260900, net260925, net261020, net261069, net261422,
         net261867, net261886, net261905, net261924, net261943, net261981,
         net262000, net262019, net262038, net262057, net262095, net262114,
         net262133, net262152, net262171, net262190, net262209, net262228,
         net262247, net262266, net262285, net262304, net262323, net262342,
         net262361, net262380, net262399, net262418, net262437, net262456,
         net262475, net262513, net262532, net262551, net262570, net262589,
         net262608, net262627, net262646, net262665, net262703, net262722,
         net262741, net262779, net262798, net262817, net262836, net262855,
         net262874, net262893, net262912, net262931, net262950, net262969,
         net262988, net263007, net263026, net263045, net263064, net263083,
         net263102, net263121, net263140, net263159, net263178, net263216,
         net263235, net263254, net263292, net263330, net263349, net263368,
         net263387, net263406, net263444, net263463, net263501, net263539,
         net263558, net263577, net263596, net263615, net263634, net263653,
         net263672, net263691, net263710, net263748, net263767, net263805,
         net263824, net263843, net263862, net263881, net263900, net263919,
         net263957, net263976, net263995, net264532, net264577, net264592,
         net264607, net264652, net264682, net264712, net264742, net264808,
         net264827, net264846, net264865, net264884, net264903, net264922,
         net264941, net264960, net264979, net264998, net265017, net265036,
         net265055, net265074, net265112, net265131, net265150, net265169,
         net265188, net265207, net265226, net265245, net265264, net265283,
         net265302, net265321, net265340, net265359, net265378, net265397,
         net265416, net265435, net265454, net265473, net265492, net265511,
         net265530, net265549, net265568, net265587, net265606, net265625,
         net265644, net265682, net265701, net265720, net265739, net265758,
         net265777, net265796, net265815, net265834, net265853, net265872,
         net265891, net265910, net265929, net265948, net265967, net266005,
         net266024, net266043, net266062, net266081, net266100, net266119,
         net266151, net266201, net266218, net266235, net266255, net266276,
         net266297, net266318, net266339, net266360, net266381, net266402,
         net266423, net266444, net266465, net266486, net266507, net266528,
         net266549, net266570, net266591, net266612, net266633, net266654,
         net266675, net266696, net266717, net266738, net266759, net266780,
         n_cell_301249_net269969, n_cell_301249_net269950,
         n_cell_301249_net269943, n_cell_301249_net269941,
         n_cell_301249_net269874, n_cell_301249_net269872,
         n_cell_301249_net269861, n_cell_301249_net269853,
         n_cell_301249_net269839, n_cell_301249_net269836,
         n_cell_301249_net269831, n_cell_301249_net269828,
         n_cell_301249_net269811, n_cell_301249_net269798,
         n_cell_301249_net269797, n_cell_301249_net269794,
         n_cell_301249_net269764, n_cell_301249_net269763,
         n_cell_301249_net269758, n_cell_301249_net269755,
         n_cell_301249_net269749, n_cell_301249_net269746,
         n_cell_301249_net269745, n_cell_301249_net269740,
         n_cell_301249_net269738, n_cell_301249_net269731,
         n_cell_301249_net269714, n_cell_301249_net269711,
         n_cell_301249_net269701, n_cell_301249_net269688,
         n_cell_301249_net269653, n_cell_301249_net269650,
         n_cell_301249_net269647, n_cell_301249_net269646,
         n_cell_301249_net269638, n_cell_301249_net269635,
         n_cell_301249_net269615, n_cell_301249_net269613,
         n_cell_301249_net269596, n_cell_301249_net269593,
         n_cell_301249_net269590, n_cell_301249_net269583,
         n_cell_301249_net269578, n_cell_301249_net269571,
         n_cell_301249_net269568, n_cell_301249_net269564,
         n_cell_301249_net269488, n_cell_301249_net269482,
         n_cell_301249_net269481, n_cell_301249_net269478,
         n_cell_301249_net269477, n_cell_301249_net269475,
         n_cell_301249_net269449, n_cell_301249_net269022,
         n_cell_301249_net268916, n_cell_301249_net268398,
         n_cell_301249_net268392, n_cell_301249_net268386,
         n_cell_301249_net268380, n_cell_301249_net268355,
         n_cell_301249_net268342, n_cell_301249_net268336,
         n_cell_301249_net268272, n_cell_301249_net268242,
         n_cell_301249_net268236, n_cell_301249_net268223,
         n_cell_301249_net268217, n_cell_301249_net268196,
         n_cell_301249_net268190, n_cell_301249_net268172,
         n_cell_301249_net268166, n_cell_301249_net268160,
         n_cell_301249_net268154, n_cell_301249_net268142,
         n_cell_301249_net268136, n_cell_301249_net268109,
         n_cell_301249_net268103, n_cell_301249_net268097,
         n_cell_301249_net268091, n_cell_301249_net268085,
         n_cell_301249_net268079, n_cell_301249_net268071,
         n_cell_301249_net268065, n_cell_301249_net268056,
         n_cell_301249_net268044, n_cell_301249_net268038,
         n_cell_301249_net268029, n_cell_301249_net268023,
         n_cell_301249_net268002, n_cell_301249_net267980,
         n_cell_301249_net267966, n_cell_301249_net267960,
         n_cell_301249_net267948, n_cell_301249_net267932,
         n_cell_301249_net267909, n_cell_301249_net267903,
         n_cell_301249_net267891, n_cell_301249_net267885,
         n_cell_301249_net267867, n_cell_301249_net267855,
         n_cell_301249_net267846, n_cell_301249_net267840,
         n_cell_301249_net267828, n_cell_301249_net267822,
         n_cell_301249_net267810, n_cell_301249_net267804,
         n_cell_301249_net267786, n_cell_301249_net267780,
         n_cell_301249_net267769, n_cell_301249_net267763,
         n_cell_301249_net267754, n_cell_301249_net267742,
         n_cell_301249_net267706, n_cell_301249_net267700,
         n_cell_301249_net267694, n_cell_301249_net267688,
         n_cell_301249_net267682, n_cell_301249_net267676,
         n_cell_301249_net267670, n_cell_301249_net267658,
         n_cell_301249_net267652, n_cell_301249_net267646,
         n_cell_301249_net267640, n_cell_301249_net267628,
         n_cell_301249_net267619, n_cell_301249_net267613,
         n_cell_301249_net267607, n_cell_301249_net267601,
         n_cell_301249_net267595, n_cell_301249_net267589,
         n_cell_301249_net267580, n_cell_301249_net267574,
         n_cell_301249_net267562, n_cell_301249_net267556,
         n_cell_301249_net267550, n_cell_301249_net267526,
         n_cell_301249_net267516, n_cell_301249_net267510,
         n_cell_301249_net267490, n_cell_301249_net267484,
         n_cell_301249_net267466, n_cell_301249_net267451,
         n_cell_301249_net267447, n_cell_301249_net267441,
         n_cell_301249_net267429, n_cell_301249_net267415,
         n_cell_301249_net267409, n_cell_301249_net267397,
         n_cell_301249_net267391, n_cell_301249_net267385,
         n_cell_301249_net267379, n_cell_301249_net267373,
         n_cell_301249_net267349, n_cell_301249_net267343,
         n_cell_301249_net267337, n_cell_301249_net267331,
         n_cell_301249_net267325, n_cell_301249_net267319,
         n_cell_301249_net267308, n_cell_301249_net267302,
         n_cell_301249_net267275, n_cell_301249_net267269,
         n_cell_301249_net267263, n_cell_301249_net267257,
         n_cell_301249_net267239, n_cell_301249_net267233,
         n_cell_301249_net267225, n_cell_301249_net267219,
         n_cell_301249_net267213, n_cell_301249_net267207,
         n_cell_301249_net267201, n_cell_301249_net267189,
         n_cell_301249_net267183, n_cell_301249_net267171,
         n_cell_301249_net267165, n_cell_301249_net267141,
         n_cell_301249_net267135, n_cell_301249_net267123,
         n_cell_301249_net267117, n_cell_301249_net267095,
         n_cell_301249_net267089, n_cell_301249_net267075,
         n_cell_301249_net267063, n_cell_301249_net266950,
         n_cell_301249_net266944, n_cell_301249_net266916, net271431,
         net271515, net271956, net271996, net271999, net272417, net272583,
         net272620, net272625, n_cell_303546_net278017,
         n_cell_303546_net277994, n_cell_303546_net277957,
         n_cell_303546_net277942, n_cell_303546_net277936,
         n_cell_303546_net277892, n_cell_303546_net277859,
         n_cell_303546_net277854, n_cell_303546_net277852,
         n_cell_303546_net277843, n_cell_303546_net277834,
         n_cell_303546_net277822, n_cell_303546_net277814,
         n_cell_303546_net277804, n_cell_303546_net277795,
         n_cell_303546_net277772, n_cell_303546_net277761,
         n_cell_303546_net277759, n_cell_303546_net277738,
         n_cell_303546_net277735, n_cell_303546_net277698,
         n_cell_303546_net277696, n_cell_303546_net277671,
         n_cell_303546_net277667, n_cell_303546_net277645,
         n_cell_303546_net277636, n_cell_303546_net277632,
         n_cell_303546_net277630, n_cell_303546_net277551,
         n_cell_303546_net277536, n_cell_303546_net277530,
         n_cell_303546_net277506, n_cell_303546_net277497,
         n_cell_303546_net277496, n_cell_303546_net277494,
         n_cell_303546_net277490, n_cell_303546_net277470,
         n_cell_303546_net277469, n_cell_303546_net277412,
         n_cell_303546_net277405, n_cell_303546_net276554,
         n_cell_303546_net276365, n_cell_303546_net276178,
         n_cell_303546_net276009, n_cell_303546_net275998,
         n_cell_303546_net275987, n_cell_303546_net275967,
         n_cell_303546_net275959, n_cell_303546_net275956,
         n_cell_303546_net275934, n_cell_303546_net275923,
         n_cell_303546_net275906, n36638, n36639, n36640, n36641, n36642,
         n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650,
         n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658,
         n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666,
         n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674,
         n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682,
         n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690,
         n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698,
         n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706,
         n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714,
         n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722,
         n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
         n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
         n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
         n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754,
         n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762,
         n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770,
         n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778,
         n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786,
         n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794,
         n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802,
         n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810,
         n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818,
         n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826,
         n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834,
         n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842,
         n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850,
         n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858,
         n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866,
         n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874,
         n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882,
         n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890,
         n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898,
         n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906,
         n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914,
         n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922,
         n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930,
         n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938,
         n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946,
         n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954,
         n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962,
         n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970,
         n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978,
         n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986,
         n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994,
         n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002,
         n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010,
         n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018,
         n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026,
         n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034,
         n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042,
         n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050,
         n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058,
         n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066,
         n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074,
         n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082,
         n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
         n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098,
         n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106,
         n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114,
         n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122,
         n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130,
         n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138,
         n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146,
         n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154,
         n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
         n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170,
         n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178,
         n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186,
         n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194,
         n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202,
         n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210,
         n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218,
         n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226,
         n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
         n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242,
         n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250,
         n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258,
         n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266,
         n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274,
         n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282,
         n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290,
         n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298,
         n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
         n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314,
         n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322,
         n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330,
         n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338,
         n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346,
         n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354,
         n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362,
         n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370,
         n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378,
         n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386,
         n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394,
         n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402,
         n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410,
         n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418,
         n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426,
         n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434,
         n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442,
         n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450,
         n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458,
         n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466,
         n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474,
         n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482,
         n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490,
         n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498,
         n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506,
         n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514,
         n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522,
         n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530,
         n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538,
         n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546,
         n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554,
         n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596,
         n37597, n37598, n37599, n37600, n37601, n39282, n39283, n39284,
         n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292,
         n39293, n39294, n39295, n39296, n39297, n39298, n39299, n39300,
         n39301, n39302, n39303, n39304, n39305, n39306, n39307, n39308,
         n39309, n39310, n39311, n39312, n39313, n39314, n39315, n39316,
         n39317, n39318, n39319, n39320, n39321, n39322, n39323, n39324,
         n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39332,
         n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340,
         n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348,
         n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356,
         n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364,
         n39365, n39366, n39367, n39368, n39369, n39370, n39371, n39372,
         n39373, n39374, n39375, n39376, n39377, n39378, n39379, n39380,
         n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388,
         n39389, n39390, n39391, n39392, n39393, n39394, n39395, n39396,
         n39397, n39398, n39399, n39400, n39401, n39402, n39403, n39404,
         n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412,
         n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420,
         n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428,
         n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436,
         n39437, n39438, n39439, n39440, n39441, n39442, n39443, n39444,
         n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452,
         n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460,
         n39461, n39462, n39463, n39464, n39465, n39466, n39467, n39468,
         n39469, n39470, n39471, n39472, n39473, n39474, n39475, n39476,
         n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484,
         n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492,
         n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500,
         n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508,
         n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516,
         n39517, n39518, n39519, n39520, n39521, n39522, n39523, n39524,
         n39525, n39526, n39527, n39528, n39529, n39530, n39531, n39532,
         n39533, n39534, n39535, n39536, n39537, n39538, n39539, n39540,
         n39541, n39542, n39543, n39544, n39545, n39546, n39547, n39548,
         n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556,
         n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564,
         n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572,
         n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580,
         n39581, n39582, n39583, n39584, n39585, n39586, n39587, n39588,
         n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596,
         n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604,
         n39605, n39606, n39607, n39608, n39609, n39610, n39611, n39612,
         n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39620,
         n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628,
         n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636,
         n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644,
         n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652,
         n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660,
         n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668,
         n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676,
         n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684,
         n39685, n39686, n39687, n39688, n39689, n39690, n39691, n39692,
         n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700,
         n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708,
         n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716,
         n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724,
         n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732,
         n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740,
         n39741, n39742, n39743, n39744, n39745, n39746, n39747, n39748,
         n39749, n39750, n39751, n39752, n39753, n39754, n39755, n39756,
         n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764,
         n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772,
         n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780,
         n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788,
         n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796,
         n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804,
         n39805, n39806, n39807, n39808, n39809, n39810, n39811, n39812,
         n39813, n39814, n39815, n39816, n39817, n39818, n39819, n39820,
         n39821, n39822, n39823, n39824, n39825, n39826, n39827, n39828,
         n39829, n39830, n39831, n39832, n39833, n39834, n39835, n39836,
         n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844,
         n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852,
         n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860,
         n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868,
         n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876,
         n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884,
         n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892,
         n39893, n39894, n39895, n39896, n39897, n39898, n39899, n39900,
         n39901, n39902, n39903, n39904, n39905, n39906, n39907, n39908,
         n39909, n39910, n39911, n39912, n39913, n39914, n39915, n39916,
         n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924,
         n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932,
         n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940,
         n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948,
         n39949, n39950, n39951, n39952, n39953, n39954, n39955, n39956,
         n39957, n39958, n39959, n39960, n39961, n39962, n39963, n39964,
         n39965, n39966, n39967, n39968, n39969, n39970, n39971, n39972,
         n39973, n39974, n39975, n39976, n39977, n39978, n39979, n39980,
         n39981, n39982, n39983, n39984, n39985, n39986, n39987, n39988,
         n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996,
         n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004,
         n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012,
         n40013, n40014, n40015, n40016, n40017, n40018, n40019, n40020,
         n40021, n40022, n40023, n40024, n40025, n40026, n40027, n40028,
         n40029, n40030, n40031, n40032, n40033, n40034, n40035, n40036,
         n40037, n40038, n40039, n40040, n40041, n40042, n40043, n40044,
         n40045, n40046, n40047, n40048, n40049, n40050, n40051, n40052,
         n40053, n40054, n40055, n40056, n40057, n40058, n40059, n40060,
         n40061, n40062, n40063, n40064, n40065, n40066, n40067, n40068,
         n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076,
         n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084,
         n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092,
         n40093, n40094, n40095, n40096, n40097, n40098, n40099, n40100,
         n40101, n40102, n40103, n40104, n40105, n40106, n40107, n40108,
         n40109, n40110, n40111, n40112, n40113, n40114, n40115, n40116,
         n40117, n40118, n40119, n40120, n40121, n40122, n40123, n40124,
         n40125, n40126, n40127, n40128, n40129, n40130, n40131, n40132,
         n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140,
         n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148,
         n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156,
         n40157, n40158, n40159, n40160, n40161, n40162, n40163, n40164,
         n40165, n40166, n40167, n40168, n40169, n40170, n40171, n40172,
         n40173, n40174, n40175, n40176, n40177, n40178, n40179, n40180,
         n40181, n40182, n40183, n40184, n40185, n40186, n40187, n40188,
         n40189, n40190, n40191, n40192, n40193, n40194, n40195, n40196,
         n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204,
         n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212,
         n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220,
         n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228,
         n40229, n40230, n40231, n40232, n40233, n40234, n40235, n40236,
         n40237, n40238, n40239, n40240, n40241, n40242, n40243, n40244,
         n40245, n40246, n40247, n40248, n40249, n40250, n40251, n40252,
         n40253, n40254, n40255, n40256, n40257, n40258, n40259, n40260,
         n40261, n40262, n40263, n40264, n40265, n40266, n40267, n40268,
         n40269, n40270, n40271, n40272, n40273, n40274, n40275, n40276,
         n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284,
         n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292,
         n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300,
         n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308,
         n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316,
         n40317, n40318, n40319, n40320, n40321, n40322, n40323, n40324,
         n40325, n40326, n40327, n40328, n40329, n40330, n40331, n40332,
         n40333, n40334, n40335, n40336, n40337, n40338, n40339, n40340,
         n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348,
         n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356,
         n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364,
         n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372,
         n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380,
         n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388,
         n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396,
         n40397, n40398, n40399, n40400, n40401, n40402, n40403, n40404,
         n40405, n40406, n40407, n40408, n40409, n40410, n40411, n40412,
         n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420,
         n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428,
         n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436,
         n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444,
         n40445, n40446, n40447, n40448, n40449, n40450, n40451, n40452,
         n40453, n40454, n40455, n40456, n40457, n40458, n40459, n40460,
         n40461, n40462, n40463, n40464, n40465, n40466, n40467, n40468,
         n40469, n40470, n40471, n40472, n40473, n40474, n40475, n40476,
         n40477, n40478, n40479, n40480, n40481, n40482, n40483, n40484,
         n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492,
         n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500,
         n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508,
         n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516,
         n40517, n40518, n40519, n40520, n40521, n40522, n40523, n40524,
         n40525, n40526, n40527, n40528, n40529, n40530, n40531, n40532,
         n40533, n40534, n40535, n40536, n40537, n40538, n40539, n40540,
         n40541, n40542, n40543, n40544, n40545, n40546, n40547, n40548,
         n40549, n40550, n40551, n40552, n40553, n40554, n40555, n40556,
         n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564,
         n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572,
         n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580,
         n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588,
         n40589, n40590, n40591, n40592, n40593, n40594, n40595, n40596,
         n40597, n40598, n40599, n40600, n40601, n40602, n40603, n40604,
         n40605, n40606, n40607, n40608, n40609, n40610, n40611, n40612,
         n40613, n40614, n40615, n40616, n40617, n40618, n40619, n40620,
         n40621, n40622, n40623, n40624, n40625, n40626, n40627, n40628,
         n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636,
         n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644,
         n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652,
         n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660,
         n40661, n40662, n40663, n40664, n40665, n40666, n40667, n40668,
         n40669, n40670, n40671, n40672, n40673, n40674, n40675, n40676,
         n40677, n40678, n40679, n40680, n40681, n40682, n40683, n40684,
         n40685, n40686, n40687, n40688, n40689, n40690, n40691, n40692,
         n40693, n40694, n40695, n40696, n40697, n40698, n40699, n40700,
         n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708,
         n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716,
         n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724,
         n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732,
         n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740,
         n40741, n40742, n40743, n40744, n40745, n40746, n40747, n40748,
         n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756,
         n40757, n40758, n40759, n40760, n40761, n40762, n40763, n40764,
         n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772,
         n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780,
         n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788,
         n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796,
         n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804,
         n40805, n40806, n40807, n40808, n40809, n40810, n40811, n40812,
         n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820,
         n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40828,
         n40829, n40830, n40831, n40832, n40833, n40834, n40835, n40836,
         n40837, n40838, n40839, n40840, n40841, n40842, n40843, n40844,
         n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852,
         n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860,
         n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868,
         n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876,
         n40877, n40878, n40879, n40880, n40881, n40882, n40883, n40884,
         n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892,
         n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900,
         n40901, n40902, n40903, n40904, n40905, n40906, n40907, n40908,
         n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916,
         n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924,
         n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932,
         n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940,
         n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948,
         n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956,
         n40957, n40958, n40959, n40960, n40961, n40962, n40963, n40964,
         n40965, n40966, n40967, n40968, n40969, n40970, n40971, n40972,
         n40973, n40974, n40975, n40976, n40977, n40978, n40979, n40980,
         n40981, n40982, n40983, n40984, n40985, n40986, n40987, n40988,
         n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996,
         n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004,
         n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012,
         n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020,
         n41021, n41022, n41023, n41024, n41025, n41026, n41027, n41028,
         n41029, n41030, n41031, n41032, n41033, n41034, n41035, n41036,
         n41037, n41038, n41039, n41040, n41041, n41042, n41043, n41044,
         n41045, n41046, n41047, n41048, n41049, n41050, n41051, n41052,
         n41053, n41054, n41055, n41056, n41057, n41058, n41059, n41060,
         n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068,
         n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076,
         n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084,
         n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092,
         n41093, n41094, n41095, n41096, n41097, n41098, n41099, n41100,
         n41101, n41102, n41103, n41104, n41105, n41106, n41107, n41108,
         n41109, n41110, n41111, n41112, n41113, n41114, n41115, n41116,
         n41117, n41118, n41119, n41120, n41121, n41122, n41123, n41124,
         n41125, n41126, n41127, n41128, n41129, n41130, n41131, n41132,
         n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140,
         n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148,
         n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156,
         n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164,
         n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172,
         n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180,
         n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188,
         n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41196,
         n41198, n41199, n41200, n41201, n41202, n41203, n41204, n41205,
         n41206, n41207, n41208, n41209, n41210, n41211, n41212, n41213,
         n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221,
         n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229,
         n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237,
         n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245,
         n41246, n41247, n41248, n41249, n41250, n41251, n41252, n41253,
         n41254, n41255, n41256, n41257, n41258, n41259, n41260, n41261,
         n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269,
         n41270, n41271, n41272, n41273, n41274, n41275, n41276, n41277,
         n41278, n41279, n41280, n41281, n41282, n41283, n41284, n41285,
         n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293,
         n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301,
         n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309,
         n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317,
         n41318, n41319, n41320, n41321, n41322, n41323, n41324, n41325,
         n41326, n41327, n41328, n41329, n41330, n41331, n41332, n41333,
         n41334, n41335, n41343, n41344, n41345, n41346, n41347, n41348,
         n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356,
         n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364,
         n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372,
         n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380,
         n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388,
         n41389, n41390, n41629, n41630, n41631, n41632, n41633, n41634,
         n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642,
         n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650,
         n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658,
         n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666,
         n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674,
         n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682,
         n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690,
         n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698,
         n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706,
         n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714,
         n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726,
         n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734,
         n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742,
         n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750,
         n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758,
         n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766,
         n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774,
         n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782,
         n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790,
         n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798,
         n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806,
         n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814,
         n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822,
         n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830,
         n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838,
         n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846,
         n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854,
         n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862,
         n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870,
         n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878,
         n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886,
         n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894,
         n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902,
         n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910,
         n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918,
         n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926,
         n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934,
         n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942,
         n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950,
         n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958,
         n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966,
         n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974,
         n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982,
         n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990,
         n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998,
         n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006,
         n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014,
         n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022,
         n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030,
         n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038,
         n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046,
         n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054,
         n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062,
         n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070,
         n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078,
         n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086,
         n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094,
         n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102,
         n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110,
         n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118,
         n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126,
         n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134,
         n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142,
         n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150,
         n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158,
         n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166,
         n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174,
         n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182,
         n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190,
         n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198,
         n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206,
         n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214,
         n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222,
         n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230,
         n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238,
         n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246,
         n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254,
         n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262,
         n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270,
         n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278,
         n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286,
         n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294,
         n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302,
         n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310,
         n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318,
         n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326,
         n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334,
         n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342,
         n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350,
         n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358,
         n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366,
         n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374,
         n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382,
         n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390,
         n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398,
         n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406,
         n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414,
         n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422,
         n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430,
         n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438,
         n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446,
         n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454,
         n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462,
         n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470,
         n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478,
         n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486,
         n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494,
         n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502,
         n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510,
         n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518,
         n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526,
         n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534,
         n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542,
         n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550,
         n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558,
         n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566,
         n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574,
         n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582,
         n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590,
         n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
         n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606,
         n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614,
         n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622,
         n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630,
         n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638,
         n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646,
         n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654,
         n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662,
         n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670,
         n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678,
         n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686,
         n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694,
         n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702,
         n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710,
         n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718,
         n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726,
         n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734,
         n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742,
         n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750,
         n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758,
         n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766,
         n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774,
         n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782,
         n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790,
         n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798,
         n42799, n42800, n42801, n42802, n42803, n42804, n42805, n42806,
         n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814,
         n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822,
         n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830,
         n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838,
         n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846,
         n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854,
         n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862,
         n42863, n42864, n42865, n42866, n42867, n42868, n42869, n42870,
         n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878,
         n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886,
         n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894,
         n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902,
         n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910,
         n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918,
         n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926,
         n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934,
         n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942,
         n42943, n42944, n42945, n42946, n42947, n42948, n42949, n42950,
         n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958,
         n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966,
         n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974,
         n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982,
         n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990,
         n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998,
         n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006,
         n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014,
         n43015, n43016, n43017, n43018, n43019, n43020, n43021, n43022,
         n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030,
         n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038,
         n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046,
         n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054,
         n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062,
         n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070,
         n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078,
         n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086,
         n43087, n43088, n43089, n43090, n43091, n43092, n43093, n43094,
         n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102,
         n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110,
         n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118,
         n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126,
         n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134,
         n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142,
         n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150,
         n43151, n43152, n43153, n43154, n43155, n43156, n43157, n43158,
         n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43166,
         n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174,
         n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182,
         n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190,
         n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198,
         n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206,
         n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214,
         n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222,
         n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230,
         n43231, n43232, n43233, n43234, n43235, n43236, n43237, n43238,
         n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246,
         n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254,
         n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262,
         n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270,
         n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278,
         n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286,
         n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294,
         n43295, n43296, n43297, n43298, n43299, n43300, n43301, n43302,
         n43303, n43304, n43305, n43306, n43307, n43308, n43309, n43310,
         n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318,
         n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326,
         n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334,
         n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342,
         n43343, n43344, n43345, n43346, n43347, n43348, n43349, n43350,
         n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358,
         n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366,
         n43367, n43368, n43369, n43370, n43371, n43372, n43373, n43374,
         n43375, n43376, n43377, n43378, n43379, n43380, n43381, n43382,
         n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390,
         n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398,
         n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406,
         n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414,
         n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422,
         n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430,
         n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438,
         n43439, n43440, n43441, n43442, n43443, n43444, n43445, n43446,
         n43447, n43448, n43449, n43450, n43451, n43452, n43453, n43454,
         n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462,
         n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470,
         n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478,
         n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486,
         n43487, n43488, n43489, n43490, n43491, n43492, n43493, n43494,
         n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502,
         n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510,
         n43511, n43512, n43513, n43514, n43515, n43516, n43517, n43518,
         n43519, n43520, n43521, n43522, n43523, n43524, n43525, n43526,
         n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534,
         n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542,
         n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550,
         n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558,
         n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566,
         n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574,
         n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582,
         n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590,
         n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598,
         n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606,
         n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614,
         n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622,
         n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630,
         n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638,
         n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646,
         n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654,
         n43655, n43656, n43657, n43658, n43659, n43660, n43661, n43662,
         n43663, n43664, n43665, n43666, n43667, n43668, n43669, n43670,
         n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678,
         n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686,
         n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694,
         n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702,
         n43703, n43704, n43705, n43706, n43707, n43708, n43709, n43710,
         n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718,
         n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726,
         n43727, n43728, n43729, n43730, n43731, n43732, n43733, n43734,
         n43735, n43736, n43737, n43738, n43739, n43740, n43741, n43742,
         n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750,
         n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758,
         n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766,
         n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774,
         n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782,
         n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790,
         n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798,
         n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806,
         n43807, n43808, n43809, n43810, n43811, n43812, n43813, n43814,
         n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822,
         n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830,
         n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838,
         n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846,
         n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854,
         n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862,
         n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870,
         n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878,
         n43879, n43880, n43881, n43882, n43883, n43884, n43885, n43886,
         n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894,
         n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902,
         n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910,
         n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918,
         n43919, n43920, n43921, n43922, n43923, n43924, n43925, n43926,
         n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934,
         n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942,
         n43943, n43944, n43945, n43946, n43947, n43948, n43949, n43950,
         n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958,
         n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966,
         n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974,
         n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982,
         n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990,
         n43991, n43992, n43993, n43994, n43995, n43996, n43997, n43998,
         n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006,
         n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014,
         n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022,
         n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030,
         n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038,
         n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046,
         n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054,
         n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062,
         n44063, n44064, n44065, n44066, n44067, n44068, n44069, n44070,
         n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078,
         n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086,
         n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094,
         n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102,
         n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110,
         n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118,
         n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126,
         n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134,
         n44135, n44136, n44137, n44138, n44139, n44140, n44141, n44142,
         n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150,
         n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158,
         n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166,
         n44167, n44168, n44169, n44170, n44171, n44172, n44173, n44174,
         n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182,
         n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190,
         n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198,
         n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206,
         n44207, n44208, n44209, n44210, n44211, n44212, n44213, n44214,
         n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222,
         n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230,
         n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238,
         n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246,
         n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254,
         n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262,
         n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270,
         n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278,
         n44279, n44280, n44281, n44282, n44283, n44284, n44285, n44286,
         n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294,
         n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302,
         n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310,
         n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318,
         n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326,
         n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334,
         n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342,
         n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350,
         n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358,
         n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366,
         n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374,
         n44375, n44376, n44377, n44378, n44379, n44380, n44381, n44382,
         n44383, n44384, n44385, n44386, n44387, n44388, n44389, n44390,
         n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398,
         n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406,
         n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414,
         n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422,
         n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430,
         n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438,
         n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446,
         n44447, n44448, n44449, n44450, n44451, n44452, n44453, n44454,
         n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462,
         n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470,
         n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478,
         n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486,
         n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494,
         n44495, n44496, n44497, n44498, n44499, n44500, n44501, n44502,
         n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510,
         n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518,
         n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526,
         n44527, n44528, n44529, n44530, n44531, n44532, n44533, n44534,
         n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542,
         n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550,
         n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558,
         n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566,
         n44567, n44568, n44569, n44570, n44571, n44572, n44573, n44574,
         n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582,
         n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590,
         n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598,
         n44599, n44600, n44601, n44602, n44603, n44604, n44605, n44606,
         n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614,
         n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622,
         n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630,
         n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638,
         n44639, n44640, n44641, n44642, n44643, n44644, n44645, n44646,
         n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654,
         n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662,
         n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670,
         n44671, n44672, n44673, n44674, n44675, n44676, n44677, n44678,
         n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686,
         n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694,
         n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702,
         n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710,
         n44711, n44712, n44713, n44714, n44715, n44716, n44717, n44718,
         n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726,
         n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734,
         n44735, n44736, n44737, n44738, n44739, n44740, n44741, n44742,
         n44743, n44744, n44745, n44746, n44747, n44748, n44749, n44750,
         n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758,
         n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766,
         n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774,
         n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782,
         n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790,
         n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798,
         n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806,
         n44807, n44808, n44809, n44810, n44811, n44812, n44813, n44814,
         n44815, n44816, n44817, n44818, n44819, n44820, n44821, n44822,
         n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830,
         n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838,
         n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846,
         n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854,
         n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862,
         n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870,
         n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878,
         n44879, n44880, n44881, n44882, n44883, n44884, n44885, n44886,
         n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894,
         n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902,
         n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910,
         n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918,
         n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926,
         n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934,
         n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942,
         n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950,
         n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44958,
         n44959, n44960, n44961, n44962, n44963, n44964, n44965, n44966,
         n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974,
         n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982,
         n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990,
         n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998,
         n44999, n45000, n45001, n45002, n45003, n45004, n45005, n45006,
         n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014,
         n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022,
         n45023, n45024, n45025, n45026, n45027, n45028, n45029, n45030,
         n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038,
         n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046,
         n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054,
         n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062,
         n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070,
         n45071, n45072, n45073, n45074, n45075, n45076, n45077, n45078,
         n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086,
         n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094,
         n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102,
         n45103, n45104, n45105, n45106, n45107, n45108, n45109, n45110,
         n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118,
         n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126,
         n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134,
         n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142,
         n45143, n45144, n45145, n45146, n45147, n45148, n45149, n45150,
         n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158,
         n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166,
         n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174,
         n45175, n45176, n45177, n45178, n45179, n45180, n45181, n45182,
         n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190,
         n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198,
         n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206,
         n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214,
         n45215, n45216, n45217, n45218, n45219, n45220, n45221, n45222,
         n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230,
         n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238,
         n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246,
         n45247, n45248, n45249, n45250, n45251, n45252, n45253, n45254,
         n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262,
         n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270,
         n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278,
         n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286,
         n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294,
         n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302,
         n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310,
         n45311, n45312, n45313, n45314, n45315, n45316, n45317, n45318,
         n45319, n45320, n45321, n45322, n45323, n45324, n45325, n45326,
         n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334,
         n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342,
         n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350,
         n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358,
         n45359, n45360, n45361, n45362, n45363, n45364, n45365, n45366,
         n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374,
         n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382,
         n45383, n45384, n45385, n45386, n45387, n45388, n45389, n45390,
         n45391, n45392, n45393, n45394, n45395, n45396, n45397, n45398,
         n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406,
         n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414,
         n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422,
         n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430,
         n45431, n45432, n45433, n45434, n45435, n45436, n45437, n45438,
         n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446,
         n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454,
         n45455, n45456, n45457, n45458, n45459, n45460, n45461, n45462,
         n45463, n45464, n45465, n45466, n45467, n45468, n45469, n45470,
         n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478,
         n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486,
         n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494,
         n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502,
         n45503, n45504, n45505, n45506, n45507, n45508, n45509, n45510,
         n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518,
         n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526,
         n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534,
         n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542,
         n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550,
         n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558,
         n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566,
         n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574,
         n45575, n45576, n45577, n45578, n45579, n45580, n45581, n45582,
         n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590,
         n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598,
         n45599, n45600, n45601, n45602, n45603, n45604, n45605, n45606,
         n45607, n45608, n45609, n45610, n45611, n45612, n45613, n45614,
         n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622,
         n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630,
         n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638,
         n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646,
         n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654,
         n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662,
         n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670,
         n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678,
         n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686,
         n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694,
         n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702,
         n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710,
         n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718,
         n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726,
         n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734,
         n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742,
         n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750,
         n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758,
         n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766,
         n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774,
         n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782,
         n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790,
         n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798,
         n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806,
         n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814,
         n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822,
         n45823, n45824, n45825, n45826, n45827, n45828, n45829, n45830,
         n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838,
         n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846,
         n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854,
         n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862,
         n45863, n45864, n45865, n45866, n45867, n45868, n45869, n45870,
         n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878,
         n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886,
         n45887, n45888, n45889, n45890, n45891, n45892, n45893, n45894,
         n45895, n45896, n45897, n45898, n45899, n45900, n45901, n45902,
         n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910,
         n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918,
         n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926,
         n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934,
         n45935, n45936, n45937, n45938, n45939, n45940, n45941, n45942,
         n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950,
         n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958,
         n45959, n45960, n45961, n45962, n45963, n45964, n45965, n45966,
         n45967, n45968, n45969, n45970, n45971, n45972, n45973, n45974,
         n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982,
         n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990,
         n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998,
         n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006,
         n46007, n46008, n46009, n46010, n46011, n46012, n46013, n46014,
         n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022,
         n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030,
         n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038,
         n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046,
         n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054,
         n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062,
         n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070,
         n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078,
         n46079, n46080, n46081, n46082, n46083, n46084, n46085, n46086,
         n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094,
         n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102,
         n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110,
         n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118,
         n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126,
         n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134,
         n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142,
         n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150,
         n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158,
         n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166,
         n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174,
         n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182,
         n46183, n46184, n46185, n46186, n46187, n46188, n46189, n46190,
         n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198,
         n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206,
         n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214,
         n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222,
         n46223, n46224, n46225, n46226, n46227, n46228, n46229, n46230,
         n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238,
         n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246,
         n46247, n46248, n46249, n46250, n46251, n46252, n46253, n46254,
         n46255, n46256, n46257, n46258, n46259, n46260, n46261, n46262,
         n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270,
         n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278,
         n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286,
         n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294,
         n46295, n46296, n46297, n46298, n46299, n46300, n46301, n46302,
         n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310,
         n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318,
         n46319, n46320, n46321, n46322, n46323, n46324, n46325, n46326,
         n46327, n46328, n46329, n46330, n46331, n46332, n46333, n46334,
         n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342,
         n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350,
         n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358,
         n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366,
         n46367, n46368, n46369, n46370, n46371, n46372, n46373, n46374,
         n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382,
         n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390,
         n46391, n46392, n46393, n46394, n46395, n46396, n46397, n46398,
         n46399, n46400, n46401, n46402, n46403, n46404, n46405, n46406,
         n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414,
         n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422,
         n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430,
         n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438,
         n46439, n46440, n46441, n46442, n46443, n46444, n46445, n46446,
         n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454,
         n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462,
         n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470,
         n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478,
         n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486,
         n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494,
         n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502,
         n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510,
         n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518,
         n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526,
         n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534,
         n46535, n46536, n46537, n46538, n46539, n46540, n46541, n46542,
         n46543, n46544, n46545, n46546, n46547, n46548, n46549, n46550,
         n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558,
         n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566,
         n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574,
         n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582,
         n46583, n46584, n46585, n46586, n46587, n46588, n46589, n46590,
         n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598,
         n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606,
         n46607, n46608, n46609, n46610, n46611, n46612, n46613, n46614,
         n46615, n46616, n46617, n46618, n46619, n46620, n46621, n46622,
         n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630,
         n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638,
         n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646,
         n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654,
         n46655, n46656, n46657, n46658, n46659, n46660, n46661, n46662,
         n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670,
         n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678,
         n46679, n46680, n46681, n46682, n46683, n46684, n46685, n46686,
         n46687, n46688, n46689, n46690, n46691, n46692, n46693, n46694,
         n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702,
         n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710,
         n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718,
         n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726,
         n46727, n46728, n46729, n46730, n46731, n46732, n46733, n46734,
         n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742,
         n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750,
         n46751, n46752, n46753, n46754, n46755, n46756, n46757, n46758,
         n46759, n46760, n46761, n46762, n46763, n46764, n46765, n46766,
         n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774,
         n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782,
         n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790,
         n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798,
         n46799, n46800, n46801, n46802, n46803, n46804, n46805, n46806,
         n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814,
         n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822,
         n46823, n46824, n46825, n46826, n46827, n46828, n46829, n46830,
         n46831, n46832, n46833, n46834, n46835, n46836, n46837, n46838,
         n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846,
         n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854,
         n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862,
         n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870,
         n46871, n46872, n46873, n46874, n46875, n46876, n46877, n46878,
         n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886,
         n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894,
         n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902,
         n46903, n46904, n46905, n46906, n46907, n46908, n46909, n46910,
         n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918,
         n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926,
         n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934,
         n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942,
         n46943, n46944, n46945, n46946, n46947, n46948, n46949, n46950,
         n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958,
         n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966,
         n46967, n46968, n46969, n46970, n46971, n46972, n46973, n46974,
         n46975, n46976, n46977, n46978, n46979, n46980, n46981, n46982,
         n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990,
         n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998,
         n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006,
         n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014,
         n47015, n47016, n47017, n47018, n47019, n47020, n47021, n47022,
         n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030,
         n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038,
         n47039, n47040, n47041, n47042, n47043, n47044, n47045, n47046,
         n47047, n47048, n47049, n47050, n47051, n47052, n47053, n47054,
         n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062,
         n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070,
         n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078,
         n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086,
         n47087, n47088, n47089, n47090, n47091, n47092, n47093, n47094,
         n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102,
         n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110,
         n47111, n47112, n47113, n47114, n47115, n47116, n47117, n47118,
         n47119, n47120, n47121, n47122, n47123, n47124, n47125, n47126,
         n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134,
         n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142,
         n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150,
         n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158,
         n47159, n47160, n47161, n47162, n47163, n47164, n47165, n47166,
         n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174,
         n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182,
         n47183, n47184, n47185, n47186, n47187, n47188, n47189, n47190,
         n47191, n47192, n47193, n47194, n47195, n47196, n47197, n47198,
         n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206,
         n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214,
         n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222,
         n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230,
         n47231, n47232, n47233, n47234, n47235, n47236, n47237, n47238,
         n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246,
         n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254,
         n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262,
         n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270,
         n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278,
         n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286,
         n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294,
         n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302,
         n47303, n47304, n47305, n47306, n47307, n47308, n47309, n47310,
         n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318,
         n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326,
         n47327, n47328, n47329, n47330, n47331, n47332, n47333, n47334,
         n47335, n47336, n47337, n47338, n47339, n47340, n47341, n47342,
         n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350,
         n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358,
         n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366,
         n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374,
         n47375, n47376, n47377, n47378, n47379, n47380, n47381, n47382,
         n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390,
         n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398,
         n47399, n47400, n47401, n47402, n47403, n47404, n47405, n47406,
         n47407, n47408, n47409, n47410, n47411, n47412, n47413, n47414,
         n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422,
         n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430,
         n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438,
         n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446,
         n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454,
         n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462,
         n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470,
         n47471, n47472, n47473, n47474, n47475, n47476, n47477, n47478,
         n47479, n47480, n47481, n47482, n47483, n47484, n47485, n47486,
         n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494,
         n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502,
         n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510,
         n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518,
         n47519, n47520, n47521, n47522, n47523, n47524, n47525, n47526,
         n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534,
         n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542,
         n47543, n47544, n47545, n47546, n47547, n47548, n47549, n47550,
         n47551, n47552, n47553, n47554, n47555, n47556, n47557, n47558,
         n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566,
         n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574,
         n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582,
         n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590,
         n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598,
         n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606,
         n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614,
         n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622,
         n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47630,
         n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638,
         n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646,
         n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654,
         n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662,
         n47663, n47664, n47665, n47666, n47667, n47668, n47669, n47670,
         n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678,
         n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686,
         n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47694,
         n47695, n47696, n47697, n47698, n47699, n47700, n47701, n47702,
         n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710,
         n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718,
         n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726,
         n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734,
         n47735, n47736, n47737, n47738, n47739, n47740, n47741, n47742,
         n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750,
         n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758,
         n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47766,
         n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774,
         n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782,
         n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790,
         n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798,
         n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806,
         n47807, n47808, n47809, n47810, n47811, n47812, n47813, n47814,
         n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822,
         n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830,
         n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838,
         n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846,
         n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854,
         n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862,
         n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870,
         n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878,
         n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886,
         n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894,
         n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902,
         n47903, n47904, n47905, n47906, n47907, n47908, n47909, n47910,
         n47911, n47912, n47913, n47914, n47915, n47916, n47917, n47918,
         n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926,
         n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934,
         n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942,
         n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950,
         n47951, n47952, n47953, n47954, n47955, n47956, n47957, n47958,
         n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966,
         n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974,
         n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982,
         n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990,
         n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998,
         n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006,
         n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014,
         n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022,
         n48023, n48024, n48025, n48026, n48027, n48028, n48029, n48030,
         n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038,
         n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046,
         n48047, n48048, n48049, n48050, n48051, n48052, n48053, n48054,
         n48055, n48056, n48057, n48058, n48059, n48060, n48061, n48062,
         n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070,
         n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078,
         n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086,
         n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094,
         n48095, n48096, n48097, n48098, n48099, n48100, n48101, n48102,
         n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110,
         n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118,
         n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126,
         n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134,
         n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142,
         n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150,
         n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158,
         n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166,
         n48167, n48168, n48169, n48170, n48171, n48172, n48173, n48174,
         n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182,
         n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190,
         n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198,
         n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206,
         n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214,
         n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222,
         n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230,
         n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238,
         n48239, n48240, n48241, n48242, n48243, n48244, n48245, n48246,
         n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254,
         n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262,
         n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270,
         n48271, n48272, n48273, n48274, n48275, n48276, n48277, n48278,
         n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286,
         n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294,
         n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302,
         n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310,
         n48311, n48312, n48313, n48314, n48315, n48316, n48317, n48318,
         n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326,
         n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334,
         n48335, n48336, n48337, n48338, n48339, n48340, n48341, n48342,
         n48343, n48344, n48345, n48346, n48347, n48348, n48349, n48350,
         n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358,
         n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366,
         n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374,
         n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382,
         n48383, n48384, n48385, n48386, n48387, n48388, n48389, n48390,
         n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398,
         n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406,
         n48407, n48408, n48409, n48410, n48411, n48412, n48413, n48414,
         n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422,
         n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430,
         n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438,
         n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446,
         n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454,
         n48455, n48456, n48457, n48458, n48459, n48460, n48461, n48462,
         n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470,
         n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478,
         n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486,
         n48487, n48488, n48489, n48490, n48491, n48492, n48493, n48494,
         n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502,
         n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510,
         n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518,
         n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526,
         n48527, n48528, n48529, n48530, n48531, n48532, n48533, n48534,
         n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542,
         n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550,
         n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558,
         n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566,
         n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574,
         n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582,
         n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590,
         n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598,
         n48599, n48600, n48601, n48602, n48603, n48604, n48605, n48606,
         n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614,
         n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622,
         n48623, n48624, n48625, n48626, n48627, n48628, n48629, n48630,
         n48631, n48632, n48633, n48634, n48635, n48636, n48637, n48638,
         n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646,
         n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654,
         n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662,
         n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670,
         n48671, n48672, n48673, n48674, n48675, n48676, n48677, n48678,
         n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686,
         n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694,
         n48695, n48696, n48697, n48698, n48699, n48700, n48701, n48702,
         n48703, n48704, n48705, n48706, n48707, n48708, n48709, n48710,
         n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718,
         n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726,
         n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734,
         n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742,
         n48743, n48744, n48745, n48746, n48747, n48748, n48749, n48750,
         n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758,
         n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766,
         n48767, n48768, n48769, n48770, n48771, n48772, n48773, n48774,
         n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782,
         n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790,
         n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798,
         n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806,
         n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814,
         n48815, n48816, n48817, n48818, n48819, n48820, n48821, n48822,
         n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830,
         n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838,
         n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846,
         n48847, n48848, n48849, n48850, n48851, n48852, n48853, n48854,
         n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862,
         n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870,
         n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878,
         n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886,
         n48887, n48888, n48889, n48890, n48891, n48892, n48893, n48894,
         n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902,
         n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910,
         n48911, n48912, n48913, n48914, n48915, n48916, n48917, n48918,
         n48919, n48920, n48921, n48922, n48923, n48924, n48925, n48926,
         n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934,
         n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942,
         n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950,
         n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958,
         n48959, n48960, n48961, n48962, n48963, n48964, n48965, n48966,
         n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974,
         n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982,
         n48983, n48984, n48985, n48986, n48987, n48988, n48989, n48990,
         n48991, n48992, n48993, n48994, n48995, n48996, n48997, n48998,
         n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006,
         n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014,
         n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022,
         n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030,
         n49031, n49032, n49033, n49034, n49035, n49036, n49037, n49038,
         n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046,
         n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054,
         n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062,
         n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070,
         n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078,
         n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086,
         n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094,
         n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102,
         n49103, n49104, n49105, n49106, n49107, n49108, n49109, n49110,
         n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118,
         n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126,
         n49127, n49128, n49129, n49130, n49131, n49132, n49133, n49134,
         n49135, n49136, n49137, n49138, n49139, n49140, n49141, n49142,
         n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150,
         n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158,
         n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166,
         n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174,
         n49175, n49176, n49177, n49178, n49179, n49180, n49181, n49182,
         n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190,
         n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198,
         n49199, n49200, n49201, n49202, n49203, n49204, n49205, n49206,
         n49207, n49208, n49209, n49210, n49211, n49212, n49213, n49214,
         n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222,
         n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230,
         n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238,
         n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246,
         n49247, n49248, n49249, n49250, n49251, n49252, n49253, n49254,
         n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262,
         n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270,
         n49271, n49272, n49273, n49274, n49275, n49276, n49277, n49278,
         n49279, n49280, n49281, n49282, n49283, n49284, n49285, n49286,
         n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294,
         n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302,
         n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310,
         n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318,
         n49319, n49320, n49321, n49322, n49323, n49324, n49325, n49326,
         n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334,
         n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342,
         n49343, n49344, n49345, n49346, n49347, n49348, n49349, n49350,
         n49351, n49352, n49353, n49354, n49355, n49356, n49357, n49358,
         n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366,
         n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374,
         n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382,
         n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390,
         n49391, n49392, n49393, n49394, n49395, n49396, n49397, n49398,
         n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406,
         n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414,
         n49415, n49416, n49417, n49418, n49419, n49420, n49421, n49422,
         n49423, n49424, n49425, n49426, n49427, n49428, n49429, n49430,
         n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438,
         n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446,
         n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454,
         n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462,
         n49463, n49464, n49465, n49466, n49467, n49468, n49469, n49470,
         n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478,
         n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486,
         n49487, n49488, n49489, n49490, n49491, n49492, n49493, n49494,
         n49495, n49496, n49497, n49498, n49499, n49500, n49501, n49502,
         n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510,
         n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518,
         n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526,
         n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534,
         n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542,
         n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550,
         n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558,
         n49559, n49560, n49561, n49562, n49563, n49564, n49565, n49566,
         n49567, n49568, n49569, n49570, n49571, n49572, n49573, n49574,
         n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582,
         n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590,
         n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598,
         n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606,
         n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614,
         n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622,
         n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630,
         n49631, n49632, n49633, n49634, n49635, n49636, n49637, n49638,
         n49639, n49640, n49641, n49642, n49643, n49644, n49645, n49646,
         n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654,
         n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662,
         n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670,
         n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678,
         n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686,
         n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694,
         n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702,
         n49703, n49704, n49705, n49706, n49707, n49708, n49709, n49710,
         n49711, n49712, n49713, n49714, n49715, n49716, n49717, n49718,
         n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726,
         n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734,
         n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742,
         n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750,
         n49751, n49752, n49753, n49754, n49755, n49756, n49757, n49758,
         n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766,
         n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774,
         n49775, n49776, n49777, n49778, n49779, n49780, n49781, n49782,
         n49783, n49784, n49785, n49786, n49787, n49788, n49789, n49790,
         n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798,
         n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806,
         n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814,
         n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822,
         n49823, n49824, n49825, n49826, n49827, n49828, n49829, n49830,
         n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838,
         n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846,
         n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854,
         n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862,
         n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870,
         n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878,
         n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886,
         n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894,
         n49895, n49896, n49897, n49898, n49899, n49900, n49901, n49902,
         n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910,
         n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918,
         n49919, n49920, n49921, n49922, n49923, n49924, n49925, n49926,
         n49927, n49928, n49929, n49930, n49931, n49932, n49933, n49934,
         n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942,
         n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950,
         n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958,
         n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966,
         n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974,
         n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982,
         n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990,
         n49991, n49992, n49993, n49994, n49995, n49996, n49997, n49998,
         n49999, n50000, n50001, n50002, n50003, n50004, n50005, n50006,
         n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014,
         n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022,
         n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030,
         n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038,
         n50039, n50040, n50041, n50042, n50043, n50044, n50045, n50046,
         n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054,
         n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062,
         n50063, n50064, n50065, n50066, n50067, n50068, n50069, n50070,
         n50071, n50072, n50073, n50074, n50075, n50076, n50077, n50078,
         n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086,
         n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094,
         n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102,
         n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110,
         n50111, n50112, n50113, n50114, n50115, n50116, n50117, n50118,
         n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126,
         n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134,
         n50135, n50136, n50137, n50138, n50139, n50140, n50141, n50142,
         n50143, n50144, n50145, n50146, n50147, n50148, n50149, n50150,
         n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158,
         n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166,
         n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174,
         n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182,
         n50183, n50184, n50185, n50186, n50187, n50188, n50189, n50190,
         n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198,
         n50199, n50200, n50201, n50202, n50203, n50204, n50205, n50206,
         n50207, n50208, n50209, n50210, n50211, n50212, n50213, n50214,
         n50215, n50216, n50217, n50218, n50219, n50220, n50221, n50222,
         n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230,
         n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238,
         n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246,
         n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254,
         n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262,
         n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270,
         n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278,
         n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286,
         n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294,
         n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302,
         n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310,
         n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318,
         n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326,
         n50327, n50328, n50329, n50330, n50331, n50332, n50333, n50334,
         n50335, n50336, n50337, n50338, n50339, n50340, n50341, n50342,
         n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350,
         n50351, n50352, n50353, n50354, n50355, n50356, n50357, n50358,
         n50359, n50360, n50361, n50362, n50363, n50364, n50365, n50366,
         n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374,
         n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382,
         n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390,
         n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398,
         n50399, n50400, n50401, n50402, n50403, n50404, n50405, n50406,
         n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414,
         n50415, n50416, n50417, n50418, n50419, n50420, n50421, n50422,
         n50423, n50424, n50425, n50426, n50427, n50428, n50429, n50430,
         n50431, n50432, n50433, n50434, n50435, n50436, n50437, n50438,
         n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446,
         n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454,
         n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462,
         n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470,
         n50471, n50472, n50473, n50474, n50475, n50476, n50477, n50478,
         n50479, n50480, n50481, n50482, n50483, n50484, n50485, n50486,
         n50487, n50488, n50489, n50490, n50491, n50492, n50493, n50494,
         n50495, n50496, n50497, n50498, n50499, n50500, n50501, n50502,
         n50503, n50504, n50505, n50506, n50507, n50508, n50509, n50510,
         n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518,
         n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526,
         n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534,
         n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542,
         n50543, n50544, n50545, n50546, n50547, n50548, n50549, n50550,
         n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558,
         n50559, n50560, n50561, n50562, n50563, n50564, n50565, n50566,
         n50567, n50568, n50569, n50570, n50571, n50572, n50573, n50574,
         n50575, n50576, n50577, n50578, n50579, n50580, n50581, n50582,
         n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590,
         n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598,
         n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606,
         n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614,
         n50615, n50616, n50617, n50618, n50619, n50620, n50621, n50622,
         n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630,
         n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638,
         n50639, n50640, n50641, n50642, n50643, n50644, n50645, n50646,
         n50647, n50648, n50649, n50650, n50651, n50652, n50653, n50654,
         n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662,
         n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670,
         n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678,
         n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686,
         n50687, n50688, n50689, n50690, n50691, n50692, n50693, n50694,
         n50695, n50696, n50697, n50698, n50699, n50700, n50701, n50702,
         n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710,
         n50711, n50712, n50713, n50714, n50715, n50716, n50717, n50718,
         n50719, n50720, n50721, n50722, n50723, n50724, n50725, n50726,
         n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734,
         n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742,
         n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750,
         n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758,
         n50759, n50760, n50761, n50762, n50763, n50764, n50765, n50766,
         n50767, n50768, n50769, n50770, n50771, n50772, n50773, n50774,
         n50775, n50776, n50777, n50778, n50779, n50780, n50781, n50782,
         n50783, n50784, n50785, n50786, n50787, n50788, n50789, n50790,
         n50791, n50792, n50793, n50794, n50795, n50796, n50797, n50798,
         n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806,
         n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814,
         n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822,
         n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830,
         n50831, n50832, n50833, n50834, n50835, n50836, n50837, n50838,
         n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846,
         n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854,
         n50855, n50856, n50857, n50858, n50859, n50860, n50861, n50862,
         n50863, n50864, n50865, n50866, n50867, n50868, n50869, n50870,
         n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878,
         n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886,
         n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894,
         n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902,
         n50903, n50904, n50905, n50906, n50907, n50908, n50909, n50910,
         n50911, n50912, n50913, n50914, n50915, n50916, n50917, n50918,
         n50919, n50920, n50921, n50922, n50923, n50924, n50925, n50926,
         n50927, n50928, n50929, n50930, n50931, n50932, n50933, n50934,
         n50935, n50936, n50937, n50938, n50939, n50940, n50941, n50942,
         n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950,
         n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958,
         n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966,
         n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974,
         n50975, n50976, n50977, n50978, n50979, n50980, n50981, n50982,
         n50983, n50984, n50985, n50986, n50987, n50988, n50989, n50990,
         n50991, n50992, n50993, n50994, n50995, n50996, n50997, n50998,
         n50999, n51000, n51001, n51002, n51003, n51004, n51005, n51006,
         n51007, n51008, n51009, n51010, n51011, n51012, n51013, n51014,
         n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022,
         n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030,
         n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038,
         n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046,
         n51047, n51048, n51049, n51050, n51051, n51052, n51053, n51054,
         n51055, n51056, n51057, n51058, n51059, n51060, n51061, n51062,
         n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070,
         n51071, n51072, n51073, n51074, n51075, n51076, n51077, n51078,
         n51079, n51080, n51081, n51082, n51083, n51084, n51085, n51086,
         n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094,
         n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102,
         n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110,
         n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118,
         n51119, n51120, n51121, n51122, n51123, n51124, n51125, n51126,
         n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51134,
         n51135, n51136, n51137, n51138, n51139, n51140, n51141, n51142,
         n51143, n51144, n51145, n51146, n51147, n51148, n51149, n51150,
         n51151, n51152, n51153, n51154, n51155, n51156, n51157, n51158,
         n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166,
         n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174,
         n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182,
         n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190,
         n51191, n51192, n51193, n51194, n51195, n51196, n51197, n51198,
         n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206,
         n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214,
         n51215, n51216, n51217, n51218, n51219, n51220, n51221, n51222,
         n51223, n51224, n51225, n51226, n51227, n51228, n51229, n51230,
         n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238,
         n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246,
         n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254,
         n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262,
         n51263, n51264, n51265, n51266, n51267, n51268, n51269, n51270,
         n51271, n51272, n51273, n51274, n51275, n51276, n51277, n51278,
         n51279, n51280, n51281, n51282, n51283, n51284, n51285, n51286,
         n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294,
         n51295, n51296, n51297, n51298, n51299, n51300, n51301, n51302,
         n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310,
         n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318,
         n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326,
         n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334,
         n51335, n51336, n51337, n51338, n51339, n51340, n51341, n51342,
         n51343, n51344, n51345, n51346, n51347, n51348, n51349, n51350,
         n51351, n51352, n51353, n51354, n51355, n51356, n51357, n51358,
         n51359, n51360, n51361, n51362, n51363, n51364, n51365, n51366,
         n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374,
         n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382,
         n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390,
         n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398,
         n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406,
         n51407, n51408, n51409, n51410, n51411, n51412, n51413, n51414,
         n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422,
         n51423, n51424, n51425, n51426, n51427, n51428, n51429, n51430,
         n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438;
  wire   [1:0] state;
  wire   [1:0] nxt_state;
  wire   [3:0] nxt_data_num;

  LZSS_DW01_inc_0 add_203 ( .A({n37194, n37191, n37192, n37193, n37187, n37188,
        n37189, n37190, n37184, n37185, n37186, n36933}), .SUM({N23562, N23561,
        N23560, N23559, N23558, N23557, N23556, N23555, N23554, N23553, N23552,
        N23551}) );
  DFFRX1 dict_reg_75__4_ ( .D(n35129), .CK(clk), .RN(n42401), .QN(n33004) );
  DFFRX1 dict_reg_76__4_ ( .D(n35137), .CK(clk), .RN(n42401), .QN(n33012) );
  DFFRX1 dict_reg_74__7_ ( .D(n35118), .CK(clk), .RN(n42339), .Q(n37245), .QN(
        n32993) );
  DFFRX1 dict_reg_75__7_ ( .D(n35126), .CK(clk), .RN(n42339), .Q(n36925), .QN(
        n33001) );
  DFFRX1 dict_reg_76__7_ ( .D(n35134), .CK(clk), .RN(n42339), .Q(n37020), .QN(
        n33009) );
  DFFRX1 dict_reg_73__7_ ( .D(n35110), .CK(clk), .RN(n42339), .Q(n36946), .QN(
        n32985) );
  DFFRX1 dict_reg_77__4_ ( .D(n35145), .CK(clk), .RN(n42401), .QN(n33020) );
  DFFRX1 dict_reg_78__4_ ( .D(n35153), .CK(clk), .RN(n42401), .QN(n33028) );
  DFFRX1 dict_reg_77__7_ ( .D(n35142), .CK(clk), .RN(n42339), .Q(n37244), .QN(
        n33017) );
  DFFRX1 dict_reg_78__7_ ( .D(n35150), .CK(clk), .RN(n42339), .Q(n36931), .QN(
        n33025) );
  DFFRX1 dict_reg_84__7_ ( .D(n35198), .CK(clk), .RN(n42340), .Q(n37243), .QN(
        n33073) );
  DFFRX1 dict_reg_85__7_ ( .D(n35206), .CK(clk), .RN(n42340), .Q(n50456), .QN(
        n33081) );
  DFFRX1 dict_reg_88__7_ ( .D(n35230), .CK(clk), .RN(n42340), .Q(n50459), .QN(
        n33105) );
  DFFRX1 dict_reg_81__4_ ( .D(n35177), .CK(clk), .RN(n42401), .Q(n37242), .QN(
        n33052) );
  DFFRX1 dict_reg_82__7_ ( .D(n35182), .CK(clk), .RN(n42339), .Q(n36930), .QN(
        n33057) );
  DFFRX1 dict_reg_83__7_ ( .D(n35190), .CK(clk), .RN(n42339), .Q(n37019), .QN(
        n33065) );
  DFFRX1 dict_reg_86__7_ ( .D(n35214), .CK(clk), .RN(n42340), .Q(n50457), .QN(
        n33089) );
  DFFRX1 dict_reg_87__7_ ( .D(n35222), .CK(clk), .RN(n42340), .Q(n50458), .QN(
        n33097) );
  DFFRX1 dict_reg_89__7_ ( .D(n35238), .CK(clk), .RN(n42340), .Q(n50460), .QN(
        n33113) );
  DFFRX1 dict_reg_90__7_ ( .D(n35246), .CK(clk), .RN(n42340), .Q(n50461), .QN(
        n33121) );
  DFFRX1 dict_reg_91__7_ ( .D(n35254), .CK(clk), .RN(n42340), .Q(n50462), .QN(
        n33129) );
  DFFRX1 dict_reg_93__7_ ( .D(n35270), .CK(clk), .RN(n42340), .Q(n50464), .QN(
        n33145) );
  DFFRX1 dict_reg_92__7_ ( .D(n35262), .CK(clk), .RN(n42340), .Q(n50463), .QN(
        n33137) );
  DFFRX1 dict_reg_249__1_ ( .D(n36524), .CK(clk), .RN(n42374), .Q(n37200),
        .QN(n34399) );
  DFFRX1 dict_reg_94__7_ ( .D(n35278), .CK(clk), .RN(n42340), .Q(n50465), .QN(
        n33153) );
  DFFRX1 dict_reg_116__7_ ( .D(n35454), .CK(clk), .RN(n42341), .Q(n50487),
        .QN(n33329) );
  DFFRX1 dict_reg_117__7_ ( .D(n35462), .CK(clk), .RN(n42341), .Q(n37252),
        .QN(n33337) );
  DFFRX1 dict_reg_120__7_ ( .D(n35486), .CK(clk), .RN(n42342), .Q(n50490),
        .QN(n33361) );
  DFFRX1 dict_reg_121__7_ ( .D(n35494), .CK(clk), .RN(n42342), .Q(n50491),
        .QN(n33369) );
  DFFRX1 dict_reg_119__7_ ( .D(n35478), .CK(clk), .RN(n42341), .Q(n50489),
        .QN(n33353) );
  DFFRX1 dict_reg_114__7_ ( .D(n35438), .CK(clk), .RN(n42341), .Q(n50485),
        .QN(n33313) );
  DFFRX1 dict_reg_199__4_ ( .D(n36121), .CK(clk), .RN(n42410), .QN(n33996) );
  DFFRX1 dict_reg_200__4_ ( .D(n36129), .CK(clk), .RN(n42410), .QN(n34004) );
  DFFRX1 dict_reg_122__4_ ( .D(n35505), .CK(clk), .RN(n42404), .QN(n33380) );
  DFFRX1 dict_reg_123__4_ ( .D(n35513), .CK(clk), .RN(n42404), .QN(n33388) );
  DFFRX1 dict_reg_122__7_ ( .D(n35502), .CK(clk), .RN(n42342), .Q(n50492),
        .QN(n33377) );
  DFFRX1 dict_reg_123__7_ ( .D(n35510), .CK(clk), .RN(n42342), .Q(n50493),
        .QN(n33385) );
  DFFRX1 dict_reg_124__7_ ( .D(n35518), .CK(clk), .RN(n42342), .Q(n50494),
        .QN(n33393) );
  DFFRX1 dict_reg_125__7_ ( .D(n35526), .CK(clk), .RN(n42342), .Q(n37251),
        .QN(n33401) );
  DFFRX1 dict_reg_216__6_ ( .D(n36255), .CK(clk), .RN(n37595), .Q(n37195),
        .QN(n34130) );
  DFFRX1 dict_reg_251__6_ ( .D(n36535), .CK(clk), .RN(n42338), .Q(n37553),
        .QN(n34410) );
  DFFRX1 dict_reg_216__7_ ( .D(n36254), .CK(clk), .RN(n42349), .Q(n37543),
        .QN(n34129) );
  DFFRX1 dict_reg_217__7_ ( .D(n36262), .CK(clk), .RN(n42349), .Q(n37542),
        .QN(n34137) );
  DFFRX1 dict_reg_251__7_ ( .D(n36534), .CK(clk), .RN(n37594), .Q(n37552),
        .QN(n34409) );
  DFFRX1 dict_reg_216__0_ ( .D(n36261), .CK(clk), .RN(n42362), .Q(n37541),
        .QN(n34136) );
  DFFRX1 dict_reg_216__2_ ( .D(n36259), .CK(clk), .RN(n42387), .Q(n37548),
        .QN(n34134) );
  DFFRX1 dict_reg_217__2_ ( .D(n36267), .CK(clk), .RN(n42387), .Q(n37547),
        .QN(n34142) );
  DFFRX1 dict_reg_251__2_ ( .D(n36539), .CK(clk), .RN(n42388), .Q(n37550),
        .QN(n34414) );
  DFFRX1 dict_reg_216__3_ ( .D(n36258), .CK(clk), .RN(n42399), .Q(n37546),
        .QN(n34133) );
  DFFRX1 dict_reg_217__3_ ( .D(n36266), .CK(clk), .RN(n42399), .Q(n37545),
        .QN(n34141) );
  DFFRX1 dict_reg_251__3_ ( .D(n36538), .CK(clk), .RN(n42400), .Q(n37549),
        .QN(n34413) );
  DFFRX1 dict_reg_216__4_ ( .D(n36257), .CK(clk), .RN(n37595), .Q(n37544),
        .QN(n34132) );
  DFFRX1 dict_reg_251__4_ ( .D(n36537), .CK(clk), .RN(n42412), .Q(n37554),
        .QN(n34412) );
  DFFRX1 dict_reg_254__7_ ( .D(n36558), .CK(clk), .RN(n37596), .QN(n9659) );
  DFFRX1 dict_reg_254__3_ ( .D(n36562), .CK(clk), .RN(n42400), .QN(n9667) );
  DFFRX1 dict_reg_254__4_ ( .D(n36561), .CK(clk), .RN(n42412), .QN(n9669) );
  DFFRX1 dict_reg_254__5_ ( .D(n36560), .CK(clk), .RN(n42337), .QN(n9655) );
  DFFRX1 dict_reg_254__2_ ( .D(n36563), .CK(clk), .RN(n42388), .QN(n9665) );
  DFFRX1 dict_reg_214__3_ ( .D(n36242), .CK(clk), .RN(n42399), .Q(n49516),
        .QN(n34117) );
  DFFRX1 dict_reg_214__0_ ( .D(n36245), .CK(clk), .RN(n42362), .QN(n34120) );
  DFFRX1 dict_reg_212__4_ ( .D(n36225), .CK(clk), .RN(n42411), .Q(n37540),
        .QN(n34100) );
  DFFRX1 dict_reg_157__4_ ( .D(n35785), .CK(clk), .RN(n42407), .QN(n33660) );
  DFFRX1 dict_reg_168__4_ ( .D(n35873), .CK(clk), .RN(n42408), .QN(n33748) );
  DFFRX1 dict_reg_171__4_ ( .D(n35897), .CK(clk), .RN(n42408), .QN(n33772) );
  DFFRX1 dict_reg_172__4_ ( .D(n35905), .CK(clk), .RN(n42408), .QN(n33780) );
  DFFRX1 dict_reg_178__4_ ( .D(n35953), .CK(clk), .RN(n42408), .QN(n33828) );
  DFFRX1 dict_reg_184__4_ ( .D(n36001), .CK(clk), .RN(n42409), .QN(n33876) );
  DFFRX1 dict_reg_201__4_ ( .D(n36137), .CK(clk), .RN(n42410), .QN(n34012) );
  DFFRX1 dict_reg_211__4_ ( .D(n36217), .CK(clk), .RN(n42411), .QN(n34092) );
  DFFRX1 dict_reg_186__4_ ( .D(n36017), .CK(clk), .RN(n42409), .QN(n33892) );
  DFFRX1 dict_reg_155__4_ ( .D(n35769), .CK(clk), .RN(n42407), .QN(n33644) );
  DFFRX1 dict_reg_187__4_ ( .D(n36025), .CK(clk), .RN(n42409), .QN(n33900) );
  DFFRX1 dict_reg_150__4_ ( .D(n35729), .CK(clk), .RN(n42406), .QN(n33604) );
  DFFRX1 dict_reg_189__4_ ( .D(n36041), .CK(clk), .RN(n42409), .QN(n33916) );
  DFFRX1 dict_reg_188__4_ ( .D(n36033), .CK(clk), .RN(n42409), .QN(n33908) );
  DFFRX1 dict_reg_111__5_ ( .D(n35416), .CK(clk), .RN(n42325), .QN(n33291) );
  DFFRX1 dict_reg_112__5_ ( .D(n35424), .CK(clk), .RN(n42325), .QN(n33299) );
  DFFRX1 dict_reg_111__1_ ( .D(n35420), .CK(clk), .RN(n42363), .QN(n33295) );
  DFFRX1 dict_reg_112__1_ ( .D(n35428), .CK(clk), .RN(n42363), .QN(n33303) );
  DFFRX1 dict_reg_113__5_ ( .D(n35432), .CK(clk), .RN(n42325), .QN(n33307) );
  DFFRX1 dict_reg_114__5_ ( .D(n35440), .CK(clk), .RN(n42325), .QN(n33315) );
  DFFRX1 dict_reg_115__5_ ( .D(n35448), .CK(clk), .RN(n42325), .QN(n33323) );
  DFFRX1 dict_reg_119__5_ ( .D(n35480), .CK(clk), .RN(n42325), .QN(n33355) );
  DFFRX1 dict_reg_120__5_ ( .D(n35488), .CK(clk), .RN(n42325), .QN(n33363) );
  DFFRX1 dict_reg_121__5_ ( .D(n35496), .CK(clk), .RN(n42325), .QN(n33371) );
  DFFRX1 dict_reg_122__5_ ( .D(n35504), .CK(clk), .RN(n42326), .QN(n33379) );
  DFFRX1 dict_reg_123__5_ ( .D(n35512), .CK(clk), .RN(n42326), .QN(n33387) );
  DFFRX1 dict_reg_124__5_ ( .D(n35520), .CK(clk), .RN(n42326), .QN(n33395) );
  DFFRX1 dict_reg_127__5_ ( .D(n35544), .CK(clk), .RN(n42326), .QN(n33419) );
  DFFRX1 dict_reg_128__5_ ( .D(n35552), .CK(clk), .RN(n42326), .QN(n33427) );
  DFFRX1 dict_reg_131__5_ ( .D(n35576), .CK(clk), .RN(n42326), .QN(n33451) );
  DFFRX1 dict_reg_113__1_ ( .D(n35436), .CK(clk), .RN(n42363), .QN(n33311) );
  DFFRX1 dict_reg_119__1_ ( .D(n35484), .CK(clk), .RN(n42363), .QN(n33359) );
  DFFRX1 dict_reg_120__1_ ( .D(n35492), .CK(clk), .RN(n42363), .QN(n33367) );
  DFFRX1 dict_reg_121__1_ ( .D(n35500), .CK(clk), .RN(n42363), .QN(n33375) );
  DFFRX1 dict_reg_122__1_ ( .D(n35508), .CK(clk), .RN(n42364), .QN(n33383) );
  DFFRX1 dict_reg_123__1_ ( .D(n35516), .CK(clk), .RN(n42364), .QN(n33391) );
  DFFRX1 dict_reg_124__1_ ( .D(n35524), .CK(clk), .RN(n42364), .QN(n33399) );
  DFFRX1 dict_reg_127__1_ ( .D(n35548), .CK(clk), .RN(n42364), .QN(n33423) );
  DFFRX1 dict_reg_128__1_ ( .D(n35556), .CK(clk), .RN(n42364), .QN(n33431) );
  DFFRX1 dict_reg_131__1_ ( .D(n35580), .CK(clk), .RN(n42364), .QN(n33455) );
  DFFRX1 dict_reg_129__5_ ( .D(n35560), .CK(clk), .RN(n42326), .QN(n33435) );
  DFFRX1 dict_reg_130__5_ ( .D(n35568), .CK(clk), .RN(n42326), .QN(n33443) );
  DFFRX1 dict_reg_135__5_ ( .D(n35608), .CK(clk), .RN(n42327), .QN(n33483) );
  DFFRX1 dict_reg_139__5_ ( .D(n35640), .CK(clk), .RN(n42327), .QN(n33515) );
  DFFRX1 dict_reg_146__5_ ( .D(n35696), .CK(clk), .RN(n42328), .QN(n33571) );
  DFFRX1 dict_reg_152__5_ ( .D(n35744), .CK(clk), .RN(n42328), .QN(n33619) );
  DFFRX1 dict_reg_153__5_ ( .D(n35752), .CK(clk), .RN(n42328), .QN(n33627) );
  DFFRX1 dict_reg_154__5_ ( .D(n35760), .CK(clk), .RN(n42328), .Q(n37247),
        .QN(n33635) );
  DFFRX1 dict_reg_155__5_ ( .D(n35768), .CK(clk), .RN(n42328), .QN(n33643) );
  DFFRX1 dict_reg_156__5_ ( .D(n35776), .CK(clk), .RN(n42328), .QN(n33651) );
  DFFRX1 dict_reg_157__5_ ( .D(n35784), .CK(clk), .RN(n42328), .QN(n33659) );
  DFFRX1 dict_reg_158__5_ ( .D(n35792), .CK(clk), .RN(n42329), .QN(n33667) );
  DFFRX1 dict_reg_159__5_ ( .D(n35800), .CK(clk), .RN(n42329), .QN(n33675) );
  DFFRX1 dict_reg_160__5_ ( .D(n35808), .CK(clk), .RN(n42329), .QN(n33683) );
  DFFRX1 dict_reg_161__5_ ( .D(n35816), .CK(clk), .RN(n42329), .QN(n33691) );
  DFFRX1 dict_reg_162__5_ ( .D(n35824), .CK(clk), .RN(n42329), .QN(n33699) );
  DFFRX1 dict_reg_163__5_ ( .D(n35832), .CK(clk), .RN(n42329), .QN(n33707) );
  DFFRX1 dict_reg_172__5_ ( .D(n35904), .CK(clk), .RN(n42330), .QN(n33779) );
  DFFRX1 dict_reg_173__5_ ( .D(n35912), .CK(clk), .RN(n42330), .QN(n33787) );
  DFFRX1 dict_reg_175__5_ ( .D(n35928), .CK(clk), .RN(n42330), .QN(n33803) );
  DFFRX1 dict_reg_190__5_ ( .D(n36048), .CK(clk), .RN(n42331), .QN(n33923) );
  DFFRX1 dict_reg_191__5_ ( .D(n36056), .CK(clk), .RN(n42331), .QN(n33931) );
  DFFRX1 dict_reg_194__5_ ( .D(n36080), .CK(clk), .RN(n42332), .QN(n33955) );
  DFFRX1 dict_reg_195__5_ ( .D(n36088), .CK(clk), .RN(n42332), .QN(n33963) );
  DFFRX1 dict_reg_196__5_ ( .D(n36096), .CK(clk), .RN(n42332), .QN(n33971) );
  DFFRX1 dict_reg_197__5_ ( .D(n36104), .CK(clk), .RN(n42332), .QN(n33979) );
  DFFRX1 dict_reg_198__5_ ( .D(n36112), .CK(clk), .RN(n42332), .QN(n33987) );
  DFFRX1 dict_reg_199__5_ ( .D(n36120), .CK(clk), .RN(n42332), .QN(n33995) );
  DFFRX1 dict_reg_210__5_ ( .D(n36208), .CK(clk), .RN(n42333), .QN(n34083) );
  DFFRX1 dict_reg_220__5_ ( .D(n36288), .CK(clk), .RN(n42334), .QN(n34163) );
  DFFRX1 dict_reg_129__1_ ( .D(n35564), .CK(clk), .RN(n42364), .QN(n33439) );
  DFFRX1 dict_reg_130__1_ ( .D(n35572), .CK(clk), .RN(n42364), .QN(n33447) );
  DFFRX1 dict_reg_135__1_ ( .D(n35612), .CK(clk), .RN(n42365), .QN(n33487) );
  DFFRX1 dict_reg_139__1_ ( .D(n35644), .CK(clk), .RN(n42365), .QN(n33519) );
  DFFRX1 dict_reg_152__1_ ( .D(n35748), .CK(clk), .RN(n42366), .QN(n33623) );
  DFFRX1 dict_reg_153__1_ ( .D(n35756), .CK(clk), .RN(n42366), .QN(n33631) );
  DFFRX1 dict_reg_156__1_ ( .D(n35780), .CK(clk), .RN(n42366), .QN(n33655) );
  DFFRX1 dict_reg_157__1_ ( .D(n35788), .CK(clk), .RN(n42366), .QN(n33663) );
  DFFRX1 dict_reg_158__1_ ( .D(n35796), .CK(clk), .RN(n42367), .QN(n33671) );
  DFFRX1 dict_reg_159__1_ ( .D(n35804), .CK(clk), .RN(n42367), .QN(n33679) );
  DFFRX1 dict_reg_160__1_ ( .D(n35812), .CK(clk), .RN(n42367), .QN(n33687) );
  DFFRX1 dict_reg_161__1_ ( .D(n35820), .CK(clk), .RN(n42367), .QN(n33695) );
  DFFRX1 dict_reg_162__1_ ( .D(n35828), .CK(clk), .RN(n42367), .QN(n33703) );
  DFFRX1 dict_reg_163__1_ ( .D(n35836), .CK(clk), .RN(n42367), .QN(n33711) );
  DFFRX1 dict_reg_172__1_ ( .D(n35908), .CK(clk), .RN(n42368), .QN(n33783) );
  DFFRX1 dict_reg_191__1_ ( .D(n36060), .CK(clk), .RN(n42369), .QN(n33935) );
  DFFRX1 dict_reg_198__1_ ( .D(n36116), .CK(clk), .RN(n42370), .QN(n33991) );
  DFFRX1 dict_reg_212__1_ ( .D(n36228), .CK(clk), .RN(n42371), .QN(n34103) );
  DFFRX1 dict_reg_200__5_ ( .D(n36128), .CK(clk), .RN(n42332), .QN(n34003) );
  DFFRX1 dict_reg_207__5_ ( .D(n36184), .CK(clk), .RN(n42333), .QN(n34059) );
  DFFRX1 dict_reg_200__1_ ( .D(n36132), .CK(clk), .RN(n42370), .QN(n34007) );
  DFFRX1 dict_reg_207__1_ ( .D(n36188), .CK(clk), .RN(n42371), .QN(n34063) );
  DFFRX1 dict_reg_132__5_ ( .D(n35584), .CK(clk), .RN(n42326), .QN(n33459) );
  DFFRX1 dict_reg_133__5_ ( .D(n35592), .CK(clk), .RN(n42326), .QN(n33467) );
  DFFRX1 dict_reg_134__5_ ( .D(n35600), .CK(clk), .RN(n42327), .QN(n33475) );
  DFFRX1 dict_reg_136__5_ ( .D(n35616), .CK(clk), .RN(n42327), .QN(n33491) );
  DFFRX1 dict_reg_137__5_ ( .D(n35624), .CK(clk), .RN(n42327), .QN(n33499) );
  DFFRX1 dict_reg_140__5_ ( .D(n35648), .CK(clk), .RN(n42327), .QN(n33523) );
  DFFRX1 dict_reg_141__5_ ( .D(n35656), .CK(clk), .RN(n42327), .QN(n33531) );
  DFFRX1 dict_reg_143__5_ ( .D(n35672), .CK(clk), .RN(n42327), .QN(n33547) );
  DFFRX1 dict_reg_164__5_ ( .D(n35840), .CK(clk), .RN(n42329), .QN(n33715) );
  DFFRX1 dict_reg_165__5_ ( .D(n35848), .CK(clk), .RN(n42329), .QN(n33723) );
  DFFRX1 dict_reg_166__5_ ( .D(n35856), .CK(clk), .RN(n42329), .QN(n33731) );
  DFFRX1 dict_reg_176__5_ ( .D(n35936), .CK(clk), .RN(n42330), .QN(n33811) );
  DFFRX1 dict_reg_178__5_ ( .D(n35952), .CK(clk), .RN(n42330), .QN(n33827) );
  DFFRX1 dict_reg_179__5_ ( .D(n35960), .CK(clk), .RN(n42330), .QN(n33835) );
  DFFRX1 dict_reg_180__5_ ( .D(n35968), .CK(clk), .RN(n42330), .QN(n33843) );
  DFFRX1 dict_reg_181__5_ ( .D(n35976), .CK(clk), .RN(n42330), .QN(n33851) );
  DFFRX1 dict_reg_182__5_ ( .D(n35984), .CK(clk), .RN(n42331), .QN(n33859) );
  DFFRX1 dict_reg_183__5_ ( .D(n35992), .CK(clk), .RN(n42331), .QN(n33867) );
  DFFRX1 dict_reg_184__5_ ( .D(n36000), .CK(clk), .RN(n42331), .QN(n33875) );
  DFFRX1 dict_reg_208__5_ ( .D(n36192), .CK(clk), .RN(n42333), .QN(n34067) );
  DFFRX1 dict_reg_209__5_ ( .D(n36200), .CK(clk), .RN(n42333), .QN(n34075) );
  DFFRX1 dict_reg_132__1_ ( .D(n35588), .CK(clk), .RN(n42364), .QN(n33463) );
  DFFRX1 dict_reg_133__1_ ( .D(n35596), .CK(clk), .RN(n42364), .QN(n33471) );
  DFFRX1 dict_reg_134__1_ ( .D(n35604), .CK(clk), .RN(n42365), .QN(n33479) );
  DFFRX1 dict_reg_140__1_ ( .D(n35652), .CK(clk), .RN(n42365), .QN(n33527) );
  DFFRX1 dict_reg_141__1_ ( .D(n35660), .CK(clk), .RN(n42365), .QN(n33535) );
  DFFRX1 dict_reg_164__1_ ( .D(n35844), .CK(clk), .RN(n42367), .QN(n33719) );
  DFFRX1 dict_reg_165__1_ ( .D(n35852), .CK(clk), .RN(n42367), .QN(n33727) );
  DFFRX1 dict_reg_166__1_ ( .D(n35860), .CK(clk), .RN(n42367), .QN(n33735) );
  DFFRX1 dict_reg_183__1_ ( .D(n35996), .CK(clk), .RN(n42369), .QN(n33871) );
  DFFRX1 dict_reg_208__1_ ( .D(n36196), .CK(clk), .RN(n42371), .QN(n34071) );
  DFFRX1 dict_reg_209__1_ ( .D(n36204), .CK(clk), .RN(n42371), .QN(n34079) );
  DFFRX1 dict_reg_144__5_ ( .D(n35680), .CK(clk), .RN(n42327), .QN(n33555) );
  DFFRX1 dict_reg_145__5_ ( .D(n35688), .CK(clk), .RN(n42327), .QN(n33563) );
  DFFRX1 dict_reg_147__5_ ( .D(n35704), .CK(clk), .RN(n42328), .QN(n33579) );
  DFFRX1 dict_reg_148__5_ ( .D(n35712), .CK(clk), .RN(n42328), .QN(n33587) );
  DFFRX1 dict_reg_149__5_ ( .D(n35720), .CK(clk), .RN(n42328), .QN(n33595) );
  DFFRX1 dict_reg_188__5_ ( .D(n36032), .CK(clk), .RN(n42331), .QN(n33907) );
  DFFRX1 dict_reg_189__5_ ( .D(n36040), .CK(clk), .RN(n42331), .QN(n33915) );
  DFFRX1 dict_reg_192__5_ ( .D(n36064), .CK(clk), .RN(n42331), .QN(n33939) );
  DFFRX1 dict_reg_202__5_ ( .D(n36144), .CK(clk), .RN(n42332), .QN(n34019) );
  DFFRX1 dict_reg_203__5_ ( .D(n36152), .CK(clk), .RN(n42332), .QN(n34027) );
  DFFRX1 dict_reg_205__5_ ( .D(n36168), .CK(clk), .RN(n42332), .QN(n34043) );
  DFFRX1 dict_reg_206__5_ ( .D(n36176), .CK(clk), .RN(n42333), .QN(n34051) );
  DFFRX1 dict_reg_213__5_ ( .D(n36232), .CK(clk), .RN(n42333), .QN(n34107) );
  DFFRX1 dict_reg_214__5_ ( .D(n36240), .CK(clk), .RN(n42333), .QN(n34115) );
  DFFRX1 dict_reg_215__5_ ( .D(n36248), .CK(clk), .RN(n42333), .QN(n34123) );
  DFFRX1 dict_reg_216__5_ ( .D(n36256), .CK(clk), .RN(n42333), .QN(n34131) );
  DFFRX1 dict_reg_217__5_ ( .D(n36264), .CK(clk), .RN(n42333), .QN(n34139) );
  DFFRX1 dict_reg_218__5_ ( .D(n36272), .CK(clk), .RN(n42334), .QN(n34147) );
  DFFRX1 dict_reg_219__5_ ( .D(n36280), .CK(clk), .RN(n42334), .QN(n34155) );
  DFFRX1 dict_reg_221__5_ ( .D(n36296), .CK(clk), .RN(n42334), .QN(n34171) );
  DFFRX1 dict_reg_222__5_ ( .D(n36304), .CK(clk), .RN(n42334), .QN(n34179) );
  DFFRX1 dict_reg_223__5_ ( .D(n36312), .CK(clk), .RN(n42334), .QN(n34187) );
  DFFRX1 dict_reg_224__5_ ( .D(n36320), .CK(clk), .RN(n42334), .QN(n34195) );
  DFFRX1 dict_reg_225__5_ ( .D(n36328), .CK(clk), .RN(n42334), .QN(n34203) );
  DFFRX1 dict_reg_226__5_ ( .D(n36336), .CK(clk), .RN(n42334), .QN(n34211) );
  DFFRX1 dict_reg_227__5_ ( .D(n36344), .CK(clk), .RN(n42334), .QN(n34219) );
  DFFRX1 dict_reg_228__5_ ( .D(n36352), .CK(clk), .RN(n42334), .QN(n34227) );
  DFFRX1 dict_reg_229__5_ ( .D(n36360), .CK(clk), .RN(n42334), .QN(n34235) );
  DFFRX1 dict_reg_230__5_ ( .D(n36368), .CK(clk), .RN(n42335), .QN(n34243) );
  DFFRX1 dict_reg_231__5_ ( .D(n36376), .CK(clk), .RN(n42335), .QN(n34251) );
  DFFRX1 dict_reg_232__5_ ( .D(n36384), .CK(clk), .RN(n42335), .QN(n34259) );
  DFFRX1 dict_reg_233__5_ ( .D(n36392), .CK(clk), .RN(n42335), .QN(n34267) );
  DFFRX1 dict_reg_234__5_ ( .D(n36400), .CK(clk), .RN(n42335), .QN(n34275) );
  DFFRX1 dict_reg_235__5_ ( .D(n36408), .CK(clk), .RN(n42335), .QN(n34283) );
  DFFRX1 dict_reg_236__5_ ( .D(n36416), .CK(clk), .RN(n42335), .QN(n34291) );
  DFFRX1 dict_reg_237__5_ ( .D(n36424), .CK(clk), .RN(n42335), .QN(n34299) );
  DFFRX1 dict_reg_238__5_ ( .D(n36432), .CK(clk), .RN(n42335), .QN(n34307) );
  DFFRX1 dict_reg_239__5_ ( .D(n36440), .CK(clk), .RN(n42335), .QN(n34315) );
  DFFRX1 dict_reg_242__5_ ( .D(n36464), .CK(clk), .RN(n42336), .Q(n37202),
        .QN(n34339) );
  DFFRX1 dict_reg_243__5_ ( .D(n36472), .CK(clk), .RN(n42336), .QN(n34347) );
  DFFRX1 dict_reg_244__5_ ( .D(n36480), .CK(clk), .RN(n42336), .QN(n34355) );
  DFFRX1 dict_reg_245__5_ ( .D(n36488), .CK(clk), .RN(n42336), .QN(n34363) );
  DFFRX1 dict_reg_246__5_ ( .D(n36496), .CK(clk), .RN(n42336), .QN(n34371) );
  DFFRX1 dict_reg_247__5_ ( .D(n36504), .CK(clk), .RN(n42336), .QN(n34379) );
  DFFRX1 dict_reg_248__5_ ( .D(n36512), .CK(clk), .RN(n42336), .QN(n34387) );
  DFFRX1 dict_reg_251__5_ ( .D(n36536), .CK(clk), .RN(n42336), .Q(n37201),
        .QN(n34411) );
  DFFRX1 dict_reg_144__1_ ( .D(n35684), .CK(clk), .RN(n42365), .QN(n33559) );
  DFFRX1 dict_reg_145__1_ ( .D(n35692), .CK(clk), .RN(n42365), .Q(n37203),
        .QN(n33567) );
  DFFRX1 dict_reg_188__1_ ( .D(n36036), .CK(clk), .RN(n42369), .QN(n33911) );
  DFFRX1 dict_reg_189__1_ ( .D(n36044), .CK(clk), .RN(n42369), .QN(n33919) );
  DFFRX1 dict_reg_192__1_ ( .D(n36068), .CK(clk), .RN(n42369), .QN(n33943) );
  DFFRX1 dict_reg_203__1_ ( .D(n36156), .CK(clk), .RN(n42370), .QN(n34031) );
  DFFRX1 dict_reg_205__1_ ( .D(n36172), .CK(clk), .RN(n42370), .QN(n34047) );
  DFFRX1 dict_reg_206__1_ ( .D(n36180), .CK(clk), .RN(n42371), .QN(n34055) );
  DFFRX1 dict_reg_213__1_ ( .D(n36236), .CK(clk), .RN(n42371), .QN(n34111) );
  DFFRX1 dict_reg_214__1_ ( .D(n36244), .CK(clk), .RN(n42371), .QN(n34119) );
  DFFRX1 dict_reg_215__1_ ( .D(n36252), .CK(clk), .RN(n42371), .QN(n34127) );
  DFFRX1 dict_reg_216__1_ ( .D(n36260), .CK(clk), .RN(n42371), .QN(n34135) );
  DFFRX1 dict_reg_217__1_ ( .D(n36268), .CK(clk), .RN(n42371), .QN(n34143) );
  DFFRX1 dict_reg_218__1_ ( .D(n36276), .CK(clk), .RN(n42372), .QN(n34151) );
  DFFRX1 dict_reg_219__1_ ( .D(n36284), .CK(clk), .RN(n42372), .QN(n34159) );
  DFFRX1 dict_reg_220__1_ ( .D(n36292), .CK(clk), .RN(n42372), .QN(n34167) );
  DFFRX1 dict_reg_222__1_ ( .D(n36308), .CK(clk), .RN(n42372), .QN(n34183) );
  DFFRX1 dict_reg_223__1_ ( .D(n36316), .CK(clk), .RN(n42372), .QN(n34191) );
  DFFRX1 dict_reg_225__1_ ( .D(n36332), .CK(clk), .RN(n42372), .QN(n34207) );
  DFFRX1 dict_reg_226__1_ ( .D(n36340), .CK(clk), .RN(n42372), .QN(n34215) );
  DFFRX1 dict_reg_228__1_ ( .D(n36356), .CK(clk), .RN(n42372), .QN(n34231) );
  DFFRX1 dict_reg_229__1_ ( .D(n36364), .CK(clk), .RN(n42372), .QN(n34239) );
  DFFRX1 dict_reg_230__1_ ( .D(n36372), .CK(clk), .RN(n42373), .QN(n34247) );
  DFFRX1 dict_reg_232__1_ ( .D(n36388), .CK(clk), .RN(n42373), .QN(n34263) );
  DFFRX1 dict_reg_233__1_ ( .D(n36396), .CK(clk), .RN(n42373), .QN(n34271) );
  DFFRX1 dict_reg_235__1_ ( .D(n36412), .CK(clk), .RN(n42373), .QN(n34287) );
  DFFRX1 dict_reg_236__1_ ( .D(n36420), .CK(clk), .RN(n42373), .QN(n34295) );
  DFFRX1 dict_reg_237__1_ ( .D(n36428), .CK(clk), .RN(n42373), .QN(n34303) );
  DFFRX1 dict_reg_239__1_ ( .D(n36444), .CK(clk), .RN(n42373), .QN(n34319) );
  DFFRX1 dict_reg_242__1_ ( .D(n36468), .CK(clk), .RN(n42374), .QN(n34343) );
  DFFRX1 dict_reg_244__1_ ( .D(n36484), .CK(clk), .RN(n42374), .QN(n34359) );
  DFFRX1 dict_reg_246__1_ ( .D(n36500), .CK(clk), .RN(n42374), .QN(n34375) );
  DFFRX1 dict_reg_247__1_ ( .D(n36508), .CK(clk), .RN(n42374), .QN(n34383) );
  DFFRX1 dict_reg_193__5_ ( .D(n36072), .CK(clk), .RN(n42331), .Q(n37246),
        .QN(n33947) );
  DFFRX1 dict_reg_201__5_ ( .D(n36136), .CK(clk), .RN(n42332), .QN(n34011) );
  DFFRX1 dict_reg_250__5_ ( .D(n36528), .CK(clk), .RN(n42336), .QN(n34403) );
  DFFRX1 dict_reg_201__1_ ( .D(n36140), .CK(clk), .RN(n42370), .QN(n34015) );
  DFFRX1 dict_reg_240__1_ ( .D(n36452), .CK(clk), .RN(n42373), .QN(n34327) );
  DFFRX1 dict_reg_142__5_ ( .D(n35664), .CK(clk), .RN(n42327), .QN(n33539) );
  DFFRX1 dict_reg_151__5_ ( .D(n35736), .CK(clk), .RN(n42328), .QN(n33611) );
  DFFRX1 dict_reg_167__5_ ( .D(n35864), .CK(clk), .RN(n42329), .QN(n33739) );
  DFFRX1 dict_reg_168__5_ ( .D(n35872), .CK(clk), .RN(n42329), .QN(n33747) );
  DFFRX1 dict_reg_169__5_ ( .D(n35880), .CK(clk), .RN(n42329), .QN(n33755) );
  DFFRX1 dict_reg_170__5_ ( .D(n35888), .CK(clk), .RN(n42330), .QN(n33763) );
  DFFRX1 dict_reg_171__5_ ( .D(n35896), .CK(clk), .RN(n42330), .QN(n33771) );
  DFFRX1 dict_reg_185__5_ ( .D(n36008), .CK(clk), .RN(n42331), .Q(n37250),
        .QN(n33883) );
  DFFRX1 dict_reg_186__5_ ( .D(n36016), .CK(clk), .RN(n42331), .QN(n33891) );
  DFFRX1 dict_reg_187__5_ ( .D(n36024), .CK(clk), .RN(n42331), .QN(n33899) );
  DFFRX1 dict_reg_240__5_ ( .D(n36448), .CK(clk), .RN(n42335), .QN(n34323) );
  DFFRX1 dict_reg_241__5_ ( .D(n36456), .CK(clk), .RN(n42335), .QN(n34331) );
  DFFRX1 dict_reg_249__5_ ( .D(n36520), .CK(clk), .RN(n42336), .QN(n34395) );
  DFFRX1 dict_reg_142__1_ ( .D(n35668), .CK(clk), .RN(n42365), .QN(n33543) );
  DFFRX1 dict_reg_143__1_ ( .D(n35676), .CK(clk), .RN(n42365), .QN(n33551) );
  DFFRX1 dict_reg_150__1_ ( .D(n35732), .CK(clk), .RN(n42366), .QN(n33607) );
  DFFRX1 dict_reg_151__1_ ( .D(n35740), .CK(clk), .RN(n42366), .QN(n33615) );
  DFFRX1 dict_reg_167__1_ ( .D(n35868), .CK(clk), .RN(n42367), .QN(n33743) );
  DFFRX1 dict_reg_168__1_ ( .D(n35876), .CK(clk), .RN(n42367), .QN(n33751) );
  DFFRX1 dict_reg_169__1_ ( .D(n35884), .CK(clk), .RN(n42367), .QN(n33759) );
  DFFRX1 dict_reg_170__1_ ( .D(n35892), .CK(clk), .RN(n42368), .QN(n33767) );
  DFFRX1 dict_reg_171__1_ ( .D(n35900), .CK(clk), .RN(n42368), .QN(n33775) );
  DFFRX1 dict_reg_185__1_ ( .D(n36012), .CK(clk), .RN(n42369), .QN(n33887) );
  DFFRX1 dict_reg_186__1_ ( .D(n36020), .CK(clk), .RN(n42369), .QN(n33895) );
  DFFRX1 dict_reg_187__1_ ( .D(n36028), .CK(clk), .RN(n42369), .QN(n33903) );
  DFFRX1 dict_reg_250__1_ ( .D(n36532), .CK(clk), .RN(n42374), .QN(n34407) );
  DFFSRX1 enc_num_reg_0_ ( .D(n32394), .CK(clk), .SN(n37591), .RN(1'b1), .Q(
        n36933), .QN(n37521) );
  DFFSRXL drop_reg ( .D(drop_done), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n9651) );
  DFFSRXL data_queue_reg_2__3_ ( .D(n36616), .CK(clk), .SN(1'b1), .RN(n37593),
        .Q(n36927), .QN(n34455) );
  DFFSRXL data_num_reg_0_ ( .D(nxt_data_num[0]), .CK(clk), .SN(1'b1), .RN(
        n37593), .QN(n32400) );
  DFFSRXL dict_reg_174__1_ ( .D(n35924), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n33799) );
  DFFSRXL dict_reg_173__1_ ( .D(n35916), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33791) );
  DFFSRXL dict_reg_79__5_ ( .D(n35160), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n33035) );
  DFFSRXL dict_reg_255__0_ ( .D(n34518), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n9662) );
  DFFSRXL dict_reg_4__5_ ( .D(n34560), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32435) );
  DFFSRXL dict_reg_4__1_ ( .D(n34564), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32439) );
  DFFSRXL dict_reg_5__5_ ( .D(n34568), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32443) );
  DFFSRXL dict_reg_29__1_ ( .D(n34764), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32639) );
  DFFSRXL dict_reg_30__5_ ( .D(n34768), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32643) );
  DFFSRXL dict_reg_30__1_ ( .D(n34772), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32647) );
  DFFSRXL dict_reg_255__7_ ( .D(n34525), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n9660) );
  DFFSRXL dict_reg_255__6_ ( .D(n34524), .CK(clk), .SN(1'b1), .RN(n37590),
        .QN(n9658) );
  DFFSRXL dict_reg_3__5_ ( .D(n34552), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32427) );
  DFFSRXL dict_reg_3__1_ ( .D(n34556), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32431) );
  DFFSRXL dict_reg_255__5_ ( .D(n34523), .CK(clk), .SN(1'b1), .RN(n37594),
        .QN(n9656) );
  DFFSRXL dict_reg_255__4_ ( .D(n34522), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n41358), .QN(n9670) );
  DFFSRXL dict_reg_255__3_ ( .D(n34521), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n9668) );
  DFFSRXL dict_reg_255__2_ ( .D(n34520), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n9666) );
  DFFSRXL dict_reg_174__5_ ( .D(n35920), .CK(clk), .SN(1'b1), .RN(n37595),
        .QN(n33795) );
  DFFSRXL dict_reg_108__5_ ( .D(n35392), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n33267) );
  DFFSRXL dict_reg_125__1_ ( .D(n35532), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n33407) );
  DFFSRXL dict_reg_105__1_ ( .D(n35372), .CK(clk), .SN(1'b1), .RN(n37590),
        .QN(n33247) );
  DFFSRXL dict_reg_99__1_ ( .D(n35324), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n33199) );
  DFFSRXL dict_reg_99__5_ ( .D(n35320), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n33195) );
  DFFSRXL dict_reg_100__5_ ( .D(n35328), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n33203) );
  DFFSRXL dict_reg_100__1_ ( .D(n35332), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33207) );
  DFFSRXL dict_reg_97__1_ ( .D(n35308), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n33183) );
  DFFSRXL dict_reg_97__5_ ( .D(n35304), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n33179) );
  DFFSRXL dict_reg_95__1_ ( .D(n35292), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n33167) );
  DFFSRXL dict_reg_98__5_ ( .D(n35312), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n33187) );
  DFFSRXL dict_reg_98__1_ ( .D(n35316), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n33191) );
  DFFSRXL dict_reg_95__5_ ( .D(n35288), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n33163) );
  DFFSRXL dict_reg_96__5_ ( .D(n35296), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n33171) );
  DFFSRXL dict_reg_96__1_ ( .D(n35300), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n33175) );
  DFFSRXL dict_reg_15__5_ ( .D(n34648), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32523) );
  DFFSRXL dict_reg_13__1_ ( .D(n34636), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32511) );
  DFFSRXL dict_reg_16__5_ ( .D(n34656), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32531) );
  DFFSRXL dict_reg_16__1_ ( .D(n34660), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32535) );
  DFFSRXL dict_reg_15__1_ ( .D(n34652), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32527) );
  DFFSRXL dict_reg_14__5_ ( .D(n34640), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32515) );
  DFFSRXL dict_reg_14__1_ ( .D(n34644), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32519) );
  DFFSRXL dict_reg_17__5_ ( .D(n34664), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32539) );
  DFFSRXL dict_reg_17__1_ ( .D(n34668), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32543) );
  DFFSRXL dict_reg_62__5_ ( .D(n35024), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32899) );
  DFFSRXL dict_reg_62__1_ ( .D(n35028), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32903) );
  DFFSRXL dict_reg_61__5_ ( .D(n35016), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32891) );
  DFFSRXL dict_reg_61__1_ ( .D(n35020), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32895) );
  DFFSRXL dict_reg_60__5_ ( .D(n35008), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32883) );
  DFFSRXL dict_reg_60__1_ ( .D(n35012), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32887) );
  DFFSRXL dict_reg_21__5_ ( .D(n34696), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32571) );
  DFFSRXL dict_reg_19__5_ ( .D(n34680), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n32555) );
  DFFSRXL dict_reg_19__1_ ( .D(n34684), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32559) );
  DFFSRXL dict_reg_18__5_ ( .D(n34672), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32547) );
  DFFSRXL dict_reg_18__1_ ( .D(n34676), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32551) );
  DFFSRXL dict_reg_35__5_ ( .D(n34808), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32683) );
  DFFSRXL dict_reg_35__1_ ( .D(n34812), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32687) );
  DFFSRXL dict_reg_34__5_ ( .D(n34800), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32675) );
  DFFSRXL dict_reg_34__1_ ( .D(n34804), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32679) );
  DFFSRXL dict_reg_33__5_ ( .D(n34792), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32667) );
  DFFSRXL dict_reg_33__1_ ( .D(n34796), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32671) );
  DFFSRXL dict_reg_31__5_ ( .D(n34776), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32651) );
  DFFSRXL dict_reg_31__1_ ( .D(n34780), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32655) );
  DFFSRXL dict_reg_51__5_ ( .D(n34936), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32811) );
  DFFSRXL dict_reg_51__1_ ( .D(n34940), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32815) );
  DFFSRXL dict_reg_50__5_ ( .D(n34928), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32803) );
  DFFSRXL dict_reg_50__1_ ( .D(n34932), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32807) );
  DFFSRXL dict_reg_49__5_ ( .D(n34920), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32795) );
  DFFSRXL dict_reg_49__1_ ( .D(n34924), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32799) );
  DFFSRXL dict_reg_48__5_ ( .D(n34912), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32787) );
  DFFSRXL dict_reg_48__1_ ( .D(n34916), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32791) );
  DFFSRXL dict_reg_20__5_ ( .D(n34688), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32563) );
  DFFSRXL dict_reg_20__1_ ( .D(n34692), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n32567) );
  DFFSRXL dict_reg_56__5_ ( .D(n34976), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32851) );
  DFFSRXL dict_reg_55__1_ ( .D(n34972), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n32847) );
  DFFSRXL dict_reg_37__5_ ( .D(n34824), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32699) );
  DFFSRXL dict_reg_36__5_ ( .D(n34816), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32691) );
  DFFSRXL dict_reg_36__1_ ( .D(n34820), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32695) );
  DFFSRXL dict_reg_32__5_ ( .D(n34784), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32659) );
  DFFSRXL dict_reg_32__1_ ( .D(n34788), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32663) );
  DFFSRXL dict_reg_59__5_ ( .D(n35000), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32875) );
  DFFSRXL dict_reg_59__1_ ( .D(n35004), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32879) );
  DFFSRXL dict_reg_58__5_ ( .D(n34992), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32867) );
  DFFSRXL dict_reg_58__1_ ( .D(n34996), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32871) );
  DFFSRXL dict_reg_57__5_ ( .D(n34984), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32859) );
  DFFSRXL dict_reg_57__1_ ( .D(n34988), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32863) );
  DFFSRXL dict_reg_56__1_ ( .D(n34980), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32855) );
  DFFSRXL dict_reg_55__5_ ( .D(n34968), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32843) );
  DFFSRXL dict_reg_54__5_ ( .D(n34960), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32835) );
  DFFSRXL dict_reg_54__1_ ( .D(n34964), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32839) );
  DFFSRXL dict_reg_53__5_ ( .D(n34952), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32827) );
  DFFSRXL dict_reg_53__1_ ( .D(n34956), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32831) );
  DFFSRXL dict_reg_52__5_ ( .D(n34944), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32819) );
  DFFSRXL dict_reg_52__1_ ( .D(n34948), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32823) );
  DFFSRXL dict_reg_47__5_ ( .D(n34904), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32779) );
  DFFSRXL dict_reg_47__1_ ( .D(n34908), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32783) );
  DFFSRXL dict_reg_255__1_ ( .D(n34519), .CK(clk), .SN(1'b1), .RN(n37590),
        .QN(n9664) );
  DFFSRXL dict_reg_117__5_ ( .D(n35464), .CK(clk), .SN(1'b1), .RN(n37595),
        .QN(n33339) );
  DFFSRXL dict_reg_117__1_ ( .D(n35468), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33343) );
  DFFSRXL dict_reg_114__1_ ( .D(n35444), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n33319) );
  DFFSRXL dict_reg_71__5_ ( .D(n35096), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32971) );
  DFFSRXL dict_reg_71__1_ ( .D(n35100), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32975) );
  DFFSRXL dict_reg_93__5_ ( .D(n35272), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n33147) );
  DFFSRXL dict_reg_91__5_ ( .D(n35256), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n33131) );
  DFFSRXL dict_reg_91__1_ ( .D(n35260), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n33135) );
  DFFSRXL dict_reg_90__1_ ( .D(n35252), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n33127) );
  DFFSRXL dict_reg_87__5_ ( .D(n35224), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n33099) );
  DFFSRXL dict_reg_82__5_ ( .D(n35184), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n33059) );
  DFFSRXL dict_reg_78__5_ ( .D(n35152), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n33027) );
  DFFSRXL dict_reg_78__1_ ( .D(n35156), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n33031) );
  DFFSRXL dict_reg_77__1_ ( .D(n35148), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n33023) );
  DFFSRXL dict_reg_92__5_ ( .D(n35264), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n33139) );
  DFFSRXL dict_reg_92__1_ ( .D(n35268), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n33143) );
  DFFSRXL dict_reg_90__5_ ( .D(n35248), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n33123) );
  DFFSRXL dict_reg_89__5_ ( .D(n35240), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n33115) );
  DFFSRXL dict_reg_89__1_ ( .D(n35244), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n33119) );
  DFFSRXL dict_reg_88__5_ ( .D(n35232), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n33107) );
  DFFSRXL dict_reg_88__1_ ( .D(n35236), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n33111) );
  DFFSRXL dict_reg_87__1_ ( .D(n35228), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n33103) );
  DFFSRXL dict_reg_86__5_ ( .D(n35216), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n33091) );
  DFFSRXL dict_reg_86__1_ ( .D(n35220), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n33095) );
  DFFSRXL dict_reg_85__5_ ( .D(n35208), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n33083) );
  DFFSRXL dict_reg_85__1_ ( .D(n35212), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n33087) );
  DFFSRXL dict_reg_84__5_ ( .D(n35200), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n33075) );
  DFFSRXL dict_reg_83__5_ ( .D(n35192), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n33067) );
  DFFSRXL dict_reg_83__1_ ( .D(n35196), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n33071) );
  DFFSRXL dict_reg_82__1_ ( .D(n35188), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n33063) );
  DFFSRXL dict_reg_81__5_ ( .D(n35176), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n33051) );
  DFFSRXL dict_reg_81__1_ ( .D(n35180), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n33055) );
  DFFSRXL dict_reg_80__5_ ( .D(n35168), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n33043) );
  DFFSRXL dict_reg_80__1_ ( .D(n35172), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n33047) );
  DFFSRXL dict_reg_94__5_ ( .D(n35280), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n33155) );
  DFFSRXL dict_reg_93__1_ ( .D(n35276), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n33151) );
  DFFSRXL dict_reg_84__1_ ( .D(n35204), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n33079) );
  DFFSRXL dict_reg_79__1_ ( .D(n35164), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n33039) );
  DFFSRXL dict_reg_94__1_ ( .D(n35284), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n33159) );
  DFFSRXL dict_reg_77__5_ ( .D(n35144), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n33019) );
  DFFSRXL dict_reg_76__5_ ( .D(n35136), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n33011) );
  DFFSRXL dict_reg_76__1_ ( .D(n35140), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n33015) );
  DFFSRXL dict_reg_75__1_ ( .D(n35132), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n33007) );
  DFFSRXL dict_reg_75__5_ ( .D(n35128), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n33003) );
  DFFSRXL dict_reg_63__5_ ( .D(n35032), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32907) );
  DFFSRXL dict_reg_74__5_ ( .D(n35120), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32995) );
  DFFSRXL dict_reg_74__1_ ( .D(n35124), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32999) );
  DFFSRXL dict_reg_73__1_ ( .D(n35116), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32991) );
  DFFSRXL dict_reg_73__5_ ( .D(n35112), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32987) );
  DFFSRXL dict_reg_70__5_ ( .D(n35088), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n32963) );
  DFFSRXL dict_reg_70__1_ ( .D(n35092), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32967) );
  DFFSRXL dict_reg_69__1_ ( .D(n35084), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32959) );
  DFFSRXL dict_reg_72__5_ ( .D(n35104), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32979) );
  DFFSRXL dict_reg_72__1_ ( .D(n35108), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32983) );
  DFFSRXL dict_reg_69__5_ ( .D(n35080), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32955) );
  DFFSRXL dict_reg_68__5_ ( .D(n35072), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32947) );
  DFFSRXL dict_reg_68__1_ ( .D(n35076), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32951) );
  DFFSRXL dict_reg_64__5_ ( .D(n35040), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32915) );
  DFFSRXL dict_reg_64__1_ ( .D(n35044), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32919) );
  DFFSRXL dict_reg_63__1_ ( .D(n35036), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32911) );
  DFFSRXL dict_reg_67__5_ ( .D(n35064), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32939) );
  DFFSRXL dict_reg_67__1_ ( .D(n35068), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32943) );
  DFFSRXL dict_reg_66__5_ ( .D(n35056), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32931) );
  DFFSRXL dict_reg_66__1_ ( .D(n35060), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32935) );
  DFFSRXL dict_reg_65__5_ ( .D(n35048), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32923) );
  DFFSRXL dict_reg_65__1_ ( .D(n35052), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32927) );
  DFFSRXL dict_reg_150__5_ ( .D(n35728), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n33603) );
  DFFSRXL dict_reg_179__1_ ( .D(n35964), .CK(clk), .SN(1'b1), .RN(n37594),
        .QN(n33839) );
  DFFSRXL dict_reg_178__1_ ( .D(n35956), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33831) );
  DFFSRXL dict_reg_177__1_ ( .D(n35948), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33823) );
  DFFSRXL dict_reg_176__1_ ( .D(n35940), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n33815) );
  DFFSRXL dict_reg_148__1_ ( .D(n35716), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n33591) );
  DFFSRXL dict_reg_177__5_ ( .D(n35944), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n33819) );
  DFFSRXL dict_reg_149__1_ ( .D(n35724), .CK(clk), .SN(1'b1), .RN(n37590),
        .QN(n33599) );
  DFFSRXL dict_reg_184__1_ ( .D(n36004), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n33879) );
  DFFSRXL dict_reg_154__1_ ( .D(n35764), .CK(clk), .SN(1'b1), .RN(n37595),
        .QN(n33639) );
  DFFSRXL dict_reg_190__1_ ( .D(n36052), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n33927) );
  DFFSRXL dict_reg_182__1_ ( .D(n35988), .CK(clk), .SN(1'b1), .RN(n37599),
        .QN(n33863) );
  DFFSRXL dict_reg_181__1_ ( .D(n35980), .CK(clk), .SN(1'b1), .RN(n37599),
        .QN(n33855) );
  DFFSRXL dict_reg_180__1_ ( .D(n35972), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n37249), .QN(n33847) );
  DFFSRXL dict_reg_175__1_ ( .D(n35932), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n33807) );
  DFFSRXL dict_reg_147__1_ ( .D(n35708), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n33583) );
  DFFSRXL dict_reg_138__5_ ( .D(n35632), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33507) );
  DFFSRXL dict_reg_138__1_ ( .D(n35636), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n33511) );
  DFFSRXL dict_reg_137__1_ ( .D(n35628), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33503) );
  DFFSRXL dict_reg_136__1_ ( .D(n35620), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n33495) );
  DFFSRXL dict_reg_155__1_ ( .D(n35772), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33647) );
  DFFSRXL dict_reg_146__1_ ( .D(n35700), .CK(clk), .SN(1'b1), .RN(n37595),
        .QN(n33575) );
  DFFSRXL dict_reg_2__5_ ( .D(n34544), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32419) );
  DFFSRXL dict_reg_2__1_ ( .D(n34548), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32423) );
  DFFSRXL dict_reg_109__5_ ( .D(n35400), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33275) );
  DFFSRXL dict_reg_108__1_ ( .D(n35396), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n33271) );
  DFFSRXL dict_reg_107__1_ ( .D(n35388), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n33263) );
  DFFSRXL dict_reg_126__5_ ( .D(n35536), .CK(clk), .SN(1'b1), .RN(n37594),
        .QN(n33411) );
  DFFSRXL dict_reg_125__5_ ( .D(n35528), .CK(clk), .SN(1'b1), .RN(n37599),
        .QN(n33403) );
  DFFSRXL dict_reg_107__5_ ( .D(n35384), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n33259) );
  DFFSRXL dict_reg_106__5_ ( .D(n35376), .CK(clk), .SN(1'b1), .RN(n37599),
        .QN(n33251) );
  DFFSRXL dict_reg_106__1_ ( .D(n35380), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n33255) );
  DFFSRXL dict_reg_105__5_ ( .D(n35368), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n33243) );
  DFFSRXL dict_reg_104__5_ ( .D(n35360), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n33235) );
  DFFSRXL dict_reg_104__1_ ( .D(n35364), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n33239) );
  DFFSRXL dict_reg_103__5_ ( .D(n35352), .CK(clk), .SN(1'b1), .RN(n37595),
        .QN(n33227) );
  DFFSRXL dict_reg_103__1_ ( .D(n35356), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n33231) );
  DFFSRXL dict_reg_102__5_ ( .D(n35344), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33219) );
  DFFSRXL dict_reg_102__1_ ( .D(n35348), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33223) );
  DFFSRXL dict_reg_101__5_ ( .D(n35336), .CK(clk), .SN(1'b1), .RN(n37594),
        .QN(n33211) );
  DFFSRXL dict_reg_101__1_ ( .D(n35340), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n33215) );
  DFFSRXL dict_reg_109__1_ ( .D(n35404), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n33279) );
  DFFSRXL dict_reg_110__5_ ( .D(n35408), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n33283) );
  DFFSRXL dict_reg_110__1_ ( .D(n35412), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n33287) );
  DFFSRXL dict_reg_1__5_ ( .D(n34536), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32411) );
  DFFSRXL dict_reg_1__1_ ( .D(n34540), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32415) );
  DFFSRXL dict_reg_0__5_ ( .D(n34528), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32403) );
  DFFSRXL dict_reg_0__1_ ( .D(n34532), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32407) );
  DFFSRXL dict_reg_13__5_ ( .D(n34632), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32507) );
  DFFSRXL dict_reg_11__5_ ( .D(n34616), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32491) );
  DFFSRXL dict_reg_11__1_ ( .D(n34620), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32495) );
  DFFSRXL dict_reg_10__5_ ( .D(n34608), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32483) );
  DFFSRXL dict_reg_10__1_ ( .D(n34612), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32487) );
  DFFSRXL dict_reg_9__5_ ( .D(n34600), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32475) );
  DFFSRXL dict_reg_9__1_ ( .D(n34604), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32479) );
  DFFSRXL dict_reg_8__5_ ( .D(n34592), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32467) );
  DFFSRXL dict_reg_8__1_ ( .D(n34596), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32471) );
  DFFSRXL dict_reg_7__5_ ( .D(n34584), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32459) );
  DFFSRXL dict_reg_7__1_ ( .D(n34588), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32463) );
  DFFSRXL dict_reg_6__5_ ( .D(n34576), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32451) );
  DFFSRXL dict_reg_6__1_ ( .D(n34580), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32455) );
  DFFSRXL dict_reg_5__1_ ( .D(n34572), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n32447) );
  DFFSRXL dict_reg_25__5_ ( .D(n34728), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32603) );
  DFFSRXL dict_reg_25__1_ ( .D(n34732), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n32607) );
  DFFSRXL dict_reg_23__5_ ( .D(n34712), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32587) );
  DFFSRXL dict_reg_23__1_ ( .D(n34716), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32591) );
  DFFSRXL dict_reg_12__5_ ( .D(n34624), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32499) );
  DFFSRXL dict_reg_12__1_ ( .D(n34628), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32503) );
  DFFSRXL dict_reg_29__5_ ( .D(n34760), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32635) );
  DFFSRXL dict_reg_28__1_ ( .D(n34756), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32631) );
  DFFSRXL dict_reg_28__5_ ( .D(n34752), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32627) );
  DFFSRXL dict_reg_27__5_ ( .D(n34744), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32619) );
  DFFSRXL dict_reg_27__1_ ( .D(n34748), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32623) );
  DFFSRXL dict_reg_26__5_ ( .D(n34736), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32611) );
  DFFSRXL dict_reg_26__1_ ( .D(n34740), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32615) );
  DFFSRXL dict_reg_24__5_ ( .D(n34720), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32595) );
  DFFSRXL dict_reg_24__1_ ( .D(n34724), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32599) );
  DFFSRXL dict_reg_22__5_ ( .D(n34704), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32579) );
  DFFSRXL dict_reg_22__1_ ( .D(n34708), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32583) );
  DFFSRXL dict_reg_21__1_ ( .D(n34700), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32575) );
  DFFSRXL dict_reg_251__1_ ( .D(n36540), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n34415) );
  DFFSRXL dict_reg_248__1_ ( .D(n36516), .CK(clk), .SN(1'b1), .RN(n37595),
        .QN(n34391) );
  DFFSRXL dict_reg_231__1_ ( .D(n36380), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n34255) );
  DFFSRXL dict_reg_227__1_ ( .D(n36348), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n34223) );
  DFFSRXL dict_reg_194__1_ ( .D(n36084), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n33959) );
  DFFSRXL dict_reg_241__1_ ( .D(n36460), .CK(clk), .SN(1'b1), .RN(n37594),
        .QN(n34335) );
  DFFSRXL dict_reg_238__1_ ( .D(n36436), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n34311) );
  DFFSRXL dict_reg_234__1_ ( .D(n36404), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n34279) );
  DFFSRXL dict_reg_224__1_ ( .D(n36324), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n34199) );
  DFFSRXL dict_reg_210__1_ ( .D(n36212), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n34087) );
  DFFSRXL dict_reg_193__1_ ( .D(n36076), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n37248), .QN(n33951) );
  DFFSRXL dict_reg_245__1_ ( .D(n36492), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n34367) );
  DFFSRXL dict_reg_211__5_ ( .D(n36216), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n34091) );
  DFFSRXL dict_reg_204__5_ ( .D(n36160), .CK(clk), .SN(1'b1), .RN(n37595),
        .QN(n34035) );
  DFFSRXL dict_reg_204__1_ ( .D(n36164), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n34039) );
  DFFSRXL dict_reg_211__1_ ( .D(n36220), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n34095) );
  DFFSRXL dict_reg_199__1_ ( .D(n36124), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n33999) );
  DFFSRXL dict_reg_196__1_ ( .D(n36100), .CK(clk), .SN(1'b1), .RN(n37594),
        .QN(n33975) );
  DFFSRXL dict_reg_195__1_ ( .D(n36092), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n33967) );
  DFFSRXL dict_reg_221__1_ ( .D(n36300), .CK(clk), .SN(1'b1), .RN(n37599),
        .QN(n34175) );
  DFFSRXL dict_reg_212__5_ ( .D(n36224), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n34099) );
  DFFSRXL dict_reg_202__1_ ( .D(n36148), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n34023) );
  DFFSRXL dict_reg_197__1_ ( .D(n36108), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n33983) );
  DFFSRXL dict_reg_40__1_ ( .D(n34852), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32727) );
  DFFSRXL dict_reg_42__5_ ( .D(n34864), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32739) );
  DFFSRXL dict_reg_41__5_ ( .D(n34856), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32731) );
  DFFSRXL dict_reg_41__1_ ( .D(n34860), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32735) );
  DFFSRXL dict_reg_46__5_ ( .D(n34896), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32771) );
  DFFSRXL dict_reg_46__1_ ( .D(n34900), .CK(clk), .SN(1'b1), .RN(n37599), .QN(
        n32775) );
  DFFSRXL dict_reg_44__5_ ( .D(n34880), .CK(clk), .SN(1'b1), .RN(n37601), .QN(
        n32755) );
  DFFSRXL dict_reg_44__1_ ( .D(n34884), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n32759) );
  DFFSRXL dict_reg_43__5_ ( .D(n34872), .CK(clk), .SN(1'b1), .RN(n37596), .QN(
        n32747) );
  DFFSRXL dict_reg_43__1_ ( .D(n34876), .CK(clk), .SN(1'b1), .RN(n37591), .QN(
        n32751) );
  DFFSRXL dict_reg_40__5_ ( .D(n34848), .CK(clk), .SN(1'b1), .RN(n37590), .QN(
        n32723) );
  DFFSRXL dict_reg_45__1_ ( .D(n34892), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32767) );
  DFFSRXL dict_reg_42__1_ ( .D(n34868), .CK(clk), .SN(1'b1), .RN(n37595), .QN(
        n32743) );
  DFFSRXL dict_reg_39__5_ ( .D(n34840), .CK(clk), .SN(1'b1), .RN(n37598), .QN(
        n32715) );
  DFFSRXL dict_reg_38__5_ ( .D(n34832), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32707) );
  DFFSRXL dict_reg_38__1_ ( .D(n34836), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n32711) );
  DFFSRXL dict_reg_37__1_ ( .D(n34828), .CK(clk), .SN(1'b1), .RN(n37594), .QN(
        n32703) );
  DFFSRXL dict_reg_45__5_ ( .D(n34888), .CK(clk), .SN(1'b1), .RN(n37593), .QN(
        n32763) );
  DFFSRXL dict_reg_39__1_ ( .D(n34844), .CK(clk), .SN(1'b1), .RN(n37592), .QN(
        n32719) );
  DFFSRXL dict_reg_126__1_ ( .D(n35540), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n33415) );
  DFFSRXL dict_reg_118__5_ ( .D(n35472), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n33347) );
  DFFSRXL dict_reg_118__1_ ( .D(n35476), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n33351) );
  DFFSRXL dict_reg_116__5_ ( .D(n35456), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n33331) );
  DFFSRXL dict_reg_116__1_ ( .D(n35460), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n33335) );
  DFFSRXL dict_reg_115__1_ ( .D(n35452), .CK(clk), .SN(1'b1), .RN(n37590),
        .QN(n33327) );
  DFFSRXL data_queue_reg_4__7_ ( .D(n36604), .CK(clk), .SN(1'b1), .RN(n37599),
        .Q(n36762), .QN(n34467) );
  DFFSRXL data_queue_reg_4__5_ ( .D(n36602), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n34469) );
  DFFSRXL data_queue_reg_4__4_ ( .D(n36601), .CK(clk), .SN(1'b1), .RN(n37600),
        .Q(n36738), .QN(n34470) );
  DFFSRXL data_queue_reg_4__3_ ( .D(n36600), .CK(clk), .SN(1'b1), .RN(n37592),
        .Q(n36712), .QN(n34471) );
  DFFSRXL data_queue_reg_4__2_ ( .D(n36599), .CK(clk), .SN(1'b1), .RN(n37594),
        .Q(n36787), .QN(n34472) );
  DFFSRXL data_queue_reg_4__1_ ( .D(n36598), .CK(clk), .SN(1'b1), .RN(n37598),
        .Q(n36751), .QN(n34473) );
  DFFSRXL data_queue_reg_4__0_ ( .D(n36597), .CK(clk), .SN(1'b1), .RN(n37599),
        .QN(n34474) );
  DFFSRXL data_queue_reg_1__1_ ( .D(n36622), .CK(clk), .SN(1'b1), .RN(n37601),
        .Q(n36919), .QN(n34449) );
  DFFSRXL data_queue_reg_3__6_ ( .D(n36611), .CK(clk), .SN(1'b1), .RN(n37598),
        .Q(n36835), .QN(n34460) );
  DFFSRXL data_queue_reg_3__0_ ( .D(n36605), .CK(clk), .SN(1'b1), .RN(n37592),
        .Q(n36848), .QN(n34466) );
  DFFSRXL dict_reg_251__0_ ( .D(n36541), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n37551), .QN(n34416) );
  DFFSRX1 enc_num_reg_5_ ( .D(n32389), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n37189), .QN(n37534) );
  DFFSRX1 enc_num_reg_4_ ( .D(n32390), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n37190), .QN(n37535) );
  DFFSRX1 enc_num_reg_3_ ( .D(n32391), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n37184), .QN(n37522) );
  DFFSRX1 enc_num_reg_2_ ( .D(n32392), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n37185), .QN(n37523) );
  DFFSRX1 enc_num_reg_1_ ( .D(n32393), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n37186), .QN(n37524) );
  DFFSRX1 enc_num_reg_6_ ( .D(n32388), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n37188), .QN(n37533) );
  DFFSRX1 enc_num_reg_7_ ( .D(n32387), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n37187), .QN(n37532) );
  DFFSRX1 enc_num_reg_8_ ( .D(n32386), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n37193), .QN(n37531) );
  DFFSRX1 enc_num_reg_9_ ( .D(n32385), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n37192), .QN(n37539) );
  DFFSRX1 enc_num_reg_10_ ( .D(n32384), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n37191), .QN(n37537) );
  DFFSRX1 enc_num_reg_11_ ( .D(n32395), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n37194), .QN(n37538) );
  DFFSRX1 codeword_reg_10_ ( .D(n34507), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51439), .QN(n9652) );
  DFFSRX1 codeword_reg_1_ ( .D(n34516), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51446), .QN(n9653) );
  DFFSRX1 codeword_reg_0_ ( .D(n34517), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51447), .QN(n9654) );
  DFFSRX1 codeword_reg_6_ ( .D(n34511), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51443), .QN(n9671) );
  DFFSRX1 codeword_reg_5_ ( .D(n34512), .CK(clk), .SN(1'b1), .RN(n37600), .QN(
        n37536) );
  DFFSRX1 codeword_reg_9_ ( .D(n34508), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51440), .QN(n9676) );
  DFFSRX1 codeword_reg_7_ ( .D(n34510), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51442), .QN(n9678) );
  DFFSRX1 codeword_reg_8_ ( .D(n34509), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51441), .QN(n9677) );
  DFFSRXL codeword_reg_4_ ( .D(n34513), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51444), .QN(n40038) );
  DFFSRXL codeword_reg_2_ ( .D(n34515), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51445), .QN(n40772) );
  DFFSRX2 dict_reg_245__4_ ( .D(n36489), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n41270), .QN(n34364) );
  DFFSRX2 dict_reg_225__0_ ( .D(n36333), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n41231), .QN(n34208) );
  DFFSRX2 dict_reg_249__2_ ( .D(n36523), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n41367), .QN(n34398) );
  DFFSRX2 dict_reg_250__0_ ( .D(n36533), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n41234), .QN(n34408) );
  DFFSRX2 dict_reg_248__6_ ( .D(n36511), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49355), .QN(n34386) );
  DFFSRX2 dict_reg_245__0_ ( .D(n36493), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n41349), .QN(n34368) );
  DFFSRX2 dict_reg_222__0_ ( .D(n36309), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n41259), .QN(n34184) );
  DFFSRX2 dict_reg_246__2_ ( .D(n36499), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n41655), .QN(n34374) );
  DFFSRX2 dict_reg_225__7_ ( .D(n36326), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n41227), .QN(n34201) );
  DFFSRX2 dict_reg_249__4_ ( .D(n36521), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n41387), .QN(n34396) );
  DFFSRX2 dict_reg_240__0_ ( .D(n36453), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49074), .QN(n34328) );
  DFFSRX2 dict_reg_230__6_ ( .D(n36367), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n41221), .QN(n34242) );
  DFFSRX2 dict_reg_240__4_ ( .D(n36449), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48606), .QN(n34324) );
  DFFSRX2 dict_reg_243__2_ ( .D(n36475), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48910), .QN(n34350) );
  DFFSRX2 dict_reg_244__2_ ( .D(n36483), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n48906), .QN(n34358) );
  DFFSRX2 dict_reg_249__3_ ( .D(n36522), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n48730), .QN(n34397) );
  DFFSRX2 dict_reg_249__6_ ( .D(n36519), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49351), .QN(n34394) );
  DFFSRX2 dict_reg_230__0_ ( .D(n36373), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49114), .QN(n34248) );
  DFFSRX2 dict_reg_249__7_ ( .D(n36518), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49196), .QN(n34393) );
  DFFSRX2 dict_reg_29__3_ ( .D(n34762), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51040), .QN(n32637) );
  DFFSRX2 dict_reg_29__2_ ( .D(n34763), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50826), .QN(n32638) );
  DFFSRX2 dict_reg_29__0_ ( .D(n34765), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50612), .QN(n32640) );
  DFFSRX2 dict_reg_55__3_ ( .D(n34970), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51066), .QN(n32845) );
  DFFSRX2 dict_reg_55__2_ ( .D(n34971), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50852), .QN(n32846) );
  DFFSRX2 dict_reg_55__0_ ( .D(n34973), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50638), .QN(n32848) );
  DFFSRX2 dict_reg_32__2_ ( .D(n34787), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50829), .QN(n32662) );
  DFFSRX2 dict_reg_32__0_ ( .D(n34789), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50615), .QN(n32664) );
  DFFSRX2 dict_reg_54__2_ ( .D(n34963), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50851), .QN(n32838) );
  DFFSRX2 dict_reg_53__3_ ( .D(n34954), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51064), .QN(n32829) );
  DFFSRX2 dict_reg_53__2_ ( .D(n34955), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50850), .QN(n32830) );
  DFFSRX2 dict_reg_53__0_ ( .D(n34957), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50636), .QN(n32832) );
  DFFSRX2 dict_reg_52__3_ ( .D(n34946), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51063), .QN(n32821) );
  DFFSRX2 dict_reg_52__2_ ( .D(n34947), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50849), .QN(n32822) );
  DFFSRX2 dict_reg_52__0_ ( .D(n34949), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50635), .QN(n32824) );
  DFFSRX2 dict_reg_51__3_ ( .D(n34938), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51062), .QN(n32813) );
  DFFSRX2 dict_reg_51__2_ ( .D(n34939), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50848), .QN(n32814) );
  DFFSRX2 dict_reg_51__0_ ( .D(n34941), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50634), .QN(n32816) );
  DFFSRX2 dict_reg_50__3_ ( .D(n34930), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51061), .QN(n32805) );
  DFFSRX2 dict_reg_50__2_ ( .D(n34931), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50847), .QN(n32806) );
  DFFSRX2 dict_reg_50__0_ ( .D(n34933), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50633), .QN(n32808) );
  DFFSRX2 dict_reg_17__3_ ( .D(n34666), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51028), .QN(n32541) );
  DFFSRX2 dict_reg_16__3_ ( .D(n34658), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51027), .QN(n32533) );
  DFFSRX2 dict_reg_27__3_ ( .D(n34746), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51038), .QN(n32621) );
  DFFSRX2 dict_reg_27__2_ ( .D(n34747), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50824), .QN(n32622) );
  DFFSRX2 dict_reg_27__0_ ( .D(n34749), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50610), .QN(n32624) );
  DFFSRX2 dict_reg_26__3_ ( .D(n34738), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51037), .QN(n32613) );
  DFFSRX2 dict_reg_26__2_ ( .D(n34739), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50823), .QN(n32614) );
  DFFSRX2 dict_reg_26__0_ ( .D(n34741), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50609), .QN(n32616) );
  DFFSRX2 dict_reg_43__3_ ( .D(n34874), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51054), .QN(n32749) );
  DFFSRX2 dict_reg_43__2_ ( .D(n34875), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50840), .QN(n32750) );
  DFFSRX2 dict_reg_43__0_ ( .D(n34877), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50626), .QN(n32752) );
  DFFSRX2 dict_reg_252__5_ ( .D(n36544), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n34419) );
  DFFSRX2 dict_reg_224__0_ ( .D(n36325), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49137), .QN(n34200) );
  DFFSRX2 dict_reg_246__0_ ( .D(n36501), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49051), .QN(n34376) );
  DFFSRX2 dict_reg_30__3_ ( .D(n34770), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51041), .QN(n32645) );
  DFFSRX2 dict_reg_30__2_ ( .D(n34771), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50827), .QN(n32646) );
  DFFSRX2 dict_reg_30__0_ ( .D(n34773), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50613), .QN(n32648) );
  DFFSRX2 dict_reg_56__3_ ( .D(n34978), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51067), .QN(n32853) );
  DFFSRX2 dict_reg_33__2_ ( .D(n34795), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50830), .QN(n32670) );
  DFFSRX2 dict_reg_33__0_ ( .D(n34797), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50616), .QN(n32672) );
  DFFSRX2 dict_reg_32__3_ ( .D(n34786), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51043), .QN(n32661) );
  DFFSRX2 dict_reg_31__3_ ( .D(n34778), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51042), .QN(n32653) );
  DFFSRX2 dict_reg_31__0_ ( .D(n34781), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50614), .QN(n32656) );
  DFFSRX2 dict_reg_56__2_ ( .D(n34979), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50853), .QN(n32854) );
  DFFSRX2 dict_reg_54__3_ ( .D(n34962), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51065), .QN(n32837) );
  DFFSRX2 dict_reg_54__0_ ( .D(n34965), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50637), .QN(n32840) );
  DFFSRX2 dict_reg_49__3_ ( .D(n34922), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51060), .QN(n32797) );
  DFFSRX2 dict_reg_49__2_ ( .D(n34923), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50846), .QN(n32798) );
  DFFSRX2 dict_reg_49__0_ ( .D(n34925), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50632), .QN(n32800) );
  DFFSRX2 dict_reg_18__3_ ( .D(n34674), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51029), .QN(n32549) );
  DFFSRX2 dict_reg_18__2_ ( .D(n34675), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50815), .QN(n32550) );
  DFFSRX2 dict_reg_18__0_ ( .D(n34677), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50601), .QN(n32552) );
  DFFSRX2 dict_reg_17__2_ ( .D(n34667), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50814), .QN(n32542) );
  DFFSRX2 dict_reg_17__0_ ( .D(n34669), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50600), .QN(n32544) );
  DFFSRX2 dict_reg_16__2_ ( .D(n34659), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50813), .QN(n32534) );
  DFFSRX2 dict_reg_16__0_ ( .D(n34661), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50599), .QN(n32536) );
  DFFSRX2 dict_reg_28__0_ ( .D(n34757), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50611), .QN(n32632) );
  DFFSRX2 dict_reg_28__3_ ( .D(n34754), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51039), .QN(n32629) );
  DFFSRX2 dict_reg_28__2_ ( .D(n34755), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50825), .QN(n32630) );
  DFFSRX2 dict_reg_24__3_ ( .D(n34722), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51035), .QN(n32597) );
  DFFSRX2 dict_reg_24__2_ ( .D(n34723), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50821), .QN(n32598) );
  DFFSRX2 dict_reg_24__0_ ( .D(n34725), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50607), .QN(n32600) );
  DFFSRX2 dict_reg_23__3_ ( .D(n34714), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51034), .QN(n32589) );
  DFFSRX2 dict_reg_23__0_ ( .D(n34717), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50606), .QN(n32592) );
  DFFSRX2 dict_reg_22__3_ ( .D(n34706), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51033), .QN(n32581) );
  DFFSRX2 dict_reg_22__2_ ( .D(n34707), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50819), .QN(n32582) );
  DFFSRX2 dict_reg_22__0_ ( .D(n34709), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50605), .QN(n32584) );
  DFFSRX2 dict_reg_41__3_ ( .D(n34858), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51052), .QN(n32733) );
  DFFSRX2 dict_reg_41__2_ ( .D(n34859), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50838), .QN(n32734) );
  DFFSRX2 dict_reg_41__0_ ( .D(n34861), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50624), .QN(n32736) );
  DFFSRX2 dict_reg_42__3_ ( .D(n34866), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51053), .QN(n32741) );
  DFFSRX2 dict_reg_46__0_ ( .D(n34901), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50629), .QN(n32776) );
  DFFSRX2 dict_reg_42__2_ ( .D(n34867), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50839), .QN(n32742) );
  DFFSRX2 dict_reg_44__2_ ( .D(n34883), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50841), .QN(n32758) );
  DFFSRX2 dict_reg_44__0_ ( .D(n34885), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50627), .QN(n32760) );
  DFFSRX2 dict_reg_42__0_ ( .D(n34869), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50625), .QN(n32744) );
  DFFSRX2 dict_reg_252__1_ ( .D(n36548), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n41205), .QN(n34423) );
  DFFSRX2 data_num_reg_2_ ( .D(nxt_data_num[2]), .CK(clk), .SN(1'b1), .RN(
        n37590), .Q(n50147), .QN(n32398) );
  DFFSRX2 dict_reg_108__3_ ( .D(n35394), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51119), .QN(n33269) );
  DFFSRX2 dict_reg_220__0_ ( .D(n36293), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49152), .QN(n34168) );
  DFFSRX2 dict_reg_174__3_ ( .D(n35922), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51185), .QN(n33797) );
  DFFSRX2 dict_reg_174__2_ ( .D(n35923), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50971), .QN(n33798) );
  DFFSRX2 dict_reg_56__0_ ( .D(n34981), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50639), .QN(n32856) );
  DFFSRX2 dict_reg_15__3_ ( .D(n34650), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51026), .QN(n32525) );
  DFFSRX2 dict_reg_35__2_ ( .D(n34811), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50832), .QN(n32686) );
  DFFSRX2 dict_reg_35__0_ ( .D(n34813), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50618), .QN(n32688) );
  DFFSRX2 dict_reg_34__2_ ( .D(n34803), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50831), .QN(n32678) );
  DFFSRX2 dict_reg_34__0_ ( .D(n34805), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50617), .QN(n32680) );
  DFFSRX2 dict_reg_33__3_ ( .D(n34794), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51044), .QN(n32669) );
  DFFSRX2 dict_reg_31__2_ ( .D(n34779), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50828), .QN(n32654) );
  DFFSRX2 dict_reg_62__3_ ( .D(n35026), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51073), .QN(n32901) );
  DFFSRX2 dict_reg_62__2_ ( .D(n35027), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50859), .QN(n32902) );
  DFFSRX2 dict_reg_62__0_ ( .D(n35029), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50645), .QN(n32904) );
  DFFSRX2 dict_reg_61__3_ ( .D(n35018), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51072), .QN(n32893) );
  DFFSRX2 dict_reg_61__2_ ( .D(n35019), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50858), .QN(n32894) );
  DFFSRX2 dict_reg_61__0_ ( .D(n35021), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50644), .QN(n32896) );
  DFFSRX2 dict_reg_60__3_ ( .D(n35010), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51071), .QN(n32885) );
  DFFSRX2 dict_reg_60__2_ ( .D(n35011), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50857), .QN(n32886) );
  DFFSRX2 dict_reg_60__0_ ( .D(n35013), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50643), .QN(n32888) );
  DFFSRX2 dict_reg_59__3_ ( .D(n35002), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51070), .QN(n32877) );
  DFFSRX2 dict_reg_59__2_ ( .D(n35003), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50856), .QN(n32878) );
  DFFSRX2 dict_reg_58__3_ ( .D(n34994), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51069), .QN(n32869) );
  DFFSRX2 dict_reg_58__2_ ( .D(n34995), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50855), .QN(n32870) );
  DFFSRX2 dict_reg_57__3_ ( .D(n34986), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51068), .QN(n32861) );
  DFFSRX2 dict_reg_48__3_ ( .D(n34914), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51059), .QN(n32789) );
  DFFSRX2 dict_reg_48__2_ ( .D(n34915), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50845), .QN(n32790) );
  DFFSRX2 dict_reg_48__0_ ( .D(n34917), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50631), .QN(n32792) );
  DFFSRX2 dict_reg_47__0_ ( .D(n34909), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50630), .QN(n32784) );
  DFFSRX2 dict_reg_21__3_ ( .D(n34698), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51032), .QN(n32573) );
  DFFSRX2 dict_reg_20__3_ ( .D(n34690), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51031), .QN(n32565) );
  DFFSRX2 dict_reg_20__2_ ( .D(n34691), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50817), .QN(n32566) );
  DFFSRX2 dict_reg_20__0_ ( .D(n34693), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50603), .QN(n32568) );
  DFFSRX2 dict_reg_15__2_ ( .D(n34651), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50812), .QN(n32526) );
  DFFSRX2 dict_reg_15__0_ ( .D(n34653), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50598), .QN(n32528) );
  DFFSRX2 dict_reg_14__3_ ( .D(n34642), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51025), .QN(n32517) );
  DFFSRX2 dict_reg_14__2_ ( .D(n34643), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50811), .QN(n32518) );
  DFFSRX2 dict_reg_14__0_ ( .D(n34645), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50597), .QN(n32520) );
  DFFSRX2 dict_reg_13__2_ ( .D(n34635), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50810), .QN(n32510) );
  DFFSRX2 dict_reg_13__0_ ( .D(n34637), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50596), .QN(n32512) );
  DFFSRX2 dict_reg_17__7_ ( .D(n34662), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50397), .QN(n32537) );
  DFFSRX2 dict_reg_15__7_ ( .D(n34646), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50395), .QN(n32521) );
  DFFSRX2 dict_reg_32__7_ ( .D(n34782), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50412), .QN(n32657) );
  DFFSRX2 dict_reg_49__7_ ( .D(n34918), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50429), .QN(n32793) );
  DFFSRX2 dict_reg_63__3_ ( .D(n35034), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51074), .QN(n32909) );
  DFFSRX2 dict_reg_63__2_ ( .D(n35035), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50860), .QN(n32910) );
  DFFSRX2 dict_reg_63__0_ ( .D(n35037), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50646), .QN(n32912) );
  DFFSRX2 dict_reg_25__3_ ( .D(n34730), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51036), .QN(n32605) );
  DFFSRX2 dict_reg_25__2_ ( .D(n34731), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50822), .QN(n32606) );
  DFFSRX2 dict_reg_25__0_ ( .D(n34733), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50608), .QN(n32608) );
  DFFSRX2 dict_reg_23__2_ ( .D(n34715), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50820), .QN(n32590) );
  DFFSRX2 dict_reg_21__2_ ( .D(n34699), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50818), .QN(n32574) );
  DFFSRX2 dict_reg_21__0_ ( .D(n34701), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50604), .QN(n32576) );
  DFFSRX2 dict_reg_13__3_ ( .D(n34634), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51024), .QN(n32509) );
  DFFSRX2 dict_reg_12__3_ ( .D(n34626), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51023), .QN(n32501) );
  DFFSRX2 dict_reg_12__2_ ( .D(n34627), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50809), .QN(n32502) );
  DFFSRX2 dict_reg_12__0_ ( .D(n34629), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50595), .QN(n32504) );
  DFFSRX2 dict_reg_11__3_ ( .D(n34618), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51022), .QN(n32493) );
  DFFSRX2 dict_reg_11__2_ ( .D(n34619), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50808), .QN(n32494) );
  DFFSRX2 dict_reg_11__0_ ( .D(n34621), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50594), .QN(n32496) );
  DFFSRX2 dict_reg_10__3_ ( .D(n34610), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51021), .QN(n32485) );
  DFFSRX2 dict_reg_10__2_ ( .D(n34611), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50807), .QN(n32486) );
  DFFSRX2 dict_reg_10__0_ ( .D(n34613), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50593), .QN(n32488) );
  DFFSRX2 dict_reg_9__3_ ( .D(n34602), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51020), .QN(n32477) );
  DFFSRX2 dict_reg_9__2_ ( .D(n34603), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50806), .QN(n32478) );
  DFFSRX2 dict_reg_9__0_ ( .D(n34605), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50592), .QN(n32480) );
  DFFSRX2 dict_reg_8__3_ ( .D(n34594), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51019), .QN(n32469) );
  DFFSRX2 dict_reg_8__2_ ( .D(n34595), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50805), .QN(n32470) );
  DFFSRX2 dict_reg_8__0_ ( .D(n34597), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50591), .QN(n32472) );
  DFFSRX2 dict_reg_7__3_ ( .D(n34586), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51018), .QN(n32461) );
  DFFSRX2 dict_reg_7__2_ ( .D(n34587), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50804), .QN(n32462) );
  DFFSRX2 dict_reg_7__0_ ( .D(n34589), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50590), .QN(n32464) );
  DFFSRX2 dict_reg_6__3_ ( .D(n34578), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51017), .QN(n32453) );
  DFFSRX2 dict_reg_6__2_ ( .D(n34579), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50803), .QN(n32454) );
  DFFSRX2 dict_reg_6__0_ ( .D(n34581), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50589), .QN(n32456) );
  DFFSRX2 dict_reg_9__7_ ( .D(n34598), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50389), .QN(n32473) );
  DFFSRX2 dict_reg_8__7_ ( .D(n34590), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50388), .QN(n32465) );
  DFFSRX2 dict_reg_7__7_ ( .D(n34582), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50387), .QN(n32457) );
  DFFSRX2 dict_reg_31__7_ ( .D(n34774), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50411), .QN(n32649) );
  DFFSRX2 dict_reg_46__3_ ( .D(n34898), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51057), .QN(n32773) );
  DFFSRX2 dict_reg_46__2_ ( .D(n34899), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50843), .QN(n32774) );
  DFFSRX2 dict_reg_45__2_ ( .D(n34891), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50842), .QN(n32766) );
  DFFSRX2 dict_reg_45__0_ ( .D(n34893), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50628), .QN(n32768) );
  DFFSRX2 dict_reg_44__3_ ( .D(n34882), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51055), .QN(n32757) );
  DFFSRX2 dict_reg_109__0_ ( .D(n35405), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50692), .QN(n33280) );
  DFFSRX2 dict_reg_247__6_ ( .D(n36503), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49359), .QN(n34378) );
  DFFSRX2 dict_reg_247__0_ ( .D(n36509), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49047), .QN(n34384) );
  DFFSRX2 dict_reg_250__2_ ( .D(n36531), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n48884), .QN(n34406) );
  DFFSRX2 dict_reg_249__0_ ( .D(n36525), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49039), .QN(n34400) );
  DFFSRX2 dict_reg_248__2_ ( .D(n36515), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48891), .QN(n34390) );
  DFFSRX2 dict_reg_5__3_ ( .D(n34570), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51016), .QN(n32445) );
  DFFSRX2 dict_reg_5__2_ ( .D(n34571), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50802), .QN(n32446) );
  DFFSRX2 dict_reg_173__3_ ( .D(n35914), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51184), .QN(n33789) );
  DFFSRX2 dict_reg_173__0_ ( .D(n35917), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50756), .QN(n33792) );
  DFFSRX2 dict_reg_37__7_ ( .D(n34822), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50417), .QN(n32697) );
  DFFSRX2 dict_reg_36__7_ ( .D(n34814), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50416), .QN(n32689) );
  DFFSRX2 dict_reg_36__2_ ( .D(n34819), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50833), .QN(n32694) );
  DFFSRX2 dict_reg_35__7_ ( .D(n34806), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50415), .QN(n32681) );
  DFFSRX2 dict_reg_35__3_ ( .D(n34810), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51046), .QN(n32685) );
  DFFSRX2 dict_reg_34__3_ ( .D(n34802), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51045), .QN(n32677) );
  DFFSRX2 dict_reg_59__0_ ( .D(n35005), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50642), .QN(n32880) );
  DFFSRX2 dict_reg_58__0_ ( .D(n34997), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50641), .QN(n32872) );
  DFFSRX2 dict_reg_57__2_ ( .D(n34987), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50854), .QN(n32862) );
  DFFSRX2 dict_reg_57__0_ ( .D(n34989), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50640), .QN(n32864) );
  DFFSRX2 dict_reg_47__3_ ( .D(n34906), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51058), .QN(n32781) );
  DFFSRX2 dict_reg_47__2_ ( .D(n34907), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50844), .QN(n32782) );
  DFFSRX2 dict_reg_19__3_ ( .D(n34682), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51030), .QN(n32557) );
  DFFSRX2 dict_reg_19__2_ ( .D(n34683), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50816), .QN(n32558) );
  DFFSRX2 dict_reg_19__0_ ( .D(n34685), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50602), .QN(n32560) );
  DFFSRX2 dict_reg_33__7_ ( .D(n34790), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50413), .QN(n32665) );
  DFFSRX2 dict_reg_16__7_ ( .D(n34654), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50396), .QN(n32529) );
  DFFSRX2 dict_reg_48__7_ ( .D(n34910), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50428), .QN(n32785) );
  DFFSRX2 dict_reg_67__3_ ( .D(n35066), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51078), .QN(n32941) );
  DFFSRX2 dict_reg_67__2_ ( .D(n35067), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50864), .QN(n32942) );
  DFFSRX2 dict_reg_64__3_ ( .D(n35042), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51075), .QN(n32917) );
  DFFSRX2 dict_reg_64__2_ ( .D(n35043), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50861), .QN(n32918) );
  DFFSRX2 dict_reg_5__0_ ( .D(n34573), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50588), .QN(n32448) );
  DFFSRX2 dict_reg_40__3_ ( .D(n34850), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51051), .QN(n32725) );
  DFFSRX2 dict_reg_40__2_ ( .D(n34851), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50837), .QN(n32726) );
  DFFSRX2 dict_reg_40__0_ ( .D(n34853), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50623), .QN(n32728) );
  DFFSRX2 dict_reg_45__3_ ( .D(n34890), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51056), .QN(n32765) );
  DFFSRX2 dict_reg_38__2_ ( .D(n34835), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50835), .QN(n32710) );
  DFFSRX2 dict_reg_38__0_ ( .D(n34837), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50621), .QN(n32712) );
  DFFSRX2 dict_reg_37__2_ ( .D(n34827), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50834), .QN(n32702) );
  DFFSRX2 dict_reg_39__2_ ( .D(n34843), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50836), .QN(n32718) );
  DFFSRX2 dict_reg_39__0_ ( .D(n34845), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50622), .QN(n32720) );
  DFFSRX2 dict_reg_47__7_ ( .D(n34902), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50427), .QN(n32777) );
  DFFSRX2 dict_reg_108__2_ ( .D(n35395), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50905), .QN(n33270) );
  DFFSRX2 dict_reg_126__3_ ( .D(n35538), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51137), .QN(n33413) );
  DFFSRX2 dict_reg_126__2_ ( .D(n35539), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50923), .QN(n33414) );
  DFFSRX2 dict_reg_125__3_ ( .D(n35530), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51136), .QN(n33405) );
  DFFSRX2 dict_reg_125__2_ ( .D(n35531), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50922), .QN(n33406) );
  DFFSRX2 dict_reg_125__0_ ( .D(n35533), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50708), .QN(n33408) );
  DFFSRX2 dict_reg_238__6_ ( .D(n36431), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49395), .QN(n34306) );
  DFFSRX2 dict_reg_250__6_ ( .D(n36527), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49347), .QN(n34402) );
  DFFSRX2 dict_reg_217__0_ ( .D(n36269), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49164), .QN(n34144) );
  DFFSRX2 dict_reg_248__3_ ( .D(n36514), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48734), .QN(n34389) );
  DFFSRX2 dict_reg_237__0_ ( .D(n36429), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49086), .QN(n34304) );
  DFFSRX2 dict_reg_239__0_ ( .D(n36445), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49078), .QN(n34320) );
  DFFSRX2 dict_reg_245__3_ ( .D(n36490), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n48746), .QN(n34365) );
  DFFSRX2 dict_reg_245__2_ ( .D(n36491), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48902), .QN(n34366) );
  DFFSRX2 dict_reg_236__6_ ( .D(n36415), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49403), .QN(n34290) );
  DFFSRX2 dict_reg_4__3_ ( .D(n34562), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51015), .QN(n32437) );
  DFFSRX2 dict_reg_4__2_ ( .D(n34563), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50801), .QN(n32438) );
  DFFSRX2 dict_reg_4__0_ ( .D(n34565), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50587), .QN(n32440) );
  DFFSRX2 dict_reg_173__2_ ( .D(n35915), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50970), .QN(n33790) );
  DFFSRX2 dict_reg_37__3_ ( .D(n34826), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51048), .QN(n32701) );
  DFFSRX2 dict_reg_36__3_ ( .D(n34818), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51047), .QN(n32693) );
  DFFSRX2 dict_reg_36__0_ ( .D(n34821), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50619), .QN(n32696) );
  DFFSRX2 dict_reg_63__7_ ( .D(n35030), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50443), .QN(n32905) );
  DFFSRX2 dict_reg_34__7_ ( .D(n34798), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50414), .QN(n32673) );
  DFFSRX2 dict_reg_71__3_ ( .D(n35098), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51082), .QN(n32973) );
  DFFSRX2 dict_reg_71__2_ ( .D(n35099), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50868), .QN(n32974) );
  DFFSRX2 dict_reg_71__0_ ( .D(n35101), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50654), .QN(n32976) );
  DFFSRX2 dict_reg_73__0_ ( .D(n35117), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50656), .QN(n32992) );
  DFFSRX2 dict_reg_70__7_ ( .D(n35086), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50450), .QN(n32961) );
  DFFSRX2 dict_reg_70__3_ ( .D(n35090), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51081), .QN(n32965) );
  DFFSRX2 dict_reg_70__2_ ( .D(n35091), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50867), .QN(n32966) );
  DFFSRX2 dict_reg_69__2_ ( .D(n35083), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50866), .QN(n32958) );
  DFFSRX2 dict_reg_72__3_ ( .D(n35106), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51083), .QN(n32981) );
  DFFSRX2 dict_reg_72__2_ ( .D(n35107), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50869), .QN(n32982) );
  DFFSRX2 dict_reg_72__0_ ( .D(n35109), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50655), .QN(n32984) );
  DFFSRX2 dict_reg_69__7_ ( .D(n35078), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50449), .QN(n32953) );
  DFFSRX2 dict_reg_67__7_ ( .D(n35062), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50447), .QN(n32937) );
  DFFSRX2 dict_reg_66__3_ ( .D(n35058), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51077), .QN(n32933) );
  DFFSRX2 dict_reg_66__2_ ( .D(n35059), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50863), .QN(n32934) );
  DFFSRX2 dict_reg_65__3_ ( .D(n35050), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51076), .QN(n32925) );
  DFFSRX2 dict_reg_65__2_ ( .D(n35051), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50862), .QN(n32926) );
  DFFSRX2 dict_reg_65__7_ ( .D(n35046), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50445), .QN(n32921) );
  DFFSRX2 dict_reg_66__7_ ( .D(n35054), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50446), .QN(n32929) );
  DFFSRX2 dict_reg_64__7_ ( .D(n35038), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50444), .QN(n32913) );
  DFFSRX2 dict_reg_2__3_ ( .D(n34546), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51013), .QN(n32421) );
  DFFSRX2 dict_reg_2__2_ ( .D(n34547), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50799), .QN(n32422) );
  DFFSRX2 dict_reg_2__0_ ( .D(n34549), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50585), .QN(n32424) );
  DFFSRX2 dict_reg_39__3_ ( .D(n34842), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51050), .QN(n32717) );
  DFFSRX2 dict_reg_38__7_ ( .D(n34830), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50418), .QN(n32705) );
  DFFSRX2 dict_reg_38__3_ ( .D(n34834), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51049), .QN(n32709) );
  DFFSRX2 dict_reg_37__0_ ( .D(n34829), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50620), .QN(n32704) );
  DFFSRX2 dict_reg_95__2_ ( .D(n35291), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50892), .QN(n33166) );
  DFFSRX2 dict_reg_109__3_ ( .D(n35402), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51120), .QN(n33277) );
  DFFSRX2 dict_reg_109__2_ ( .D(n35403), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50906), .QN(n33278) );
  DFFSRX2 dict_reg_100__0_ ( .D(n35333), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50683), .QN(n33208) );
  DFFSRX2 dict_reg_95__3_ ( .D(n35290), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51106), .QN(n33165) );
  DFFSRX2 dict_reg_95__0_ ( .D(n35293), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50678), .QN(n33168) );
  DFFSRX2 dict_reg_108__0_ ( .D(n35397), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50691), .QN(n33272) );
  DFFSRX2 dict_reg_110__0_ ( .D(n35413), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50693), .QN(n33288) );
  DFFSRX2 dict_reg_110__3_ ( .D(n35410), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51121), .QN(n33285) );
  DFFSRX2 dict_reg_110__2_ ( .D(n35411), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50907), .QN(n33286) );
  DFFSRX2 dict_reg_225__6_ ( .D(n36327), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n49446), .QN(n34202) );
  DFFSRX2 dict_reg_1__0_ ( .D(n34541), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50584), .QN(n32416) );
  DFFSRX2 dict_reg_1__2_ ( .D(n34539), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50798), .QN(n32414) );
  DFFSRX2 dict_reg_1__7_ ( .D(n34534), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50381), .QN(n32409) );
  DFFSRX2 dict_reg_243__0_ ( .D(n36477), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49062), .QN(n34352) );
  DFFSRX2 dict_reg_236__0_ ( .D(n36421), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49090), .QN(n34296) );
  DFFSRX2 dict_reg_235__0_ ( .D(n36413), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49094), .QN(n34288) );
  DFFSRX2 dict_reg_238__0_ ( .D(n36437), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49082), .QN(n34312) );
  DFFSRX2 dict_reg_239__3_ ( .D(n36442), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48770), .QN(n34317) );
  DFFSRX2 dict_reg_221__0_ ( .D(n36301), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49148), .QN(n34176) );
  DFFSRX2 dict_reg_247__3_ ( .D(n36506), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48738), .QN(n34381) );
  DFFSRX2 dict_reg_247__2_ ( .D(n36507), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n48895), .QN(n34382) );
  DFFSRX2 dict_reg_243__3_ ( .D(n36474), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48754), .QN(n34349) );
  DFFSRX2 dict_reg_3__2_ ( .D(n34555), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50800), .QN(n32430) );
  DFFSRX2 dict_reg_3__3_ ( .D(n34554), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51014), .QN(n32429) );
  DFFSRX2 dict_reg_3__0_ ( .D(n34557), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50586), .QN(n32432) );
  DFFSRX2 dict_reg_76__3_ ( .D(n35138), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51087), .QN(n33013) );
  DFFSRX2 dict_reg_76__0_ ( .D(n35141), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50659), .QN(n33016) );
  DFFSRX2 dict_reg_74__0_ ( .D(n35125), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50657), .QN(n33000) );
  DFFSRX2 dict_reg_74__3_ ( .D(n35122), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51085), .QN(n32997) );
  DFFSRX2 dict_reg_74__2_ ( .D(n35123), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50871), .QN(n32998) );
  DFFSRX2 dict_reg_73__3_ ( .D(n35114), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51084), .QN(n32989) );
  DFFSRX2 dict_reg_73__2_ ( .D(n35115), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50870), .QN(n32990) );
  DFFSRX2 dict_reg_70__0_ ( .D(n35093), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50653), .QN(n32968) );
  DFFSRX2 dict_reg_69__0_ ( .D(n35085), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50652), .QN(n32960) );
  DFFSRX2 dict_reg_69__3_ ( .D(n35082), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51080), .QN(n32957) );
  DFFSRX2 dict_reg_68__7_ ( .D(n35070), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50448), .QN(n32945) );
  DFFSRX2 dict_reg_68__3_ ( .D(n35074), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51079), .QN(n32949) );
  DFFSRX2 dict_reg_68__2_ ( .D(n35075), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50865), .QN(n32950) );
  DFFSRX2 dict_reg_68__0_ ( .D(n35077), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50651), .QN(n32952) );
  DFFSRX2 dict_reg_67__0_ ( .D(n35069), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50650), .QN(n32944) );
  DFFSRX2 dict_reg_66__0_ ( .D(n35061), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50649), .QN(n32936) );
  DFFSRX2 dict_reg_65__0_ ( .D(n35053), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50648), .QN(n32928) );
  DFFSRX2 dict_reg_64__0_ ( .D(n35045), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50647), .QN(n32920) );
  DFFSRX2 dict_reg_76__2_ ( .D(n35139), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50873), .QN(n33014) );
  DFFSRX2 dict_reg_75__2_ ( .D(n35131), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50872), .QN(n33006) );
  DFFSRX2 dict_reg_75__3_ ( .D(n35130), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51086), .QN(n33005) );
  DFFSRX2 dict_reg_75__0_ ( .D(n35133), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50658), .QN(n33008) );
  DFFSRX2 dict_reg_96__3_ ( .D(n35298), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51107), .QN(n33173) );
  DFFSRX2 dict_reg_96__2_ ( .D(n35299), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50893), .QN(n33174) );
  DFFSRX2 dict_reg_96__0_ ( .D(n35301), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50679), .QN(n33176) );
  DFFSRX2 dict_reg_107__3_ ( .D(n35386), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51118), .QN(n33261) );
  DFFSRX2 dict_reg_107__2_ ( .D(n35387), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50904), .QN(n33262) );
  DFFSRX2 dict_reg_107__0_ ( .D(n35389), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50690), .QN(n33264) );
  DFFSRX2 dict_reg_106__3_ ( .D(n35378), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51117), .QN(n33253) );
  DFFSRX2 dict_reg_106__2_ ( .D(n35379), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50903), .QN(n33254) );
  DFFSRX2 dict_reg_106__0_ ( .D(n35381), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50689), .QN(n33256) );
  DFFSRX2 dict_reg_105__3_ ( .D(n35370), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51116), .QN(n33245) );
  DFFSRX2 dict_reg_105__2_ ( .D(n35371), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50902), .QN(n33246) );
  DFFSRX2 dict_reg_105__0_ ( .D(n35373), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50688), .QN(n33248) );
  DFFSRX2 dict_reg_104__3_ ( .D(n35362), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51115), .QN(n33237) );
  DFFSRX2 dict_reg_104__2_ ( .D(n35363), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50901), .QN(n33238) );
  DFFSRX2 dict_reg_104__0_ ( .D(n35365), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50687), .QN(n33240) );
  DFFSRX2 dict_reg_103__3_ ( .D(n35354), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51114), .QN(n33229) );
  DFFSRX2 dict_reg_103__2_ ( .D(n35355), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50900), .QN(n33230) );
  DFFSRX2 dict_reg_102__3_ ( .D(n35346), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51113), .QN(n33221) );
  DFFSRX2 dict_reg_102__2_ ( .D(n35347), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50899), .QN(n33222) );
  DFFSRX2 dict_reg_102__0_ ( .D(n35349), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50685), .QN(n33224) );
  DFFSRX2 dict_reg_101__3_ ( .D(n35338), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51112), .QN(n33213) );
  DFFSRX2 dict_reg_101__2_ ( .D(n35339), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50898), .QN(n33214) );
  DFFSRX2 dict_reg_101__0_ ( .D(n35341), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50684), .QN(n33216) );
  DFFSRX2 dict_reg_99__3_ ( .D(n35322), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51110), .QN(n33197) );
  DFFSRX2 dict_reg_99__2_ ( .D(n35323), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50896), .QN(n33198) );
  DFFSRX2 dict_reg_99__0_ ( .D(n35325), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50682), .QN(n33200) );
  DFFSRX2 dict_reg_100__3_ ( .D(n35330), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51111), .QN(n33205) );
  DFFSRX2 dict_reg_100__2_ ( .D(n35331), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50897), .QN(n33206) );
  DFFSRX2 dict_reg_97__3_ ( .D(n35306), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51108), .QN(n33181) );
  DFFSRX2 dict_reg_97__2_ ( .D(n35307), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50894), .QN(n33182) );
  DFFSRX2 dict_reg_97__0_ ( .D(n35309), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50680), .QN(n33184) );
  DFFSRX2 dict_reg_98__3_ ( .D(n35314), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51109), .QN(n33189) );
  DFFSRX2 dict_reg_98__2_ ( .D(n35315), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50895), .QN(n33190) );
  DFFSRX2 dict_reg_98__0_ ( .D(n35317), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50681), .QN(n33192) );
  DFFSRX2 dict_reg_103__0_ ( .D(n35357), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50686), .QN(n33232) );
  DFFSRX2 dict_reg_95__7_ ( .D(n35286), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50466), .QN(n33161) );
  DFFSRX2 dict_reg_97__7_ ( .D(n35302), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50468), .QN(n33177) );
  DFFSRX2 dict_reg_96__7_ ( .D(n35294), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50467), .QN(n33169) );
  DFFSRX2 dict_reg_98__7_ ( .D(n35310), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50469), .QN(n33185) );
  DFFSRX2 dict_reg_228__0_ ( .D(n36357), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49122), .QN(n34232) );
  DFFSRX2 dict_reg_246__3_ ( .D(n36498), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48742), .QN(n34373) );
  DFFSRX2 dict_reg_246__7_ ( .D(n36494), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49208), .QN(n34369) );
  DFFSRX2 dict_reg_244__6_ ( .D(n36479), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49371), .QN(n34354) );
  DFFSRX2 dict_reg_1__3_ ( .D(n34538), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51012), .QN(n32413) );
  DFFSRX2 dict_reg_244__0_ ( .D(n36485), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49058), .QN(n34360) );
  DFFSRX2 dict_reg_246__4_ ( .D(n36497), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n48583), .QN(n34372) );
  DFFSRX2 dict_reg_237__3_ ( .D(n36426), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48778), .QN(n34301) );
  DFFSRX2 dict_reg_250__3_ ( .D(n36530), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48726), .QN(n34405) );
  DFFSRX2 dict_reg_250__4_ ( .D(n36529), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48568), .QN(n34404) );
  DFFSRX2 dict_reg_242__7_ ( .D(n36462), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49224), .QN(n34337) );
  DFFSRX2 dict_reg_226__2_ ( .D(n36339), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n48978), .QN(n34214) );
  DFFSRX2 dict_reg_233__0_ ( .D(n36397), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49102), .QN(n34272) );
  DFFSRX2 dict_reg_234__0_ ( .D(n36405), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49098), .QN(n34280) );
  DFFSRX2 dict_reg_242__3_ ( .D(n36466), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48758), .QN(n34341) );
  DFFSRX2 dict_reg_239__2_ ( .D(n36443), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n48926), .QN(n34318) );
  DFFSRX2 dict_reg_245__7_ ( .D(n36486), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49212), .QN(n34361) );
  DFFSRX2 dict_reg_222__6_ ( .D(n36303), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49458), .QN(n34178) );
  DFFSRX2 dict_reg_237__6_ ( .D(n36423), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49399), .QN(n34298) );
  DFFSRX2 dict_reg_232__7_ ( .D(n36382), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49264), .QN(n34257) );
  DFFSRX2 dict_reg_232__6_ ( .D(n36383), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n49419), .QN(n34258) );
  DFFSRX2 dict_reg_237__7_ ( .D(n36422), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49244), .QN(n34297) );
  DFFSRX2 dict_reg_236__7_ ( .D(n36414), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n49248), .QN(n34289) );
  DFFSRX2 dict_reg_237__4_ ( .D(n36425), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48618), .QN(n34300) );
  DFFSRX2 dict_reg_220__6_ ( .D(n36287), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49466), .QN(n34162) );
  DFFSRX2 dict_reg_239__6_ ( .D(n36439), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49391), .QN(n34314) );
  DFFSRX2 dict_reg_247__4_ ( .D(n36505), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n48579), .QN(n34380) );
  DFFSRX2 dict_reg_242__0_ ( .D(n36469), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49066), .QN(n34344) );
  DFFSRX2 dict_reg_244__7_ ( .D(n36478), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49216), .QN(n34353) );
  DFFSRX2 dict_reg_246__6_ ( .D(n36495), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49363), .QN(n34370) );
  DFFSRX2 dict_reg_238__7_ ( .D(n36430), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49240), .QN(n34305) );
  DFFSRX2 dict_reg_244__3_ ( .D(n36482), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n48750), .QN(n34357) );
  DFFSRX2 dict_reg_239__4_ ( .D(n36441), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48610), .QN(n34316) );
  DFFSRX2 dict_reg_236__4_ ( .D(n36417), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48622), .QN(n34292) );
  DFFSRX2 dict_reg_234__7_ ( .D(n36398), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49256), .QN(n34273) );
  DFFSRX2 dict_reg_228__4_ ( .D(n36353), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48654), .QN(n34228) );
  DFFSRX2 dict_reg_245__6_ ( .D(n36487), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49367), .QN(n34362) );
  DFFSRX2 dict_reg_240__2_ ( .D(n36451), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48922), .QN(n34326) );
  DFFSRX2 dict_reg_241__7_ ( .D(n36454), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49228), .QN(n34329) );
  DFFSRX2 dict_reg_244__4_ ( .D(n36481), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n48590), .QN(n34356) );
  DFFSRX2 dict_reg_250__7_ ( .D(n36526), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49192), .QN(n34401) );
  DFFSRX2 dict_reg_218__2_ ( .D(n36275), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49010), .QN(n34150) );
  DFFSRX2 dict_reg_219__0_ ( .D(n36285), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49156), .QN(n34160) );
  DFFSRX2 dict_reg_231__0_ ( .D(n36381), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49110), .QN(n34256) );
  DFFSRX2 dict_reg_227__0_ ( .D(n36349), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49126), .QN(n34224) );
  DFFSRX2 dict_reg_223__0_ ( .D(n36317), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49141), .QN(n34192) );
  DFFSRX2 dict_reg_238__3_ ( .D(n36434), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n48774), .QN(n34309) );
  DFFSRX2 dict_reg_238__4_ ( .D(n36433), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48614), .QN(n34308) );
  DFFSRX2 dict_reg_239__7_ ( .D(n36438), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49236), .QN(n34313) );
  DFFSRX2 dict_reg_233__4_ ( .D(n36393), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48634), .QN(n34268) );
  DFFSRX2 dict_reg_226__0_ ( .D(n36341), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49130), .QN(n34216) );
  DFFSRX2 dict_reg_247__7_ ( .D(n36502), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49204), .QN(n34377) );
  DFFSRX2 dict_reg_248__7_ ( .D(n36510), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49200), .QN(n34385) );
  DFFSRX2 dict_reg_229__0_ ( .D(n36365), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49118), .QN(n34240) );
  DFFSRX2 dict_reg_248__4_ ( .D(n36513), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48575), .QN(n34388) );
  DFFSRX2 dict_reg_248__0_ ( .D(n36517), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49043), .QN(n34392) );
  DFFSRX2 dict_reg_242__6_ ( .D(n36463), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49379), .QN(n34338) );
  DFFSRX2 dict_reg_215__0_ ( .D(n36253), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49171), .QN(n34128) );
  DFFSRX2 dict_reg_226__7_ ( .D(n36334), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49288), .QN(n34209) );
  DFFSRX2 dict_reg_240__6_ ( .D(n36447), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49387), .QN(n34322) );
  DFFSRX2 dict_reg_222__7_ ( .D(n36302), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49303), .QN(n34177) );
  DFFSRX2 dict_reg_222__2_ ( .D(n36307), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n48994), .QN(n34182) );
  DFFSRX2 dict_reg_238__2_ ( .D(n36435), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48930), .QN(n34310) );
  DFFSRX2 dict_reg_220__7_ ( .D(n36286), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49311), .QN(n34161) );
  DFFSRX2 dict_reg_220__2_ ( .D(n36291), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49002), .QN(n34166) );
  DFFSRX2 dict_reg_221__2_ ( .D(n36299), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48998), .QN(n34174) );
  DFFSRX2 dict_reg_218__6_ ( .D(n36271), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49474), .QN(n34146) );
  DFFSRX2 dict_reg_218__7_ ( .D(n36270), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49319), .QN(n34145) );
  DFFSRX2 dict_reg_223__7_ ( .D(n36310), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49299), .QN(n34185) );
  DFFSRX2 dict_reg_236__3_ ( .D(n36418), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48782), .QN(n34293) );
  DFFSRX2 dict_reg_235__3_ ( .D(n36410), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48786), .QN(n34285) );
  DFFSRX2 dict_reg_219__7_ ( .D(n36278), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n49315), .QN(n34153) );
  DFFSRX2 dict_reg_240__3_ ( .D(n36450), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48766), .QN(n34325) );
  DFFSRX2 dict_reg_235__7_ ( .D(n36406), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49252), .QN(n34281) );
  DFFSRX2 dict_reg_233__7_ ( .D(n36390), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49260), .QN(n34265) );
  DFFSRX2 dict_reg_233__3_ ( .D(n36394), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n48794), .QN(n34269) );
  DFFSRX2 dict_reg_230__4_ ( .D(n36369), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48646), .QN(n34244) );
  DFFSRX2 dict_reg_229__2_ ( .D(n36363), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48966), .QN(n34238) );
  DFFSRX2 dict_reg_228__2_ ( .D(n36355), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48970), .QN(n34230) );
  DFFSRX2 dict_reg_227__4_ ( .D(n36345), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48658), .QN(n34220) );
  DFFSRX2 dict_reg_227__2_ ( .D(n36347), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48974), .QN(n34222) );
  DFFSRX2 dict_reg_225__4_ ( .D(n36329), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n48666), .QN(n34204) );
  DFFSRX2 dict_reg_219__4_ ( .D(n36281), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n48690), .QN(n34156) );
  DFFSRX2 dict_reg_224__6_ ( .D(n36319), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n49450), .QN(n34194) );
  DFFSRX2 dict_reg_236__2_ ( .D(n36419), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48938), .QN(n34294) );
  DFFSRX2 dict_reg_232__2_ ( .D(n36387), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48954), .QN(n34262) );
  DFFSRX2 dict_reg_231__2_ ( .D(n36379), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48958), .QN(n34254) );
  DFFSRX2 dict_reg_229__4_ ( .D(n36361), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48650), .QN(n34236) );
  DFFSRX2 dict_reg_224__7_ ( .D(n36318), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49295), .QN(n34193) );
  DFFSRX2 dict_reg_243__7_ ( .D(n36470), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49220), .QN(n34345) );
  DFFSRX2 dict_reg_241__3_ ( .D(n36458), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48762), .QN(n34333) );
  DFFSRX2 dict_reg_241__6_ ( .D(n36455), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n49383), .QN(n34330) );
  DFFSRX2 dict_reg_218__4_ ( .D(n36273), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48694), .QN(n34148) );
  DFFSRX2 dict_reg_217__4_ ( .D(n36265), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48698), .QN(n34140) );
  DFFSRX2 dict_reg_242__4_ ( .D(n36465), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48598), .QN(n34340) );
  DFFSRX2 dict_reg_243__4_ ( .D(n36473), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48594), .QN(n34348) );
  DFFSRX2 dict_reg_232__0_ ( .D(n36389), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49106), .QN(n34264) );
  DFFSRX2 dict_reg_218__0_ ( .D(n36277), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n49160), .QN(n34152) );
  DFFSRX2 dict_reg_241__0_ ( .D(n36461), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49070), .QN(n34336) );
  DFFSRX2 dict_reg_226__6_ ( .D(n36335), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49442), .QN(n34210) );
  DFFSRX2 dict_reg_230__7_ ( .D(n36366), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49272), .QN(n34241) );
  DFFSRX2 dict_reg_222__3_ ( .D(n36306), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n48838), .QN(n34181) );
  DFFSRX2 dict_reg_222__4_ ( .D(n36305), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n48678), .QN(n34180) );
  DFFSRX2 dict_reg_237__2_ ( .D(n36427), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48934), .QN(n34302) );
  DFFSRX2 dict_reg_221__7_ ( .D(n36294), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49307), .QN(n34169) );
  DFFSRX2 dict_reg_220__4_ ( .D(n36289), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48686), .QN(n34164) );
  DFFSRX2 dict_reg_220__3_ ( .D(n36290), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48846), .QN(n34165) );
  DFFSRX2 dict_reg_234__6_ ( .D(n36399), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49411), .QN(n34274) );
  DFFSRX2 dict_reg_229__7_ ( .D(n36358), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49276), .QN(n34233) );
  DFFSRX2 dict_reg_221__3_ ( .D(n36298), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48842), .QN(n34173) );
  DFFSRX2 dict_reg_223__6_ ( .D(n36311), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49454), .QN(n34186) );
  DFFSRX2 dict_reg_217__6_ ( .D(n36263), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49478), .QN(n34138) );
  DFFSRX2 dict_reg_221__6_ ( .D(n36295), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49462), .QN(n34170) );
  DFFSRX2 dict_reg_219__6_ ( .D(n36279), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49470), .QN(n34154) );
  DFFSRX2 dict_reg_219__2_ ( .D(n36283), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49006), .QN(n34158) );
  DFFSRX2 dict_reg_241__2_ ( .D(n36459), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48918), .QN(n34334) );
  DFFSRX2 dict_reg_235__6_ ( .D(n36407), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49407), .QN(n34282) );
  DFFSRX2 dict_reg_235__4_ ( .D(n36409), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48626), .QN(n34284) );
  DFFSRX2 dict_reg_234__3_ ( .D(n36402), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n48790), .QN(n34277) );
  DFFSRX2 dict_reg_234__2_ ( .D(n36403), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48946), .QN(n34278) );
  DFFSRX2 dict_reg_233__6_ ( .D(n36391), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49415), .QN(n34266) );
  DFFSRX2 dict_reg_232__3_ ( .D(n36386), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48798), .QN(n34261) );
  DFFSRX2 dict_reg_231__7_ ( .D(n36374), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49268), .QN(n34249) );
  DFFSRX2 dict_reg_231__6_ ( .D(n36375), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49423), .QN(n34250) );
  DFFSRX2 dict_reg_231__3_ ( .D(n36378), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48802), .QN(n34253) );
  DFFSRX2 dict_reg_230__3_ ( .D(n36370), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n48806), .QN(n34245) );
  DFFSRX2 dict_reg_229__3_ ( .D(n36362), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48810), .QN(n34237) );
  DFFSRX2 dict_reg_228__3_ ( .D(n36354), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n48814), .QN(n34229) );
  DFFSRX2 dict_reg_227__6_ ( .D(n36343), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49438), .QN(n34218) );
  DFFSRX2 dict_reg_227__3_ ( .D(n36346), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48818), .QN(n34221) );
  DFFSRX2 dict_reg_226__4_ ( .D(n36337), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48662), .QN(n34212) );
  DFFSRX2 dict_reg_226__3_ ( .D(n36338), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n48822), .QN(n34213) );
  DFFSRX2 dict_reg_225__3_ ( .D(n36330), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n48826), .QN(n34205) );
  DFFSRX2 dict_reg_224__4_ ( .D(n36321), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48670), .QN(n34196) );
  DFFSRX2 dict_reg_224__3_ ( .D(n36322), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n48830), .QN(n34197) );
  DFFSRX2 dict_reg_223__3_ ( .D(n36314), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n48834), .QN(n34189) );
  DFFSRX2 dict_reg_223__2_ ( .D(n36315), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n48990), .QN(n34190) );
  DFFSRX2 dict_reg_219__3_ ( .D(n36282), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48850), .QN(n34157) );
  DFFSRX2 dict_reg_242__2_ ( .D(n36467), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48914), .QN(n34342) );
  DFFSRX2 dict_reg_235__2_ ( .D(n36411), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n48942), .QN(n34286) );
  DFFSRX2 dict_reg_233__2_ ( .D(n36395), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48950), .QN(n34270) );
  DFFSRX2 dict_reg_231__4_ ( .D(n36377), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n48642), .QN(n34252) );
  DFFSRX2 dict_reg_228__7_ ( .D(n36350), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49280), .QN(n34225) );
  DFFSRX2 dict_reg_228__6_ ( .D(n36351), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49434), .QN(n34226) );
  DFFSRX2 dict_reg_227__7_ ( .D(n36342), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49284), .QN(n34217) );
  DFFSRX2 dict_reg_225__2_ ( .D(n36331), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n48982), .QN(n34206) );
  DFFSRX2 dict_reg_224__2_ ( .D(n36323), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n48986), .QN(n34198) );
  DFFSRX2 dict_reg_223__4_ ( .D(n36313), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48674), .QN(n34188) );
  DFFSRX2 dict_reg_232__4_ ( .D(n36385), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n48638), .QN(n34260) );
  DFFSRX2 dict_reg_230__2_ ( .D(n36371), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48962), .QN(n34246) );
  DFFSRX2 dict_reg_221__4_ ( .D(n36297), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n48682), .QN(n34172) );
  DFFSRX2 dict_reg_229__6_ ( .D(n36359), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n49430), .QN(n34234) );
  DFFSRX2 dict_reg_215__4_ ( .D(n36249), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n48705), .QN(n34124) );
  DFFSRX2 dict_reg_215__3_ ( .D(n36250), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n48864), .QN(n34125) );
  DFFSRX2 dict_reg_218__3_ ( .D(n36274), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n48854), .QN(n34149) );
  DFFSRX2 dict_reg_241__4_ ( .D(n36457), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n48602), .QN(n34332) );
  DFFSRX2 dict_reg_234__4_ ( .D(n36401), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n48630), .QN(n34276) );
  DFFSRX2 dict_reg_243__6_ ( .D(n36471), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n49375), .QN(n34346) );
  DFFSRX2 dict_reg_30__4_ ( .D(n34769), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51255), .QN(n32644) );
  DFFSRX2 dict_reg_53__4_ ( .D(n34953), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51278), .QN(n32828) );
  DFFSRX2 dict_reg_52__4_ ( .D(n34945), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51277), .QN(n32820) );
  DFFSRX2 dict_reg_51__4_ ( .D(n34937), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51276), .QN(n32812) );
  DFFSRX2 dict_reg_55__4_ ( .D(n34969), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51280), .QN(n32844) );
  DFFSRX2 dict_reg_54__4_ ( .D(n34961), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51279), .QN(n32836) );
  DFFSRX2 dict_reg_50__4_ ( .D(n34929), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51275), .QN(n32804) );
  DFFSRX2 dict_reg_26__4_ ( .D(n34737), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51251), .QN(n32612) );
  DFFSRX2 dict_reg_42__7_ ( .D(n34862), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50422), .QN(n32737) );
  DFFSRX2 dict_reg_43__4_ ( .D(n34873), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51268), .QN(n32748) );
  DFFSRX2 dict_reg_56__4_ ( .D(n34977), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51281), .QN(n32852) );
  DFFSRX2 dict_reg_10__7_ ( .D(n34606), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50390), .QN(n32481) );
  DFFSRX2 dict_reg_6__7_ ( .D(n34574), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50386), .QN(n32449) );
  DFFSRX2 dict_reg_28__4_ ( .D(n34753), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51253), .QN(n32628) );
  DFFSRX2 dict_reg_27__4_ ( .D(n34745), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51252), .QN(n32620) );
  DFFSRX2 dict_reg_46__4_ ( .D(n34897), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51271), .QN(n32772) );
  DFFSRX2 dict_reg_44__4_ ( .D(n34881), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51269), .QN(n32756) );
  DFFSRX2 dict_reg_5__7_ ( .D(n34566), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50385), .QN(n32441) );
  DFFSRX2 dict_reg_19__4_ ( .D(n34681), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51244), .QN(n32556) );
  DFFSRX2 dict_reg_62__4_ ( .D(n35025), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51287), .QN(n32900) );
  DFFSRX2 dict_reg_61__4_ ( .D(n35017), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51286), .QN(n32892) );
  DFFSRX2 dict_reg_60__4_ ( .D(n35009), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51285), .QN(n32884) );
  DFFSRX2 dict_reg_59__4_ ( .D(n35001), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51284), .QN(n32876) );
  DFFSRX2 dict_reg_58__4_ ( .D(n34993), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51283), .QN(n32868) );
  DFFSRX2 dict_reg_57__4_ ( .D(n34985), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51282), .QN(n32860) );
  DFFSRX2 dict_reg_18__7_ ( .D(n34670), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50398), .QN(n32545) );
  DFFSRX2 dict_reg_14__4_ ( .D(n34641), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51239), .QN(n32516) );
  DFFSRX2 dict_reg_72__4_ ( .D(n35105), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51297), .QN(n32980) );
  DFFSRX2 dict_reg_13__4_ ( .D(n34633), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51238), .QN(n32508) );
  DFFSRX2 dict_reg_12__4_ ( .D(n34625), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51237), .QN(n32500) );
  DFFSRX2 dict_reg_11__4_ ( .D(n34617), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51236), .QN(n32492) );
  DFFSRX2 dict_reg_23__4_ ( .D(n34713), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51248), .QN(n32588) );
  DFFSRX2 dict_reg_29__4_ ( .D(n34761), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51254), .QN(n32636) );
  DFFSRX2 dict_reg_25__4_ ( .D(n34729), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51250), .QN(n32604) );
  DFFSRX2 dict_reg_24__4_ ( .D(n34721), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51249), .QN(n32596) );
  DFFSRX2 dict_reg_22__4_ ( .D(n34705), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51247), .QN(n32580) );
  DFFSRX2 dict_reg_41__7_ ( .D(n34854), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50421), .QN(n32729) );
  DFFSRX2 dict_reg_40__7_ ( .D(n34846), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50420), .QN(n32721) );
  DFFSRX2 dict_reg_45__4_ ( .D(n34889), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51270), .QN(n32764) );
  DFFSRX2 dict_reg_126__4_ ( .D(n35537), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51350), .QN(n33412) );
  DFFSRX2 dict_reg_110__4_ ( .D(n35409), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51334), .QN(n33284) );
  DFFSRX2 dict_reg_3__7_ ( .D(n34550), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50383), .QN(n32425) );
  DFFSRX2 dict_reg_4__7_ ( .D(n34558), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50384), .QN(n32433) );
  DFFSRX2 dict_reg_174__4_ ( .D(n35921), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51398), .QN(n33796) );
  DFFSRX2 dict_reg_173__4_ ( .D(n35913), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51397), .QN(n33788) );
  DFFSRX2 dict_reg_20__4_ ( .D(n34689), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51245), .QN(n32564) );
  DFFSRX2 dict_reg_21__4_ ( .D(n34697), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51246), .QN(n32572) );
  DFFSRX2 dict_reg_73__4_ ( .D(n35113), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51298), .QN(n32988) );
  DFFSRX2 dict_reg_2__7_ ( .D(n34542), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50382), .QN(n32417) );
  DFFSRX2 dict_reg_39__7_ ( .D(n34838), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50419), .QN(n32713) );
  DFFSRX2 dict_reg_109__4_ ( .D(n35401), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51333), .QN(n33276) );
  DFFSRX2 dict_reg_125__4_ ( .D(n35529), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51349), .QN(n33404) );
  DFFSRX2 dict_reg_209__7_ ( .D(n36198), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50578), .QN(n34073) );
  DFFSRX2 dict_reg_0__0_ ( .D(n34533), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50583), .QN(n32408) );
  DFFSRX2 dict_reg_0__3_ ( .D(n34530), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51011), .QN(n32405) );
  DFFSRX2 dict_reg_0__2_ ( .D(n34531), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50797), .QN(n32406) );
  DFFSRX2 dict_reg_74__4_ ( .D(n35121), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51299), .QN(n32996) );
  DFFSRX2 dict_reg_102__4_ ( .D(n35345), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51326), .QN(n33220) );
  DFFSRX2 dict_reg_101__4_ ( .D(n35337), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51325), .QN(n33212) );
  DFFSRX2 dict_reg_99__4_ ( .D(n35321), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51323), .QN(n33196) );
  DFFSRX2 dict_reg_100__4_ ( .D(n35329), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51324), .QN(n33204) );
  DFFSRX2 dict_reg_103__4_ ( .D(n35353), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51327), .QN(n33228) );
  DFFSRX2 dict_reg_107__4_ ( .D(n35385), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51331), .QN(n33260) );
  DFFSRX2 dict_reg_108__4_ ( .D(n35393), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51332), .QN(n33268) );
  DFFSRX2 dict_reg_106__4_ ( .D(n35377), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51330), .QN(n33252) );
  DFFSRX2 dict_reg_105__4_ ( .D(n35369), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51329), .QN(n33244) );
  DFFSRX2 dict_reg_104__4_ ( .D(n35361), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51328), .QN(n33236) );
  DFFSRX2 dict_reg_71__4_ ( .D(n35097), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51296), .QN(n32972) );
  DFFSRX2 dict_reg_0__7_ ( .D(n34526), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50380), .QN(n32401) );
  DFFSRX1 dict_reg_215__6_ ( .D(n36247), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n49510), .QN(n34122) );
  DFFSRX1 dict_reg_215__2_ ( .D(n36251), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n49515), .QN(n34126) );
  DFFSRX1 dict_reg_215__7_ ( .D(n36246), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49512), .QN(n34121) );
  DFFSRX1 dict_reg_253__1_ ( .D(n36556), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n34431) );
  DFFRX2 dict_reg_189__0_ ( .D(n36045), .CK(clk), .RN(n42360), .Q(n50772),
        .QN(n33920) );
  DFFRX2 dict_reg_145__7_ ( .D(n35686), .CK(clk), .RN(n42344), .Q(n50514),
        .QN(n33561) );
  DFFRX2 dict_reg_174__0_ ( .D(n35925), .CK(clk), .RN(n42358), .Q(n50757),
        .QN(n33800) );
  DFFSRX1 dict_reg_252__4_ ( .D(n36545), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48561), .QN(n34420) );
  DFFRX2 dict_reg_145__3_ ( .D(n35690), .CK(clk), .RN(n42393), .Q(n51156),
        .QN(n33565) );
  DFFRX2 dict_reg_171__2_ ( .D(n35899), .CK(clk), .RN(n42383), .Q(n50968),
        .QN(n33774) );
  DFFRX2 dict_reg_171__3_ ( .D(n35898), .CK(clk), .RN(n42395), .Q(n51182),
        .QN(n33773) );
  DFFSRX1 dict_reg_253__5_ ( .D(n36552), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n34427) );
  DFFSRX1 dict_reg_172__6_ ( .D(n35903), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50337), .QN(n33778) );
  DFFSRX1 dict_reg_30__7_ ( .D(n34766), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50410), .QN(n32641) );
  DFFSRX1 dict_reg_53__7_ ( .D(n34950), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50433), .QN(n32825) );
  DFFSRX1 dict_reg_52__7_ ( .D(n34942), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50432), .QN(n32817) );
  DFFSRX1 dict_reg_51__7_ ( .D(n34934), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50431), .QN(n32809) );
  DFFSRX1 dict_reg_14__7_ ( .D(n34638), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50394), .QN(n32513) );
  DFFSRX1 dict_reg_55__7_ ( .D(n34966), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50435), .QN(n32841) );
  DFFSRX1 dict_reg_54__7_ ( .D(n34958), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50434), .QN(n32833) );
  DFFSRX1 dict_reg_50__7_ ( .D(n34926), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50430), .QN(n32801) );
  DFFSRX1 dict_reg_56__7_ ( .D(n34974), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50436), .QN(n32849) );
  DFFSRX1 dict_reg_13__7_ ( .D(n34630), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50393), .QN(n32505) );
  DFFSRX1 dict_reg_12__7_ ( .D(n34622), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50392), .QN(n32497) );
  DFFSRX1 dict_reg_11__7_ ( .D(n34614), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50391), .QN(n32489) );
  DFFSRX1 dict_reg_22__7_ ( .D(n34702), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50402), .QN(n32577) );
  DFFSRX1 dict_reg_27__7_ ( .D(n34742), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50407), .QN(n32617) );
  DFFSRX1 dict_reg_29__7_ ( .D(n34758), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50409), .QN(n32633) );
  DFFSRX1 dict_reg_28__7_ ( .D(n34750), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50408), .QN(n32625) );
  DFFSRX1 dict_reg_24__7_ ( .D(n34718), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50404), .QN(n32593) );
  DFFSRX1 dict_reg_6__4_ ( .D(n34577), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51231), .QN(n32452) );
  DFFSRX1 dict_reg_26__7_ ( .D(n34734), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50406), .QN(n32609) );
  DFFSRX1 dict_reg_44__7_ ( .D(n34878), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50424), .QN(n32753) );
  DFFSRX1 dict_reg_43__7_ ( .D(n34870), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50423), .QN(n32745) );
  DFFSRX1 dict_reg_174__7_ ( .D(n35918), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50543), .QN(n33793) );
  DFFSRX1 dict_reg_156__7_ ( .D(n35774), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50525), .QN(n33649) );
  DFFSRX1 dict_reg_252__7_ ( .D(n36542), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n49185), .QN(n34417) );
  DFFSRX1 dict_reg_155__7_ ( .D(n35766), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50524), .QN(n33641) );
  DFFSRX1 dict_reg_204__6_ ( .D(n36159), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50369), .QN(n34034) );
  DFFSRX1 dict_reg_79__6_ ( .D(n35159), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50244), .QN(n33034) );
  DFFSRX1 dict_reg_101__6_ ( .D(n35335), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50266), .QN(n33210) );
  DFFSRX1 dict_reg_107__6_ ( .D(n35383), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50272), .QN(n33258) );
  DFFSRX1 dict_reg_106__6_ ( .D(n35375), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50271), .QN(n33250) );
  DFFSRX1 dict_reg_102__6_ ( .D(n35343), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50267), .QN(n33218) );
  DFFSRX1 dict_reg_110__6_ ( .D(n35407), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50275), .QN(n33282) );
  DFFSRX1 dict_reg_100__6_ ( .D(n35327), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50265), .QN(n33202) );
  DFFSRX1 dict_reg_96__6_ ( .D(n35295), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50261), .QN(n33170) );
  DFFSRX1 dict_reg_95__6_ ( .D(n35287), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50260), .QN(n33162) );
  DFFSRX1 dict_reg_116__6_ ( .D(n35455), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50281), .QN(n33330) );
  DFFSRX1 dict_reg_91__6_ ( .D(n35255), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50256), .QN(n33130) );
  DFFSRX1 dict_reg_85__6_ ( .D(n35207), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50250), .QN(n33082) );
  DFFSRX1 dict_reg_77__6_ ( .D(n35143), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50242), .QN(n33018) );
  DFFSRX1 dict_reg_153__6_ ( .D(n35751), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50318), .QN(n33626) );
  DFFSRX1 dict_reg_154__6_ ( .D(n35759), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50319), .QN(n33634) );
  DFFSRX1 dict_reg_185__6_ ( .D(n36007), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50350), .QN(n33882) );
  DFFSRX1 dict_reg_152__6_ ( .D(n35743), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50317), .QN(n33618) );
  DFFSRX1 dict_reg_186__6_ ( .D(n36015), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50351), .QN(n33890) );
  DFFSRX1 dict_reg_108__6_ ( .D(n35391), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50273), .QN(n33266) );
  DFFSRX1 dict_reg_205__6_ ( .D(n36167), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50370), .QN(n34042) );
  DFFSRX1 dict_reg_195__6_ ( .D(n36087), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50360), .QN(n33962) );
  DFFSRX1 dict_reg_206__6_ ( .D(n36175), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50371), .QN(n34050) );
  DFFSRX1 dict_reg_200__6_ ( .D(n36127), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50365), .QN(n34002) );
  DFFSRX1 dict_reg_156__6_ ( .D(n35775), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50321), .QN(n33650) );
  DFFSRX1 dict_reg_21__7_ ( .D(n34694), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50401), .QN(n32569) );
  DFFSRX1 dict_reg_57__7_ ( .D(n34982), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50437), .QN(n32857) );
  DFFSRX1 dict_reg_18__4_ ( .D(n34673), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51243), .QN(n32548) );
  DFFSRX1 dict_reg_2__4_ ( .D(n34545), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51227), .QN(n32420) );
  DFFSRX1 dict_reg_23__7_ ( .D(n34710), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50403), .QN(n32585) );
  DFFSRX1 dict_reg_25__7_ ( .D(n34726), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50405), .QN(n32601) );
  DFFSRX1 dict_reg_10__4_ ( .D(n34609), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51235), .QN(n32484) );
  DFFSRX1 dict_reg_41__4_ ( .D(n34857), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51266), .QN(n32732) );
  DFFSRX1 dict_reg_42__4_ ( .D(n34865), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51267), .QN(n32740) );
  DFFSRX1 dict_reg_46__7_ ( .D(n34894), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50426), .QN(n32769) );
  DFFSRX1 dict_reg_45__7_ ( .D(n34886), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50425), .QN(n32761) );
  DFFSRX1 dict_reg_71__7_ ( .D(n35094), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50451), .QN(n32969) );
  DFFSRX1 dict_reg_151__7_ ( .D(n35734), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50520), .QN(n33609) );
  DFFSRX1 dict_reg_152__7_ ( .D(n35742), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50521), .QN(n33617) );
  DFFSRX1 dict_reg_189__7_ ( .D(n36038), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50558), .QN(n33913) );
  DFFSRX1 dict_reg_187__7_ ( .D(n36022), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50556), .QN(n33897) );
  DFFSRX1 dict_reg_181__7_ ( .D(n35974), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50550), .QN(n33849) );
  DFFSRX1 dict_reg_149__7_ ( .D(n35718), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50518), .QN(n33593) );
  DFFSRX1 dict_reg_148__7_ ( .D(n35710), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50517), .QN(n33585) );
  DFFSRX1 dict_reg_206__7_ ( .D(n36174), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50575), .QN(n34049) );
  DFFSRX1 dict_reg_205__7_ ( .D(n36166), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50574), .QN(n34041) );
  DFFSRX1 dict_reg_204__7_ ( .D(n36158), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50573), .QN(n34033) );
  DFFSRX1 dict_reg_209__4_ ( .D(n36201), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51433), .QN(n34076) );
  DFFSRX1 dict_reg_172__7_ ( .D(n35902), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50541), .QN(n33777) );
  DFFSRX1 dict_reg_170__7_ ( .D(n35886), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50539), .QN(n33761) );
  DFFSRX1 dict_reg_173__6_ ( .D(n35911), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50338), .QN(n33786) );
  DFFSRX1 dict_reg_105__6_ ( .D(n35367), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50270), .QN(n33242) );
  DFFSRX1 dict_reg_98__6_ ( .D(n35311), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50263), .QN(n33186) );
  DFFSRX1 dict_reg_93__6_ ( .D(n35271), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50258), .QN(n33146) );
  DFFSRX1 dict_reg_92__6_ ( .D(n35263), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50257), .QN(n33138) );
  DFFSRX1 dict_reg_136__6_ ( .D(n35615), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50301), .QN(n33490) );
  DFFSRX1 dict_reg_35__6_ ( .D(n34807), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50200), .QN(n32682) );
  DFFSRX1 dict_reg_33__6_ ( .D(n34791), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50198), .QN(n32666) );
  DFFSRX1 dict_reg_50__6_ ( .D(n34927), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50215), .QN(n32802) );
  DFFSRX1 dict_reg_52__6_ ( .D(n34943), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50217), .QN(n32818) );
  DFFSRX1 dict_reg_51__6_ ( .D(n34935), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50216), .QN(n32810) );
  DFFSRX1 dict_reg_140__6_ ( .D(n35647), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50305), .QN(n33522) );
  DFFSRX1 dict_reg_138__6_ ( .D(n35631), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50303), .QN(n33506) );
  DFFSRX1 dict_reg_103__6_ ( .D(n35351), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50268), .QN(n33226) );
  DFFSRX1 dict_reg_150__6_ ( .D(n35727), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50315), .QN(n33602) );
  DFFSRX1 dict_reg_208__6_ ( .D(n36191), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50373), .QN(n34066) );
  DFFSRX1 dict_reg_160__6_ ( .D(n35807), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50325), .QN(n33682) );
  DFFSRX1 dict_reg_158__6_ ( .D(n35791), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50323), .QN(n33666) );
  DFFSRX1 dict_reg_134__6_ ( .D(n35599), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50299), .QN(n33474) );
  DFFSRX1 dict_reg_207__6_ ( .D(n36183), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50372), .QN(n34058) );
  DFFSRX1 dict_reg_170__6_ ( .D(n35887), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50335), .QN(n33762) );
  DFFSRX1 dict_reg_169__6_ ( .D(n35879), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50334), .QN(n33754) );
  DFFSRX1 dict_reg_175__6_ ( .D(n35927), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50340), .QN(n33802) );
  DFFSRX1 dict_reg_191__4_ ( .D(n36057), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51415), .QN(n33932) );
  DFFSRX1 dict_reg_159__4_ ( .D(n35801), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51383), .QN(n33676) );
  DFFSRX1 dict_reg_125__6_ ( .D(n35527), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50290), .QN(n33402) );
  DFFSRX1 dict_reg_120__6_ ( .D(n35487), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50285), .QN(n33362) );
  DFFSRX1 dict_reg_78__6_ ( .D(n35151), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50243), .QN(n33026) );
  DFFSRX1 dict_reg_84__6_ ( .D(n35199), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50249), .QN(n33074) );
  DFFSRX1 dict_reg_80__6_ ( .D(n35167), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50245), .QN(n33042) );
  DFFSRX1 dict_reg_94__6_ ( .D(n35279), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50259), .QN(n33154) );
  DFFSRX1 dict_reg_141__6_ ( .D(n35655), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50306), .QN(n33530) );
  DFFSRX1 dict_reg_128__6_ ( .D(n35551), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50293), .QN(n33426) );
  DFFSRX1 dict_reg_130__6_ ( .D(n35567), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50295), .QN(n33442) );
  DFFSRX1 dict_reg_165__6_ ( .D(n35847), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50330), .QN(n33722) );
  DFFSRX1 dict_reg_184__6_ ( .D(n35999), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50349), .QN(n33874) );
  DFFSRX1 dict_reg_119__6_ ( .D(n35479), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50284), .QN(n33354) );
  DFFSRX1 dict_reg_87__6_ ( .D(n35223), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50252), .QN(n33098) );
  DFFSRX1 dict_reg_112__6_ ( .D(n35423), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50277), .QN(n33298) );
  DFFSRX1 dict_reg_86__6_ ( .D(n35215), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50251), .QN(n33090) );
  DFFSRX1 dict_reg_111__6_ ( .D(n35415), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50276), .QN(n33290) );
  DFFSRX1 dict_reg_139__6_ ( .D(n35639), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50304), .QN(n33514) );
  DFFSRX1 dict_reg_196__6_ ( .D(n36095), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50361), .QN(n33970) );
  DFFSRX1 dict_reg_5__4_ ( .D(n34569), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51230), .QN(n32444) );
  DFFSRX1 dict_reg_3__4_ ( .D(n34553), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51228), .QN(n32428) );
  DFFSRX1 dict_reg_20__7_ ( .D(n34686), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50400), .QN(n32561) );
  DFFSRX1 dict_reg_19__7_ ( .D(n34678), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50399), .QN(n32553) );
  DFFSRX1 dict_reg_61__7_ ( .D(n35014), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50441), .QN(n32889) );
  DFFSRX1 dict_reg_59__7_ ( .D(n34998), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50439), .QN(n32873) );
  DFFSRX1 dict_reg_58__7_ ( .D(n34990), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50438), .QN(n32865) );
  DFFSRX1 dict_reg_60__7_ ( .D(n35006), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50440), .QN(n32881) );
  DFFSRX1 dict_reg_62__7_ ( .D(n35022), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50442), .QN(n32897) );
  DFFSRX1 dict_reg_72__7_ ( .D(n35102), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50452), .QN(n32977) );
  DFFSRX1 dict_reg_126__7_ ( .D(n35534), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50495), .QN(n33409) );
  DFFSRX1 dict_reg_108__7_ ( .D(n35390), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50479), .QN(n33265) );
  DFFSRX1 dict_reg_109__7_ ( .D(n35398), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50480), .QN(n33273) );
  DFFSRX1 dict_reg_153__7_ ( .D(n35750), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50522), .QN(n33625) );
  DFFSRX1 dict_reg_154__7_ ( .D(n35758), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50523), .QN(n33633) );
  DFFSRX1 dict_reg_182__7_ ( .D(n35982), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50551), .QN(n33857) );
  DFFSRX1 dict_reg_178__7_ ( .D(n35950), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50547), .QN(n33825) );
  DFFSRX1 dict_reg_188__7_ ( .D(n36030), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50557), .QN(n33905) );
  DFFSRX1 dict_reg_186__7_ ( .D(n36014), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50555), .QN(n33889) );
  DFFSRX1 dict_reg_157__7_ ( .D(n35782), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50526), .QN(n33657) );
  DFFSRX1 dict_reg_150__7_ ( .D(n35726), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50519), .QN(n33601) );
  DFFSRX1 dict_reg_184__7_ ( .D(n35998), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50553), .QN(n33873) );
  DFFSRX1 dict_reg_180__7_ ( .D(n35966), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50549), .QN(n33841) );
  DFFSRX1 dict_reg_179__7_ ( .D(n35958), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50548), .QN(n33833) );
  DFFSRX1 dict_reg_147__7_ ( .D(n35702), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50516), .QN(n33577) );
  DFFSRX1 dict_reg_210__7_ ( .D(n36206), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50579), .QN(n34081) );
  DFFSRX1 dict_reg_211__7_ ( .D(n36214), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50580), .QN(n34089) );
  DFFSRX1 dict_reg_201__7_ ( .D(n36134), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50570), .QN(n34009) );
  DFFSRX1 dict_reg_200__7_ ( .D(n36126), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50569), .QN(n34001) );
  DFFSRX1 dict_reg_202__7_ ( .D(n36142), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50571), .QN(n34017) );
  DFFSRX1 dict_reg_199__7_ ( .D(n36118), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50568), .QN(n33993) );
  DFFSRX1 dict_reg_173__7_ ( .D(n35910), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50542), .QN(n33785) );
  DFFSRX1 dict_reg_171__7_ ( .D(n35894), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50540), .QN(n33769) );
  DFFSRX1 dict_reg_190__7_ ( .D(n36046), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50559), .QN(n33921) );
  DFFSRX1 dict_reg_169__7_ ( .D(n35878), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50538), .QN(n33753) );
  DFFSRX1 dict_reg_168__7_ ( .D(n35870), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50537), .QN(n33745) );
  DFFSRX1 dict_reg_118__6_ ( .D(n35471), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50283), .QN(n33346) );
  DFFSRX1 dict_reg_188__6_ ( .D(n36031), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50353), .QN(n33906) );
  DFFSRX1 dict_reg_252__6_ ( .D(n36543), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n49340), .QN(n34418) );
  DFFSRX1 dict_reg_32__6_ ( .D(n34783), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50197), .QN(n32658) );
  DFFSRX1 dict_reg_149__6_ ( .D(n35719), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50314), .QN(n33594) );
  DFFSRX1 dict_reg_201__6_ ( .D(n36135), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50366), .QN(n34010) );
  DFFSRX1 dict_reg_197__6_ ( .D(n36103), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50362), .QN(n33978) );
  DFFSRX1 dict_reg_155__6_ ( .D(n35767), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50320), .QN(n33642) );
  DFFSRX1 dict_reg_113__6_ ( .D(n35431), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50278), .QN(n33306) );
  DFFSRX1 dict_reg_133__6_ ( .D(n35591), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50298), .QN(n33466) );
  DFFSRX1 dict_reg_171__6_ ( .D(n35895), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50336), .QN(n33770) );
  DFFSRX1 dict_reg_174__6_ ( .D(n35919), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50339), .QN(n33794) );
  DFFSRX1 dict_reg_157__6_ ( .D(n35783), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50322), .QN(n33658) );
  DFFSRX1 dict_reg_96__4_ ( .D(n35297), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51320), .QN(n33172) );
  DFFSRX1 dict_reg_112__4_ ( .D(n35425), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51336), .QN(n33300) );
  DFFSRX1 dict_reg_90__6_ ( .D(n35247), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50255), .QN(n33122) );
  DFFSRX1 dict_reg_76__6_ ( .D(n35135), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50241), .QN(n33010) );
  DFFSRX1 dict_reg_202__6_ ( .D(n36143), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50367), .QN(n34018) );
  DFFSRX1 dict_reg_181__6_ ( .D(n35975), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50346), .QN(n33850) );
  DFFSRX1 dict_reg_193__6_ ( .D(n36071), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50358), .QN(n33946) );
  DFFSRX1 dict_reg_163__6_ ( .D(n35831), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50328), .QN(n33706) );
  DFFSRX1 dict_reg_115__6_ ( .D(n35447), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50280), .QN(n33322) );
  DFFSRX1 dict_reg_34__6_ ( .D(n34799), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50199), .QN(n32674) );
  DFFSRX1 dict_reg_37__6_ ( .D(n34823), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50202), .QN(n32698) );
  DFFSRX1 dict_reg_60__6_ ( .D(n35007), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50225), .QN(n32882) );
  DFFSRX1 dict_reg_19__6_ ( .D(n34679), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50184), .QN(n32554) );
  DFFSRX1 dict_reg_18__6_ ( .D(n34671), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50183), .QN(n32546) );
  DFFSRX1 dict_reg_62__6_ ( .D(n35023), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50227), .QN(n32898) );
  DFFSRX1 dict_reg_61__6_ ( .D(n35015), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50226), .QN(n32890) );
  DFFSRX1 dict_reg_53__6_ ( .D(n34951), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50218), .QN(n32826) );
  DFFSRX1 dict_reg_20__6_ ( .D(n34687), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50185), .QN(n32562) );
  DFFSRX1 dict_reg_55__6_ ( .D(n34967), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50220), .QN(n32842) );
  DFFSRX1 dict_reg_63__6_ ( .D(n35031), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50228), .QN(n32906) );
  DFFSRX1 dict_reg_25__6_ ( .D(n34727), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50190), .QN(n32602) );
  DFFSRX1 dict_reg_28__6_ ( .D(n34751), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50193), .QN(n32626) );
  DFFSRX1 dict_reg_24__6_ ( .D(n34719), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50189), .QN(n32594) );
  DFFSRX1 dict_reg_42__6_ ( .D(n34863), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50207), .QN(n32738) );
  DFFSRX1 dict_reg_41__6_ ( .D(n34855), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50206), .QN(n32730) );
  DFFSRX1 dict_reg_43__6_ ( .D(n34871), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50208), .QN(n32746) );
  DFFSRX1 dict_reg_210__6_ ( .D(n36207), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50375), .QN(n34082) );
  DFFSRX1 dict_reg_26__6_ ( .D(n34735), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50191), .QN(n32610) );
  DFFSRX1 dict_reg_97__6_ ( .D(n35303), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50262), .QN(n33178) );
  DFFSRX1 dict_reg_89__6_ ( .D(n35239), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50254), .QN(n33114) );
  DFFSRX1 dict_reg_117__6_ ( .D(n35463), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50282), .QN(n33338) );
  DFFSRX1 dict_reg_167__6_ ( .D(n35863), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50332), .QN(n33738) );
  DFFSRX1 dict_reg_183__6_ ( .D(n35991), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50348), .QN(n33866) );
  DFFSRX1 dict_reg_99__6_ ( .D(n35319), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50264), .QN(n33194) );
  DFFSRX1 dict_reg_122__6_ ( .D(n35503), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50287), .QN(n33378) );
  DFFSRX1 dict_reg_81__6_ ( .D(n35175), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50246), .QN(n33050) );
  DFFSRX1 dict_reg_146__6_ ( .D(n35695), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50311), .QN(n33570) );
  DFFSRX1 dict_reg_36__6_ ( .D(n34815), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50201), .QN(n32690) );
  DFFSRX1 dict_reg_121__6_ ( .D(n35495), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50286), .QN(n33370) );
  DFFSRX1 dict_reg_187__6_ ( .D(n36023), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50352), .QN(n33898) );
  DFFSRX1 dict_reg_148__6_ ( .D(n35711), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50313), .QN(n33586) );
  DFFSRX1 dict_reg_27__6_ ( .D(n34743), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50192), .QN(n32618) );
  DFFSRX1 dict_reg_129__6_ ( .D(n35559), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50294), .QN(n33434) );
  DFFSRX1 dict_reg_4__4_ ( .D(n34561), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51229), .QN(n32436) );
  DFFSRX1 dict_reg_39__4_ ( .D(n34841), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51264), .QN(n32716) );
  DFFSRX1 dict_reg_40__4_ ( .D(n34849), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51265), .QN(n32724) );
  DFFSRX1 dict_reg_102__7_ ( .D(n35342), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50473), .QN(n33217) );
  DFFSRX1 dict_reg_101__7_ ( .D(n35334), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50472), .QN(n33209) );
  DFFSRX1 dict_reg_99__7_ ( .D(n35318), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50470), .QN(n33193) );
  DFFSRX1 dict_reg_110__7_ ( .D(n35406), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50481), .QN(n33281) );
  DFFSRX1 dict_reg_107__7_ ( .D(n35382), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50478), .QN(n33257) );
  DFFSRX1 dict_reg_105__7_ ( .D(n35366), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50476), .QN(n33241) );
  DFFSRX1 dict_reg_103__7_ ( .D(n35350), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50474), .QN(n33225) );
  DFFSRX1 dict_reg_106__7_ ( .D(n35374), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50477), .QN(n33249) );
  DFFSRX1 dict_reg_104__7_ ( .D(n35358), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50475), .QN(n33233) );
  DFFSRX1 dict_reg_100__7_ ( .D(n35326), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50471), .QN(n33201) );
  DFFSRX1 dict_reg_115__7_ ( .D(n35446), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50486), .QN(n33321) );
  DFFSRX1 dict_reg_118__7_ ( .D(n35470), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50488), .QN(n33345) );
  DFFSRX1 dict_reg_183__7_ ( .D(n35990), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50552), .QN(n33865) );
  DFFSRX1 dict_reg_185__7_ ( .D(n36006), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50554), .QN(n33881) );
  DFFSRX1 dict_reg_158__7_ ( .D(n35790), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50527), .QN(n33665) );
  DFFSRX1 dict_reg_139__7_ ( .D(n35638), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50508), .QN(n33513) );
  DFFSRX1 dict_reg_142__7_ ( .D(n35662), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50511), .QN(n33537) );
  DFFSRX1 dict_reg_141__7_ ( .D(n35654), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50510), .QN(n33529) );
  DFFSRX1 dict_reg_140__7_ ( .D(n35646), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50509), .QN(n33521) );
  DFFSRX1 dict_reg_213__7_ ( .D(n36230), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50582), .QN(n34105) );
  DFFSRX1 dict_reg_203__7_ ( .D(n36150), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50572), .QN(n34025) );
  DFFSRX1 dict_reg_212__7_ ( .D(n36222), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50581), .QN(n34097) );
  DFFSRX1 dict_reg_167__7_ ( .D(n35862), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50536), .QN(n33737) );
  DFFSRX1 dict_reg_109__6_ ( .D(n35399), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50274), .QN(n33274) );
  DFFSRX1 dict_reg_104__6_ ( .D(n35359), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50269), .QN(n33234) );
  DFFSRX1 dict_reg_88__6_ ( .D(n35231), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50253), .QN(n33106) );
  DFFSRX1 dict_reg_189__6_ ( .D(n36039), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50354), .QN(n33914) );
  DFFSRX1 dict_reg_209__6_ ( .D(n36199), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50374), .QN(n34074) );
  DFFSRX1 dict_reg_180__6_ ( .D(n35967), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50345), .QN(n33842) );
  DFFSRX1 dict_reg_178__6_ ( .D(n35951), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50343), .QN(n33826) );
  DFFSRX1 dict_reg_137__6_ ( .D(n35623), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50302), .QN(n33498) );
  DFFSRX1 dict_reg_179__6_ ( .D(n35959), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50344), .QN(n33834) );
  DFFSRX1 dict_reg_161__6_ ( .D(n35815), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50326), .QN(n33690) );
  DFFSRX1 dict_reg_162__6_ ( .D(n35823), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50327), .QN(n33698) );
  DFFSRX1 dict_reg_191__6_ ( .D(n36055), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50356), .QN(n33930) );
  DFFSRX1 dict_reg_159__6_ ( .D(n35799), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50324), .QN(n33674) );
  DFFSRX1 dict_reg_54__6_ ( .D(n34959), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50219), .QN(n32834) );
  DFFSRX1 dict_reg_5__6_ ( .D(n34567), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50170), .QN(n32442) );
  DFFSRX1 dict_reg_182__6_ ( .D(n35983), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50347), .QN(n33858) );
  DFFSRX1 dict_reg_145__6_ ( .D(n35687), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50310), .QN(n33562) );
  DFFSRX1 dict_reg_144__6_ ( .D(n35679), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50309), .QN(n33554) );
  DFFSRX1 dict_reg_194__4_ ( .D(n36081), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51418), .QN(n33956) );
  DFFSRX1 dict_reg_95__4_ ( .D(n35289), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51319), .QN(n33164) );
  DFFSRX1 dict_reg_132__4_ ( .D(n35585), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51356), .QN(n33460) );
  DFFSRX1 dict_reg_195__4_ ( .D(n36089), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51419), .QN(n33964) );
  DFFSRX1 dict_reg_190__6_ ( .D(n36047), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50355), .QN(n33922) );
  DFFSRX1 dict_reg_97__4_ ( .D(n35305), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51321), .QN(n33180) );
  DFFSRX1 dict_reg_98__4_ ( .D(n35313), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51322), .QN(n33188) );
  DFFSRX1 dict_reg_113__4_ ( .D(n35433), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51337), .QN(n33308) );
  DFFSRX1 dict_reg_111__4_ ( .D(n35417), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51335), .QN(n33292) );
  DFFSRX1 dict_reg_207__4_ ( .D(n36185), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51431), .QN(n34060) );
  DFFSRX1 dict_reg_177__4_ ( .D(n35945), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51401), .QN(n33820) );
  DFFSRX1 dict_reg_196__4_ ( .D(n36097), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51420), .QN(n33972) );
  DFFSRX1 dict_reg_164__4_ ( .D(n35841), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51388), .QN(n33716) );
  DFFSRX1 dict_reg_124__6_ ( .D(n35519), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50289), .QN(n33394) );
  DFFSRX1 dict_reg_132__6_ ( .D(n35583), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50297), .QN(n33458) );
  DFFSRX1 dict_reg_31__4_ ( .D(n34777), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51256), .QN(n32652) );
  DFFSRX1 dict_reg_143__4_ ( .D(n35673), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51367), .QN(n33548) );
  DFFSRX1 dict_reg_4__6_ ( .D(n34559), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50169), .QN(n32434) );
  DFFSRX1 dict_reg_13__6_ ( .D(n34631), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50178), .QN(n32506) );
  DFFSRX1 dict_reg_12__6_ ( .D(n34623), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50177), .QN(n32498) );
  DFFSRX1 dict_reg_114__6_ ( .D(n35439), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50279), .QN(n33314) );
  DFFSRX1 data_queue_reg_5__7_ ( .D(n36596), .CK(clk), .SN(1'b1), .RN(n37594),
        .QN(n34475) );
  DFFSRX1 data_queue_reg_5__6_ ( .D(n36595), .CK(clk), .SN(1'b1), .RN(n37593),
        .QN(n34476) );
  DFFSRX1 data_queue_reg_5__5_ ( .D(n36594), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n34477) );
  DFFSRX1 data_queue_reg_5__4_ ( .D(n36593), .CK(clk), .SN(1'b1), .RN(n37590),
        .QN(n34478) );
  DFFSRX1 data_queue_reg_5__3_ ( .D(n36592), .CK(clk), .SN(1'b1), .RN(n37596),
        .QN(n34479) );
  DFFSRX1 data_queue_reg_5__2_ ( .D(n36591), .CK(clk), .SN(1'b1), .RN(n37590),
        .QN(n34480) );
  DFFSRX1 data_queue_reg_5__1_ ( .D(n36590), .CK(clk), .SN(1'b1), .RN(n37591),
        .QN(n34481) );
  DFFSRX1 data_queue_reg_5__0_ ( .D(n36589), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n34482) );
  DFFSRX1 dict_reg_31__6_ ( .D(n34775), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50196), .QN(n32650) );
  DFFSRX1 dict_reg_49__6_ ( .D(n34919), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50214), .QN(n32794) );
  DFFSRX1 dict_reg_48__6_ ( .D(n34911), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50213), .QN(n32786) );
  DFFSRX1 dict_reg_59__6_ ( .D(n34999), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50224), .QN(n32874) );
  DFFSRX1 dict_reg_58__6_ ( .D(n34991), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50223), .QN(n32866) );
  DFFSRX1 dict_reg_47__6_ ( .D(n34903), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50212), .QN(n32778) );
  DFFSRX1 dict_reg_17__6_ ( .D(n34663), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50182), .QN(n32538) );
  DFFSRX1 dict_reg_16__6_ ( .D(n34655), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50181), .QN(n32530) );
  DFFSRX1 dict_reg_40__6_ ( .D(n34847), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50205), .QN(n32722) );
  DFFSRX1 dict_reg_127__6_ ( .D(n35543), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50292), .QN(n33418) );
  DFFSRX1 dict_reg_131__6_ ( .D(n35575), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50296), .QN(n33450) );
  DFFSRX1 dict_reg_147__6_ ( .D(n35703), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50312), .QN(n33578) );
  DFFSRX1 dict_reg_30__6_ ( .D(n34767), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50195), .QN(n32642) );
  DFFSRX1 dict_reg_75__6_ ( .D(n35127), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50240), .QN(n33002) );
  DFFSRX1 dict_reg_38__6_ ( .D(n34831), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50203), .QN(n32706) );
  DFFSRX1 dict_reg_123__6_ ( .D(n35511), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50288), .QN(n33386) );
  DFFSRX1 dict_reg_135__6_ ( .D(n35607), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50300), .QN(n33482) );
  DFFSRX1 dict_reg_29__6_ ( .D(n34759), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50194), .QN(n32634) );
  DFFSRX1 dict_reg_176__6_ ( .D(n35935), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50341), .QN(n33810) );
  DFFSRX1 dict_reg_212__6_ ( .D(n36223), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50377), .QN(n34098) );
  DFFSRX1 dict_reg_198__4_ ( .D(n36113), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51422), .QN(n33988) );
  DFFSRX1 dict_reg_166__4_ ( .D(n35857), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51390), .QN(n33732) );
  DFFSRX1 dict_reg_146__4_ ( .D(n35697), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51370), .QN(n33572) );
  DFFSRX1 dict_reg_144__4_ ( .D(n35681), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51368), .QN(n33556) );
  DFFSRX1 dict_reg_145__4_ ( .D(n35689), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51369), .QN(n33564) );
  DFFSRX1 dict_reg_83__6_ ( .D(n35191), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50248), .QN(n33066) );
  DFFSRX1 dict_reg_198__6_ ( .D(n36111), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50363), .QN(n33986) );
  DFFSRX1 dict_reg_166__6_ ( .D(n35855), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50331), .QN(n33730) );
  DFFSRX1 dict_reg_3__6_ ( .D(n34551), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50168), .QN(n32426) );
  DFFSRX1 dict_reg_70__6_ ( .D(n35087), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50235), .QN(n32962) );
  DFFSRX1 dict_reg_69__6_ ( .D(n35079), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50234), .QN(n32954) );
  DFFSRX1 dict_reg_65__6_ ( .D(n35047), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50230), .QN(n32922) );
  DFFSRX1 dict_reg_11__6_ ( .D(n34615), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50176), .QN(n32490) );
  DFFSRX1 dict_reg_71__6_ ( .D(n35095), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50236), .QN(n32970) );
  DFFSRX1 dict_reg_7__6_ ( .D(n34583), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50172), .QN(n32458) );
  DFFSRX1 dict_reg_74__6_ ( .D(n35119), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50239), .QN(n32994) );
  DFFSRX1 dict_reg_203__6_ ( .D(n36151), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50368), .QN(n34026) );
  DFFSRX1 dict_reg_126__6_ ( .D(n35535), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50291), .QN(n33410) );
  DFFSRX1 dict_reg_164__6_ ( .D(n35839), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50329), .QN(n33714) );
  DFFSRX1 data_queue_reg_7__0_ ( .D(n36573), .CK(clk), .SN(1'b1), .RN(n37595),
        .QN(n34498) );
  DFFSRX1 data_queue_reg_7__7_ ( .D(n36580), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n34491) );
  DFFSRX1 data_queue_reg_7__6_ ( .D(n36579), .CK(clk), .SN(1'b1), .RN(n37599),
        .QN(n34492) );
  DFFSRX1 data_queue_reg_7__5_ ( .D(n36578), .CK(clk), .SN(1'b1), .RN(n37599),
        .QN(n34493) );
  DFFSRX1 data_queue_reg_7__4_ ( .D(n36577), .CK(clk), .SN(1'b1), .RN(n37594),
        .QN(n34494) );
  DFFSRX1 data_queue_reg_7__3_ ( .D(n36576), .CK(clk), .SN(1'b1), .RN(n37601),
        .QN(n34495) );
  DFFSRX1 data_queue_reg_7__2_ ( .D(n36575), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n34496) );
  DFFSRX1 data_queue_reg_7__1_ ( .D(n36574), .CK(clk), .SN(1'b1), .RN(n37598),
        .QN(n34497) );
  DFFSRX1 dict_reg_35__4_ ( .D(n34809), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51260), .QN(n32684) );
  DFFSRX1 dict_reg_34__4_ ( .D(n34801), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51259), .QN(n32676) );
  DFFSRX1 dict_reg_67__4_ ( .D(n35065), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51292), .QN(n32940) );
  DFFSRX1 dict_reg_63__4_ ( .D(n35033), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51288), .QN(n32908) );
  DFFSRX1 dict_reg_66__4_ ( .D(n35057), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51291), .QN(n32932) );
  DFFSRX1 dict_reg_127__4_ ( .D(n35545), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51351), .QN(n33420) );
  DFFSRX1 dict_reg_130__4_ ( .D(n35569), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51354), .QN(n33444) );
  DFFSRX1 dict_reg_6__6_ ( .D(n34575), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50171), .QN(n32450) );
  DFFSRX1 dict_reg_142__6_ ( .D(n35663), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50307), .QN(n33538) );
  DFFSRX1 dict_reg_143__6_ ( .D(n35671), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50308), .QN(n33546) );
  DFFSRX1 dict_reg_168__6_ ( .D(n35871), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50333), .QN(n33746) );
  DFFSRX1 dict_reg_177__6_ ( .D(n35943), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50342), .QN(n33818) );
  DFFSRX1 dict_reg_194__6_ ( .D(n36079), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50359), .QN(n33954) );
  DFFSRX1 dict_reg_192__6_ ( .D(n36063), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50357), .QN(n33938) );
  DFFSRX1 dict_reg_82__6_ ( .D(n35183), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n50247), .QN(n33058) );
  DFFSRX1 dict_reg_33__4_ ( .D(n34793), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51258), .QN(n32668) );
  DFFSRX1 dict_reg_65__4_ ( .D(n35049), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51290), .QN(n32924) );
  DFFSRX1 dict_reg_128__4_ ( .D(n35553), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51352), .QN(n33428) );
  DFFSRX1 dict_reg_64__6_ ( .D(n35039), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50229), .QN(n32914) );
  DFFSRX1 dict_reg_131__4_ ( .D(n35577), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51355), .QN(n33452) );
  DFFSRX1 dict_reg_7__4_ ( .D(n34585), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51232), .QN(n32460) );
  DFFSRX1 dict_reg_162__4_ ( .D(n35825), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51386), .QN(n33700) );
  DFFSRX1 dict_reg_1__4_ ( .D(n34537), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51226), .QN(n32412) );
  DFFSRX1 dict_reg_15__4_ ( .D(n34649), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51240), .QN(n32524) );
  DFFSRX1 dict_reg_17__4_ ( .D(n34665), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51242), .QN(n32540) );
  DFFSRX1 dict_reg_9__4_ ( .D(n34601), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n51234), .QN(n32476) );
  DFFSRX1 dict_reg_213__6_ ( .D(n36231), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50378), .QN(n34106) );
  DFFSRX1 dict_reg_79__4_ ( .D(n35161), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51304), .QN(n33036) );
  DFFSRX1 dict_reg_134__4_ ( .D(n35601), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51358), .QN(n33476) );
  DFFSRX1 dict_reg_8__4_ ( .D(n34593), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51233), .QN(n32468) );
  DFFSRX1 dict_reg_208__4_ ( .D(n36193), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51432), .QN(n34068) );
  DFFSRX1 dict_reg_137__4_ ( .D(n35625), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51361), .QN(n33500) );
  DFFSRX1 dict_reg_57__6_ ( .D(n34983), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50222), .QN(n32858) );
  DFFRX2 dict_reg_155__2_ ( .D(n35771), .CK(clk), .RN(n42382), .Q(n50952),
        .QN(n33646) );
  DFFSRX1 dict_reg_1__6_ ( .D(n34535), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50166), .QN(n32410) );
  DFFSRX1 dict_reg_14__6_ ( .D(n34639), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50179), .QN(n32514) );
  DFFSRX1 dict_reg_21__6_ ( .D(n34695), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50186), .QN(n32570) );
  DFFSRX1 dict_reg_68__6_ ( .D(n35071), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n50233), .QN(n32946) );
  DFFSRX1 dict_reg_10__6_ ( .D(n34607), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50175), .QN(n32482) );
  DFFSRX1 dict_reg_46__6_ ( .D(n34895), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50211), .QN(n32770) );
  DFFSRX1 dict_reg_44__6_ ( .D(n34879), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50209), .QN(n32754) );
  DFFSRX1 dict_reg_23__6_ ( .D(n34711), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50188), .QN(n32586) );
  DFFSRX1 dict_reg_37__4_ ( .D(n34825), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51262), .QN(n32700) );
  DFFSRX1 dict_reg_49__4_ ( .D(n34921), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n51274), .QN(n32796) );
  DFFSRX1 dict_reg_47__4_ ( .D(n34905), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51272), .QN(n32780) );
  DFFSRX1 dict_reg_69__4_ ( .D(n35081), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51294), .QN(n32956) );
  DFFSRX1 dict_reg_73__6_ ( .D(n35111), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n50238), .QN(n32986) );
  DFFSRX1 dict_reg_67__6_ ( .D(n35063), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50232), .QN(n32938) );
  DFFSRX1 dict_reg_9__6_ ( .D(n34599), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50174), .QN(n32474) );
  DFFSRX1 dict_reg_2__6_ ( .D(n34543), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n50167), .QN(n32418) );
  DFFSRX1 dict_reg_151__6_ ( .D(n35735), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50316), .QN(n33610) );
  DFFSRX1 dict_reg_36__4_ ( .D(n34817), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51261), .QN(n32692) );
  DFFSRX1 dict_reg_68__4_ ( .D(n35073), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51293), .QN(n32948) );
  DFFSRX1 dict_reg_193__4_ ( .D(n36073), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51417), .QN(n33948) );
  DFFSRX1 dict_reg_161__4_ ( .D(n35817), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51385), .QN(n33692) );
  DFFSRX1 dict_reg_38__4_ ( .D(n34833), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51263), .QN(n32708) );
  DFFSRX1 dict_reg_138__4_ ( .D(n35633), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51362), .QN(n33508) );
  DFFSRX1 dict_reg_0__6_ ( .D(n34527), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50165), .QN(n32402) );
  DFFSRX1 dict_reg_56__6_ ( .D(n34975), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n50221), .QN(n32850) );
  DFFSRX1 dict_reg_72__6_ ( .D(n35103), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50237), .QN(n32978) );
  DFFSRX1 dict_reg_66__6_ ( .D(n35055), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n50231), .QN(n32930) );
  DFFSRX1 dict_reg_15__6_ ( .D(n34647), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50180), .QN(n32522) );
  DFFSRX1 dict_reg_8__6_ ( .D(n34591), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50173), .QN(n32466) );
  DFFSRX1 dict_reg_45__6_ ( .D(n34887), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50210), .QN(n32762) );
  DFFSRX1 dict_reg_22__6_ ( .D(n34703), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n50187), .QN(n32578) );
  DFFSRX1 dict_reg_199__6_ ( .D(n36119), .CK(clk), .SN(1'b1), .RN(n37595), .Q(
        n50364), .QN(n33994) );
  DFFSRX1 dict_reg_39__6_ ( .D(n34839), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n50204), .QN(n32714) );
  DFFSRX1 dict_reg_48__4_ ( .D(n34913), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51273), .QN(n32788) );
  DFFSRX1 dict_reg_16__4_ ( .D(n34657), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51241), .QN(n32532) );
  DFFSRX1 dict_reg_32__4_ ( .D(n34785), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51257), .QN(n32660) );
  DFFSRX1 dict_reg_70__4_ ( .D(n35089), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51295), .QN(n32964) );
  DFFSRX1 dict_reg_64__4_ ( .D(n35041), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51289), .QN(n32916) );
  DFFSRX1 dict_reg_135__4_ ( .D(n35609), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51359), .QN(n33484) );
  DFFSRX1 dict_reg_133__4_ ( .D(n35593), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51357), .QN(n33468) );
  DFFSRX1 dict_reg_129__4_ ( .D(n35561), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n51353), .QN(n33436) );
  DFFSRX1 dict_reg_197__4_ ( .D(n36105), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51421), .QN(n33980) );
  DFFSRX1 dict_reg_192__4_ ( .D(n36065), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n51416), .QN(n33940) );
  DFFSRX1 dict_reg_165__4_ ( .D(n35849), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n51389), .QN(n33724) );
  DFFSRX1 dict_reg_80__4_ ( .D(n35169), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51305), .QN(n33044) );
  DFFSRX1 dict_reg_136__4_ ( .D(n35617), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n51360), .QN(n33492) );
  DFFSRX1 dict_reg_176__4_ ( .D(n35937), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n51400), .QN(n33812) );
  DFFSRX1 dict_reg_175__4_ ( .D(n35929), .CK(clk), .SN(1'b1), .RN(n37591), .Q(
        n51399), .QN(n33804) );
  DFFSRX1 dict_reg_163__4_ ( .D(n35833), .CK(clk), .SN(1'b1), .RN(n37598), .Q(
        n51387), .QN(n33708) );
  DFFSRX1 dict_reg_160__4_ ( .D(n35809), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n51384), .QN(n33684) );
  DFFSRX1 dict_reg_0__4_ ( .D(n34529), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n51225), .QN(n32404) );
  DFFSRX1 dict_reg_214__6_ ( .D(n36239), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n50379), .QN(n34114) );
  DFFRX2 dict_reg_198__2_ ( .D(n36115), .CK(clk), .RN(n42385), .Q(n50995),
        .QN(n33990) );
  DFFRX2 dict_reg_180__2_ ( .D(n35971), .CK(clk), .RN(n42384), .Q(n50977),
        .QN(n33846) );
  DFFSRX1 dict_reg_214__7_ ( .D(n36238), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n49511), .QN(n34113) );
  DFFRX2 dict_reg_145__2_ ( .D(n35691), .CK(clk), .RN(n42381), .Q(n50942),
        .QN(n33566) );
  DFFRX2 dict_reg_212__3_ ( .D(n36226), .CK(clk), .RN(n42399), .Q(n51223),
        .QN(n34101) );
  DFFRX2 dict_reg_188__2_ ( .D(n36035), .CK(clk), .RN(n42384), .Q(n50985),
        .QN(n33910) );
  DFFRX2 dict_reg_127__7_ ( .D(n35542), .CK(clk), .RN(n42342), .Q(n50496),
        .QN(n33417) );
  DFFRX2 dict_reg_127__0_ ( .D(n35549), .CK(clk), .RN(n42355), .Q(n50710),
        .QN(n33424) );
  DFFRX2 dict_reg_127__2_ ( .D(n35547), .CK(clk), .RN(n42379), .Q(n50924),
        .QN(n33422) );
  DFFRX2 dict_reg_127__3_ ( .D(n35546), .CK(clk), .RN(n42392), .Q(n51138),
        .QN(n33421) );
  DFFRX2 dict_reg_211__3_ ( .D(n36218), .CK(clk), .RN(n42399), .Q(n51222),
        .QN(n34093) );
  DFFRX2 dict_reg_211__2_ ( .D(n36219), .CK(clk), .RN(n42386), .Q(n51008),
        .QN(n34094) );
  DFFRX2 dict_reg_148__0_ ( .D(n35717), .CK(clk), .RN(n42356), .Q(n50731),
        .QN(n33592) );
  DFFRX2 dict_reg_211__0_ ( .D(n36221), .CK(clk), .RN(n42362), .Q(n50794),
        .QN(n34096) );
  DFFRX2 dict_reg_148__3_ ( .D(n35714), .CK(clk), .RN(n42394), .Q(n51159),
        .QN(n33589) );
  DFFRX2 dict_reg_142__2_ ( .D(n35667), .CK(clk), .RN(n42381), .Q(n50939),
        .QN(n33542) );
  DFFRX2 dict_reg_196__7_ ( .D(n36094), .CK(clk), .RN(n42347), .Q(n50565),
        .QN(n33969) );
  DFFRX2 dict_reg_197__7_ ( .D(n36102), .CK(clk), .RN(n42347), .Q(n50566),
        .QN(n33977) );
  DFFRX2 dict_reg_141__0_ ( .D(n35661), .CK(clk), .RN(n42356), .Q(n50724),
        .QN(n33536) );
  DFFRX2 dict_reg_181__3_ ( .D(n35978), .CK(clk), .RN(n42396), .Q(n51192),
        .QN(n33853) );
  DFFRX2 dict_reg_212__0_ ( .D(n36229), .CK(clk), .RN(n42362), .Q(n50795),
        .QN(n34104) );
  DFFRX2 dict_reg_147__0_ ( .D(n35709), .CK(clk), .RN(n42356), .Q(n50730),
        .QN(n33584) );
  DFFRX2 dict_reg_149__0_ ( .D(n35725), .CK(clk), .RN(n42356), .Q(n50732),
        .QN(n33600) );
  DFFRX2 dict_reg_150__0_ ( .D(n35733), .CK(clk), .RN(n42356), .Q(n50733),
        .QN(n33608) );
  DFFRX2 dict_reg_187__0_ ( .D(n36029), .CK(clk), .RN(n42360), .Q(n50770),
        .QN(n33904) );
  DFFRX2 dict_reg_188__0_ ( .D(n36037), .CK(clk), .RN(n42360), .Q(n50771),
        .QN(n33912) );
  DFFRX2 dict_reg_147__2_ ( .D(n35707), .CK(clk), .RN(n42381), .Q(n50944),
        .QN(n33582) );
  DFFRX2 dict_reg_148__2_ ( .D(n35715), .CK(clk), .RN(n42381), .Q(n50945),
        .QN(n33590) );
  DFFRX2 dict_reg_187__2_ ( .D(n36027), .CK(clk), .RN(n42384), .Q(n50984),
        .QN(n33902) );
  DFFRX2 dict_reg_147__3_ ( .D(n35706), .CK(clk), .RN(n42393), .Q(n51158),
        .QN(n33581) );
  DFFRX2 dict_reg_188__3_ ( .D(n36034), .CK(clk), .RN(n42397), .Q(n51199),
        .QN(n33909) );
  DFFRX2 dict_reg_135__0_ ( .D(n35613), .CK(clk), .RN(n42355), .Q(n50718),
        .QN(n33488) );
  DFFSRX1 dict_reg_253__6_ ( .D(n36551), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n49336), .QN(n34426) );
  DFFRX2 dict_reg_122__0_ ( .D(n35509), .CK(clk), .RN(n42354), .Q(n50705),
        .QN(n33384) );
  DFFRX2 dict_reg_124__0_ ( .D(n35525), .CK(clk), .RN(n42354), .Q(n50707),
        .QN(n33400) );
  DFFRX2 dict_reg_126__0_ ( .D(n35541), .CK(clk), .RN(n42354), .Q(n50709),
        .QN(n33416) );
  DFFRX2 dict_reg_122__2_ ( .D(n35507), .CK(clk), .RN(n42379), .Q(n50919),
        .QN(n33382) );
  DFFRX2 dict_reg_124__2_ ( .D(n35523), .CK(clk), .RN(n42379), .Q(n50921),
        .QN(n33398) );
  DFFRX2 dict_reg_120__3_ ( .D(n35490), .CK(clk), .RN(n42391), .Q(n51131),
        .QN(n33365) );
  DFFRX2 dict_reg_124__3_ ( .D(n35522), .CK(clk), .RN(n42392), .Q(n51135),
        .QN(n33397) );
  DFFRX2 dict_reg_198__7_ ( .D(n36110), .CK(clk), .RN(n42347), .Q(n50567),
        .QN(n33985) );
  DFFRX2 dict_reg_128__0_ ( .D(n35557), .CK(clk), .RN(n42355), .Q(n50711),
        .QN(n33432) );
  DFFRX2 dict_reg_130__0_ ( .D(n35573), .CK(clk), .RN(n42355), .Q(n50713),
        .QN(n33448) );
  DFFRX2 dict_reg_131__0_ ( .D(n35581), .CK(clk), .RN(n42355), .Q(n50714),
        .QN(n33456) );
  DFFRX2 dict_reg_198__0_ ( .D(n36117), .CK(clk), .RN(n42360), .Q(n50781),
        .QN(n33992) );
  DFFRX2 dict_reg_199__0_ ( .D(n36125), .CK(clk), .RN(n42361), .Q(n50782),
        .QN(n34000) );
  DFFRX2 dict_reg_128__2_ ( .D(n35555), .CK(clk), .RN(n42379), .Q(n50925),
        .QN(n33430) );
  DFFRX2 dict_reg_130__2_ ( .D(n35571), .CK(clk), .RN(n42380), .Q(n50927),
        .QN(n33446) );
  DFFRX2 dict_reg_141__2_ ( .D(n35659), .CK(clk), .RN(n42381), .Q(n50938),
        .QN(n33534) );
  DFFRX2 dict_reg_199__2_ ( .D(n36123), .CK(clk), .RN(n42385), .Q(n50996),
        .QN(n33998) );
  DFFRX2 dict_reg_128__3_ ( .D(n35554), .CK(clk), .RN(n42392), .Q(n51139),
        .QN(n33429) );
  DFFRX2 dict_reg_130__3_ ( .D(n35570), .CK(clk), .RN(n42392), .Q(n51141),
        .QN(n33445) );
  DFFRX2 dict_reg_131__3_ ( .D(n35578), .CK(clk), .RN(n42392), .Q(n51142),
        .QN(n33453) );
  DFFRX2 dict_reg_141__3_ ( .D(n35658), .CK(clk), .RN(n42393), .Q(n51152),
        .QN(n33533) );
  DFFRX2 dict_reg_190__3_ ( .D(n36050), .CK(clk), .RN(n42397), .Q(n51201),
        .QN(n33925) );
  DFFRX2 dict_reg_198__3_ ( .D(n36114), .CK(clk), .RN(n42398), .Q(n51209),
        .QN(n33989) );
  DFFRX2 dict_reg_199__3_ ( .D(n36122), .CK(clk), .RN(n42398), .Q(n51210),
        .QN(n33997) );
  DFFRX2 dict_reg_134__0_ ( .D(n35605), .CK(clk), .RN(n42355), .Q(n50717),
        .QN(n33480) );
  DFFRX2 dict_reg_181__0_ ( .D(n35981), .CK(clk), .RN(n42359), .Q(n50764),
        .QN(n33856) );
  DFFRX2 dict_reg_181__2_ ( .D(n35979), .CK(clk), .RN(n42384), .Q(n50978),
        .QN(n33854) );
  DFFRX2 dict_reg_159__7_ ( .D(n35798), .CK(clk), .RN(n42345), .Q(n50528),
        .QN(n33673) );
  DFFRX2 dict_reg_163__7_ ( .D(n35830), .CK(clk), .RN(n42345), .Q(n50532),
        .QN(n33705) );
  DFFRX2 dict_reg_166__7_ ( .D(n35854), .CK(clk), .RN(n42345), .Q(n50535),
        .QN(n33729) );
  DFFRX2 dict_reg_177__7_ ( .D(n35942), .CK(clk), .RN(n42346), .Q(n50546),
        .QN(n33817) );
  DFFRX2 dict_reg_207__7_ ( .D(n36182), .CK(clk), .RN(n42348), .Q(n50576),
        .QN(n34057) );
  DFFRX2 dict_reg_208__7_ ( .D(n36190), .CK(clk), .RN(n42348), .Q(n50577),
        .QN(n34065) );
  DFFRX2 dict_reg_151__0_ ( .D(n35741), .CK(clk), .RN(n42357), .Q(n50734),
        .QN(n33616) );
  DFFRX2 dict_reg_156__0_ ( .D(n35781), .CK(clk), .RN(n42357), .Q(n50739),
        .QN(n33656) );
  DFFRX2 dict_reg_167__0_ ( .D(n35869), .CK(clk), .RN(n42358), .Q(n50750),
        .QN(n33744) );
  DFFRX2 dict_reg_177__0_ ( .D(n35949), .CK(clk), .RN(n42359), .Q(n50760),
        .QN(n33824) );
  DFFRX2 dict_reg_186__0_ ( .D(n36021), .CK(clk), .RN(n42359), .Q(n50769),
        .QN(n33896) );
  DFFRX2 dict_reg_201__0_ ( .D(n36141), .CK(clk), .RN(n42361), .Q(n50784),
        .QN(n34016) );
  DFFRX2 dict_reg_202__0_ ( .D(n36149), .CK(clk), .RN(n42361), .Q(n50785),
        .QN(n34024) );
  DFFRX2 dict_reg_204__0_ ( .D(n36165), .CK(clk), .RN(n42361), .Q(n50787),
        .QN(n34040) );
  DFFRX2 dict_reg_207__0_ ( .D(n36189), .CK(clk), .RN(n42361), .Q(n50790),
        .QN(n34064) );
  DFFRX2 dict_reg_210__0_ ( .D(n36213), .CK(clk), .RN(n42361), .Q(n50793),
        .QN(n34088) );
  DFFRX2 dict_reg_143__2_ ( .D(n35675), .CK(clk), .RN(n42381), .Q(n50940),
        .QN(n33550) );
  DFFRX2 dict_reg_149__2_ ( .D(n35723), .CK(clk), .RN(n42381), .Q(n50946),
        .QN(n33598) );
  DFFRX2 dict_reg_150__2_ ( .D(n35731), .CK(clk), .RN(n42381), .Q(n50947),
        .QN(n33606) );
  DFFRX2 dict_reg_156__2_ ( .D(n35779), .CK(clk), .RN(n42382), .Q(n50953),
        .QN(n33654) );
  DFFRX2 dict_reg_157__2_ ( .D(n35787), .CK(clk), .RN(n42382), .Q(n50954),
        .QN(n33662) );
  DFFRX2 dict_reg_167__2_ ( .D(n35867), .CK(clk), .RN(n42383), .Q(n50964),
        .QN(n33742) );
  DFFRX2 dict_reg_175__2_ ( .D(n35931), .CK(clk), .RN(n42383), .Q(n50972),
        .QN(n33806) );
  DFFRX2 dict_reg_177__2_ ( .D(n35947), .CK(clk), .RN(n42384), .Q(n50974),
        .QN(n33822) );
  DFFRX2 dict_reg_178__2_ ( .D(n35955), .CK(clk), .RN(n42384), .Q(n50975),
        .QN(n33830) );
  DFFRX2 dict_reg_191__2_ ( .D(n36059), .CK(clk), .RN(n42385), .Q(n50988),
        .QN(n33934) );
  DFFRX2 dict_reg_201__2_ ( .D(n36139), .CK(clk), .RN(n42386), .Q(n50998),
        .QN(n34014) );
  DFFRX2 dict_reg_207__2_ ( .D(n36187), .CK(clk), .RN(n42386), .Q(n51004),
        .QN(n34062) );
  DFFRX2 dict_reg_143__3_ ( .D(n35674), .CK(clk), .RN(n42393), .Q(n51154),
        .QN(n33549) );
  DFFRX2 dict_reg_144__3_ ( .D(n35682), .CK(clk), .RN(n42393), .Q(n51155),
        .QN(n33557) );
  DFFRX2 dict_reg_149__3_ ( .D(n35722), .CK(clk), .RN(n42394), .Q(n51160),
        .QN(n33597) );
  DFFRX2 dict_reg_151__3_ ( .D(n35738), .CK(clk), .RN(n42394), .Q(n51162),
        .QN(n33613) );
  DFFRX2 dict_reg_156__3_ ( .D(n35778), .CK(clk), .RN(n42394), .Q(n51167),
        .QN(n33653) );
  DFFRX2 dict_reg_167__3_ ( .D(n35866), .CK(clk), .RN(n42395), .Q(n51178),
        .QN(n33741) );
  DFFRX2 dict_reg_169__3_ ( .D(n35882), .CK(clk), .RN(n42395), .Q(n51180),
        .QN(n33757) );
  DFFRX2 dict_reg_176__3_ ( .D(n35938), .CK(clk), .RN(n42396), .Q(n51187),
        .QN(n33813) );
  DFFRX2 dict_reg_177__3_ ( .D(n35946), .CK(clk), .RN(n42396), .Q(n51188),
        .QN(n33821) );
  DFFRX2 dict_reg_179__3_ ( .D(n35962), .CK(clk), .RN(n42396), .Q(n51190),
        .QN(n33837) );
  DFFRX2 dict_reg_187__3_ ( .D(n36026), .CK(clk), .RN(n42397), .Q(n51198),
        .QN(n33901) );
  DFFRX2 dict_reg_201__3_ ( .D(n36138), .CK(clk), .RN(n42398), .Q(n51212),
        .QN(n34013) );
  DFFRX2 dict_reg_202__3_ ( .D(n36146), .CK(clk), .RN(n42398), .Q(n51213),
        .QN(n34021) );
  DFFRX2 dict_reg_205__3_ ( .D(n36170), .CK(clk), .RN(n42398), .Q(n51216),
        .QN(n34045) );
  DFFRX2 dict_reg_207__3_ ( .D(n36186), .CK(clk), .RN(n42398), .Q(n51218),
        .QN(n34061) );
  DFFRX2 dict_reg_210__3_ ( .D(n36210), .CK(clk), .RN(n42399), .Q(n51221),
        .QN(n34085) );
  DFFRX2 dict_reg_210__2_ ( .D(n36211), .CK(clk), .RN(n42386), .Q(n51007),
        .QN(n34086) );
  DFFRX2 dict_reg_212__2_ ( .D(n36227), .CK(clk), .RN(n42386), .Q(n51009),
        .QN(n34102) );
  DFFSRX1 dict_reg_253__0_ ( .D(n36557), .CK(clk), .SN(1'b1), .RN(n37593), .Q(
        n49025), .QN(n34432) );
  DFFSRX1 data_num_reg_1_ ( .D(nxt_data_num[1]), .CK(clk), .SN(1'b1), .RN(
        n37595), .Q(n50134), .QN(n32399) );
  DFFSRX1 dict_reg_253__2_ ( .D(n36555), .CK(clk), .SN(1'b1), .RN(n37592), .Q(
        n48874), .QN(n34430) );
  DFFRX2 dict_reg_93__0_ ( .D(n35277), .CK(clk), .RN(n42352), .Q(n50676), .QN(
        n33152) );
  DFFRX2 dict_reg_93__2_ ( .D(n35275), .CK(clk), .RN(n42377), .Q(n50890), .QN(
        n33150) );
  DFFRX2 dict_reg_93__3_ ( .D(n35274), .CK(clk), .RN(n42390), .Q(n51104), .QN(
        n33149) );
  DFFRX2 dict_reg_94__0_ ( .D(n35285), .CK(clk), .RN(n42352), .Q(n50677), .QN(
        n33160) );
  DFFRX2 dict_reg_94__2_ ( .D(n35283), .CK(clk), .RN(n42377), .Q(n50891), .QN(
        n33158) );
  DFFRX2 dict_reg_94__3_ ( .D(n35282), .CK(clk), .RN(n42390), .Q(n51105), .QN(
        n33157) );
  DFFRX2 dict_reg_111__3_ ( .D(n35418), .CK(clk), .RN(n37594), .Q(n51122),
        .QN(n33293) );
  DFFRX2 dict_reg_112__7_ ( .D(n35422), .CK(clk), .RN(n42341), .Q(n50483),
        .QN(n33297) );
  DFFRX2 dict_reg_113__7_ ( .D(n35430), .CK(clk), .RN(n42341), .Q(n50484),
        .QN(n33305) );
  DFFRX2 dict_reg_112__0_ ( .D(n35429), .CK(clk), .RN(n42353), .Q(n50695),
        .QN(n33304) );
  DFFRX2 dict_reg_113__0_ ( .D(n35437), .CK(clk), .RN(n42353), .Q(n50696),
        .QN(n33312) );
  DFFRX2 dict_reg_114__0_ ( .D(n35445), .CK(clk), .RN(n42353), .Q(n50697),
        .QN(n33320) );
  DFFRX2 dict_reg_115__0_ ( .D(n35453), .CK(clk), .RN(n42354), .Q(n50698),
        .QN(n33328) );
  DFFRX2 dict_reg_116__0_ ( .D(n35461), .CK(clk), .RN(n42354), .Q(n50699),
        .QN(n33336) );
  DFFRX2 dict_reg_117__0_ ( .D(n35469), .CK(clk), .RN(n42354), .Q(n50700),
        .QN(n33344) );
  DFFRX2 dict_reg_118__0_ ( .D(n35477), .CK(clk), .RN(n42354), .Q(n50701),
        .QN(n33352) );
  DFFRX2 dict_reg_120__0_ ( .D(n35493), .CK(clk), .RN(n42354), .Q(n50703),
        .QN(n33368) );
  DFFRX2 dict_reg_121__0_ ( .D(n35501), .CK(clk), .RN(n42354), .Q(n50704),
        .QN(n33376) );
  DFFRX2 dict_reg_112__2_ ( .D(n35427), .CK(clk), .RN(n42378), .Q(n50909),
        .QN(n33302) );
  DFFRX2 dict_reg_113__2_ ( .D(n35435), .CK(clk), .RN(n42378), .Q(n50910),
        .QN(n33310) );
  DFFRX2 dict_reg_114__2_ ( .D(n35443), .CK(clk), .RN(n42378), .Q(n50911),
        .QN(n33318) );
  DFFRX2 dict_reg_115__2_ ( .D(n35451), .CK(clk), .RN(n42378), .Q(n50912),
        .QN(n33326) );
  DFFRX2 dict_reg_116__2_ ( .D(n35459), .CK(clk), .RN(n42378), .Q(n50913),
        .QN(n33334) );
  DFFRX2 dict_reg_117__2_ ( .D(n35467), .CK(clk), .RN(n42379), .Q(n50914),
        .QN(n33342) );
  DFFRX2 dict_reg_118__2_ ( .D(n35475), .CK(clk), .RN(n42379), .Q(n50915),
        .QN(n33350) );
  DFFRX2 dict_reg_120__2_ ( .D(n35491), .CK(clk), .RN(n42379), .Q(n50917),
        .QN(n33366) );
  DFFRX2 dict_reg_121__2_ ( .D(n35499), .CK(clk), .RN(n42379), .Q(n50918),
        .QN(n33374) );
  DFFRX2 dict_reg_112__3_ ( .D(n35426), .CK(clk), .RN(n42391), .Q(n51123),
        .QN(n33301) );
  DFFRX2 dict_reg_113__3_ ( .D(n35434), .CK(clk), .RN(n42391), .Q(n51124),
        .QN(n33309) );
  DFFRX2 dict_reg_114__3_ ( .D(n35442), .CK(clk), .RN(n42391), .Q(n51125),
        .QN(n33317) );
  DFFRX2 dict_reg_115__3_ ( .D(n35450), .CK(clk), .RN(n42391), .Q(n51126),
        .QN(n33325) );
  DFFRX2 dict_reg_116__3_ ( .D(n35458), .CK(clk), .RN(n42391), .Q(n51127),
        .QN(n33333) );
  DFFRX2 dict_reg_117__3_ ( .D(n35466), .CK(clk), .RN(n42391), .Q(n51128),
        .QN(n33341) );
  DFFRX2 dict_reg_118__3_ ( .D(n35474), .CK(clk), .RN(n42391), .Q(n51129),
        .QN(n33349) );
  DFFRX2 dict_reg_121__3_ ( .D(n35498), .CK(clk), .RN(n42391), .Q(n51132),
        .QN(n33373) );
  DFFRX2 dict_reg_122__3_ ( .D(n35506), .CK(clk), .RN(n42391), .Q(n51133),
        .QN(n33381) );
  DFFRX2 dict_reg_128__7_ ( .D(n35550), .CK(clk), .RN(n42342), .Q(n50497),
        .QN(n33425) );
  DFFRX2 dict_reg_131__7_ ( .D(n35574), .CK(clk), .RN(n42342), .Q(n50500),
        .QN(n33449) );
  DFFRX2 dict_reg_161__7_ ( .D(n35814), .CK(clk), .RN(n42345), .Q(n50530),
        .QN(n33689) );
  DFFRX2 dict_reg_191__7_ ( .D(n36054), .CK(clk), .RN(n37596), .Q(n50560),
        .QN(n33929) );
  DFFRX2 dict_reg_194__7_ ( .D(n36078), .CK(clk), .RN(n42347), .Q(n50563),
        .QN(n33953) );
  DFFRX2 dict_reg_195__7_ ( .D(n36086), .CK(clk), .RN(n42347), .Q(n50564),
        .QN(n33961) );
  DFFRX2 dict_reg_123__0_ ( .D(n35517), .CK(clk), .RN(n42354), .Q(n50706),
        .QN(n33392) );
  DFFRX2 dict_reg_139__0_ ( .D(n35645), .CK(clk), .RN(n42356), .Q(n50722),
        .QN(n33520) );
  DFFRX2 dict_reg_152__0_ ( .D(n35749), .CK(clk), .RN(n42357), .Q(n50735),
        .QN(n33624) );
  DFFRX2 dict_reg_191__0_ ( .D(n36061), .CK(clk), .RN(n42360), .Q(n50774),
        .QN(n33936) );
  DFFRX2 dict_reg_195__0_ ( .D(n36093), .CK(clk), .RN(n42360), .Q(n50778),
        .QN(n33968) );
  DFFRX2 dict_reg_197__0_ ( .D(n36109), .CK(clk), .RN(n42360), .Q(n50780),
        .QN(n33984) );
  DFFRX2 dict_reg_200__0_ ( .D(n36133), .CK(clk), .RN(n42361), .Q(n50783),
        .QN(n34008) );
  DFFRX2 dict_reg_123__2_ ( .D(n35515), .CK(clk), .RN(n42379), .Q(n50920),
        .QN(n33390) );
  DFFRX2 dict_reg_129__2_ ( .D(n35563), .CK(clk), .RN(n42380), .Q(n50926),
        .QN(n33438) );
  DFFRX2 dict_reg_131__2_ ( .D(n35579), .CK(clk), .RN(n42380), .Q(n50928),
        .QN(n33454) );
  DFFRX2 dict_reg_139__2_ ( .D(n35643), .CK(clk), .RN(n42380), .Q(n50936),
        .QN(n33518) );
  DFFRX2 dict_reg_152__2_ ( .D(n35747), .CK(clk), .RN(n42381), .Q(n50949),
        .QN(n33622) );
  DFFRX2 dict_reg_165__2_ ( .D(n35851), .CK(clk), .RN(n42383), .Q(n50962),
        .QN(n33726) );
  DFFRX2 dict_reg_172__2_ ( .D(n35907), .CK(clk), .RN(n42383), .Q(n50969),
        .QN(n33782) );
  DFFRX2 dict_reg_182__2_ ( .D(n35987), .CK(clk), .RN(n42384), .Q(n50979),
        .QN(n33862) );
  DFFRX2 dict_reg_190__2_ ( .D(n36051), .CK(clk), .RN(n42385), .Q(n50987),
        .QN(n33926) );
  DFFRX2 dict_reg_195__2_ ( .D(n36091), .CK(clk), .RN(n42385), .Q(n50992),
        .QN(n33966) );
  DFFRX2 dict_reg_196__2_ ( .D(n36099), .CK(clk), .RN(n42385), .Q(n50993),
        .QN(n33974) );
  DFFRX2 dict_reg_197__2_ ( .D(n36107), .CK(clk), .RN(n42385), .Q(n50994),
        .QN(n33982) );
  DFFRX2 dict_reg_200__2_ ( .D(n36131), .CK(clk), .RN(n42385), .Q(n50997),
        .QN(n34006) );
  DFFRX2 dict_reg_123__3_ ( .D(n35514), .CK(clk), .RN(n42391), .Q(n51134),
        .QN(n33389) );
  DFFRX2 dict_reg_129__3_ ( .D(n35562), .CK(clk), .RN(n42392), .Q(n51140),
        .QN(n33437) );
  DFFRX2 dict_reg_139__3_ ( .D(n35642), .CK(clk), .RN(n42393), .Q(n51150),
        .QN(n33517) );
  DFFRX2 dict_reg_152__3_ ( .D(n35746), .CK(clk), .RN(n42394), .Q(n51163),
        .QN(n33621) );
  DFFRX2 dict_reg_182__3_ ( .D(n35986), .CK(clk), .RN(n42396), .Q(n51193),
        .QN(n33861) );
  DFFRX2 dict_reg_195__3_ ( .D(n36090), .CK(clk), .RN(n42397), .Q(n51206),
        .QN(n33965) );
  DFFRX2 dict_reg_196__3_ ( .D(n36098), .CK(clk), .RN(n42398), .Q(n51207),
        .QN(n33973) );
  DFFRX2 dict_reg_197__3_ ( .D(n36106), .CK(clk), .RN(n42398), .Q(n51208),
        .QN(n33981) );
  DFFRX2 dict_reg_200__3_ ( .D(n36130), .CK(clk), .RN(n42398), .Q(n51211),
        .QN(n34005) );
  DFFRX2 dict_reg_137__7_ ( .D(n35622), .CK(clk), .RN(n42343), .Q(n50506),
        .QN(n33497) );
  DFFRX2 dict_reg_132__0_ ( .D(n35589), .CK(clk), .RN(n42355), .Q(n50715),
        .QN(n33464) );
  DFFRX2 dict_reg_136__0_ ( .D(n35621), .CK(clk), .RN(n42355), .Q(n50719),
        .QN(n33496) );
  DFFRX2 dict_reg_132__2_ ( .D(n35587), .CK(clk), .RN(n42380), .Q(n50929),
        .QN(n33462) );
  DFFRX2 dict_reg_134__2_ ( .D(n35603), .CK(clk), .RN(n42380), .Q(n50931),
        .QN(n33478) );
  DFFRX2 dict_reg_136__2_ ( .D(n35619), .CK(clk), .RN(n42380), .Q(n50933),
        .QN(n33494) );
  DFFRX2 dict_reg_137__2_ ( .D(n35627), .CK(clk), .RN(n42380), .Q(n50934),
        .QN(n33502) );
  DFFRX2 dict_reg_132__3_ ( .D(n35586), .CK(clk), .RN(n42392), .Q(n51143),
        .QN(n33461) );
  DFFRX2 dict_reg_134__3_ ( .D(n35602), .CK(clk), .RN(n42392), .Q(n51145),
        .QN(n33477) );
  DFFRX2 dict_reg_136__3_ ( .D(n35618), .CK(clk), .RN(n42393), .Q(n51147),
        .QN(n33493) );
  DFFRX2 dict_reg_137__3_ ( .D(n35626), .CK(clk), .RN(n42393), .Q(n51148),
        .QN(n33501) );
  DFFRX2 dict_reg_144__7_ ( .D(n35678), .CK(clk), .RN(n42344), .Q(n50513),
        .QN(n33553) );
  DFFRX2 dict_reg_160__7_ ( .D(n35806), .CK(clk), .RN(n42345), .Q(n50529),
        .QN(n33681) );
  DFFRX2 dict_reg_162__7_ ( .D(n35822), .CK(clk), .RN(n42345), .Q(n50531),
        .QN(n33697) );
  DFFRX2 dict_reg_164__7_ ( .D(n35838), .CK(clk), .RN(n42345), .Q(n50533),
        .QN(n33713) );
  DFFRX2 dict_reg_175__7_ ( .D(n35926), .CK(clk), .RN(n42346), .Q(n50544),
        .QN(n33801) );
  DFFRX2 dict_reg_176__7_ ( .D(n35934), .CK(clk), .RN(n42346), .Q(n50545),
        .QN(n33809) );
  DFFRX2 dict_reg_142__0_ ( .D(n35669), .CK(clk), .RN(n42356), .Q(n50725),
        .QN(n33544) );
  DFFRX2 dict_reg_143__0_ ( .D(n35677), .CK(clk), .RN(n42356), .Q(n50726),
        .QN(n33552) );
  DFFRX2 dict_reg_144__0_ ( .D(n35685), .CK(clk), .RN(n42356), .Q(n50727),
        .QN(n33560) );
  DFFRX2 dict_reg_145__0_ ( .D(n35693), .CK(clk), .RN(n42356), .Q(n50728),
        .QN(n33568) );
  DFFRX2 dict_reg_146__0_ ( .D(n35701), .CK(clk), .RN(n42356), .Q(n50729),
        .QN(n33576) );
  DFFRX2 dict_reg_157__0_ ( .D(n35789), .CK(clk), .RN(n42357), .Q(n50740),
        .QN(n33664) );
  DFFRX2 dict_reg_163__0_ ( .D(n35837), .CK(clk), .RN(n42358), .Q(n50746),
        .QN(n33712) );
  DFFRX2 dict_reg_164__0_ ( .D(n35845), .CK(clk), .RN(n42358), .Q(n50747),
        .QN(n33720) );
  DFFRX2 dict_reg_165__0_ ( .D(n35853), .CK(clk), .RN(n42358), .Q(n50748),
        .QN(n33728) );
  DFFRX2 dict_reg_166__0_ ( .D(n35861), .CK(clk), .RN(n42358), .Q(n50749),
        .QN(n33736) );
  DFFRX2 dict_reg_169__0_ ( .D(n35885), .CK(clk), .RN(n42358), .Q(n50752),
        .QN(n33760) );
  DFFRX2 dict_reg_170__0_ ( .D(n35893), .CK(clk), .RN(n42358), .Q(n50753),
        .QN(n33768) );
  DFFRX2 dict_reg_176__0_ ( .D(n35941), .CK(clk), .RN(n42359), .Q(n50759),
        .QN(n33816) );
  DFFRX2 dict_reg_178__0_ ( .D(n35957), .CK(clk), .RN(n42359), .Q(n50761),
        .QN(n33832) );
  DFFRX2 dict_reg_179__0_ ( .D(n35965), .CK(clk), .RN(n42359), .Q(n50762),
        .QN(n33840) );
  DFFRX2 dict_reg_184__0_ ( .D(n36005), .CK(clk), .RN(n42359), .Q(n50767),
        .QN(n33880) );
  DFFRX2 dict_reg_185__0_ ( .D(n36013), .CK(clk), .RN(n42359), .Q(n50768),
        .QN(n33888) );
  DFFRX2 dict_reg_190__0_ ( .D(n36053), .CK(clk), .RN(n42360), .Q(n50773),
        .QN(n33928) );
  DFFRX2 dict_reg_192__0_ ( .D(n36069), .CK(clk), .RN(n42360), .Q(n50775),
        .QN(n33944) );
  DFFRX2 dict_reg_193__0_ ( .D(n36077), .CK(clk), .RN(n42360), .Q(n50776),
        .QN(n33952) );
  DFFRX2 dict_reg_203__0_ ( .D(n36157), .CK(clk), .RN(n42361), .Q(n50786),
        .QN(n34032) );
  DFFRX2 dict_reg_205__0_ ( .D(n36173), .CK(clk), .RN(n42361), .Q(n50788),
        .QN(n34048) );
  DFFRX2 dict_reg_206__0_ ( .D(n36181), .CK(clk), .RN(n42361), .Q(n50789),
        .QN(n34056) );
  DFFRX2 dict_reg_144__2_ ( .D(n35683), .CK(clk), .RN(n42381), .Q(n50941),
        .QN(n33558) );
  DFFRX2 dict_reg_151__2_ ( .D(n35739), .CK(clk), .RN(n42381), .Q(n50948),
        .QN(n33614) );
  DFFRX2 dict_reg_153__2_ ( .D(n35755), .CK(clk), .RN(n42382), .Q(n50950),
        .QN(n33630) );
  DFFRX2 dict_reg_163__2_ ( .D(n35835), .CK(clk), .RN(n42382), .Q(n50960),
        .QN(n33710) );
  DFFRX2 dict_reg_164__2_ ( .D(n35843), .CK(clk), .RN(n42382), .Q(n50961),
        .QN(n33718) );
  DFFRX2 dict_reg_169__2_ ( .D(n35883), .CK(clk), .RN(n42383), .Q(n50966),
        .QN(n33758) );
  DFFRX2 dict_reg_170__2_ ( .D(n35891), .CK(clk), .RN(n42383), .Q(n50967),
        .QN(n33766) );
  DFFRX2 dict_reg_176__2_ ( .D(n35939), .CK(clk), .RN(n42383), .Q(n50973),
        .QN(n33814) );
  DFFRX2 dict_reg_186__2_ ( .D(n36019), .CK(clk), .RN(n42384), .Q(n50983),
        .QN(n33894) );
  DFFRX2 dict_reg_189__2_ ( .D(n36043), .CK(clk), .RN(n42385), .Q(n50986),
        .QN(n33918) );
  DFFRX2 dict_reg_192__2_ ( .D(n36067), .CK(clk), .RN(n42385), .Q(n50989),
        .QN(n33942) );
  DFFRX2 dict_reg_193__2_ ( .D(n36075), .CK(clk), .RN(n42385), .Q(n50990),
        .QN(n33950) );
  DFFRX2 dict_reg_202__2_ ( .D(n36147), .CK(clk), .RN(n42386), .Q(n50999),
        .QN(n34022) );
  DFFRX2 dict_reg_206__2_ ( .D(n36179), .CK(clk), .RN(n42386), .Q(n51003),
        .QN(n34054) );
  DFFRX2 dict_reg_209__2_ ( .D(n36203), .CK(clk), .RN(n42386), .Q(n51006),
        .QN(n34078) );
  DFFRX2 dict_reg_142__3_ ( .D(n35666), .CK(clk), .RN(n42393), .Q(n51153),
        .QN(n33541) );
  DFFRX2 dict_reg_146__3_ ( .D(n35698), .CK(clk), .RN(n42393), .Q(n51157),
        .QN(n33573) );
  DFFRX2 dict_reg_150__3_ ( .D(n35730), .CK(clk), .RN(n42394), .Q(n51161),
        .QN(n33605) );
  DFFRX2 dict_reg_157__3_ ( .D(n35786), .CK(clk), .RN(n42394), .Q(n51168),
        .QN(n33661) );
  DFFRX2 dict_reg_163__3_ ( .D(n35834), .CK(clk), .RN(n42395), .Q(n51174),
        .QN(n33709) );
  DFFRX2 dict_reg_164__3_ ( .D(n35842), .CK(clk), .RN(n42395), .Q(n51175),
        .QN(n33717) );
  DFFRX2 dict_reg_165__3_ ( .D(n35850), .CK(clk), .RN(n42395), .Q(n51176),
        .QN(n33725) );
  DFFRX2 dict_reg_166__3_ ( .D(n35858), .CK(clk), .RN(n42395), .Q(n51177),
        .QN(n33733) );
  DFFRX2 dict_reg_170__3_ ( .D(n35890), .CK(clk), .RN(n42395), .Q(n51181),
        .QN(n33765) );
  DFFRX2 dict_reg_175__3_ ( .D(n35930), .CK(clk), .RN(n42396), .Q(n51186),
        .QN(n33805) );
  DFFRX2 dict_reg_178__3_ ( .D(n35954), .CK(clk), .RN(n42396), .Q(n51189),
        .QN(n33829) );
  DFFRX2 dict_reg_184__3_ ( .D(n36002), .CK(clk), .RN(n42397), .Q(n51195),
        .QN(n33877) );
  DFFRX2 dict_reg_186__3_ ( .D(n36018), .CK(clk), .RN(n42397), .Q(n51197),
        .QN(n33893) );
  DFFRX2 dict_reg_192__3_ ( .D(n36066), .CK(clk), .RN(n42397), .Q(n51203),
        .QN(n33941) );
  DFFRX2 dict_reg_193__3_ ( .D(n36074), .CK(clk), .RN(n42397), .Q(n51204),
        .QN(n33949) );
  DFFRX2 dict_reg_203__3_ ( .D(n36154), .CK(clk), .RN(n42398), .Q(n51214),
        .QN(n34029) );
  DFFRX2 dict_reg_204__3_ ( .D(n36162), .CK(clk), .RN(n42398), .Q(n51215),
        .QN(n34037) );
  DFFRX2 dict_reg_206__3_ ( .D(n36178), .CK(clk), .RN(n42398), .Q(n51217),
        .QN(n34053) );
  DFFRX2 dict_reg_143__7_ ( .D(n35670), .CK(clk), .RN(n42343), .Q(n50512),
        .QN(n33545) );
  DFFSRX1 dict_reg_253__3_ ( .D(n36554), .CK(clk), .SN(1'b1), .RN(n37590), .Q(
        n48716), .QN(n34429) );
  DFFRX2 dict_reg_213__0_ ( .D(n36237), .CK(clk), .RN(n42362), .Q(n50796),
        .QN(n34112) );
  DFFRX2 dict_reg_213__3_ ( .D(n36234), .CK(clk), .RN(n42399), .Q(n51224),
        .QN(n34109) );
  DFFRX2 dict_reg_77__0_ ( .D(n35149), .CK(clk), .RN(n42350), .Q(n50660), .QN(
        n33024) );
  DFFRX2 dict_reg_78__0_ ( .D(n35157), .CK(clk), .RN(n42350), .Q(n50661), .QN(
        n33032) );
  DFFRX2 dict_reg_77__2_ ( .D(n35147), .CK(clk), .RN(n42375), .Q(n50874), .QN(
        n33022) );
  DFFRX2 dict_reg_78__2_ ( .D(n35155), .CK(clk), .RN(n42375), .Q(n50875), .QN(
        n33030) );
  DFFRX2 dict_reg_77__3_ ( .D(n35146), .CK(clk), .RN(n42389), .Q(n51088), .QN(
        n33021) );
  DFFRX2 dict_reg_78__3_ ( .D(n35154), .CK(clk), .RN(n42389), .Q(n51089), .QN(
        n33029) );
  DFFRX2 dict_reg_79__7_ ( .D(n35158), .CK(clk), .RN(n42339), .Q(n50453), .QN(
        n33033) );
  DFFRX2 dict_reg_80__7_ ( .D(n35166), .CK(clk), .RN(n42339), .Q(n50454), .QN(
        n33041) );
  DFFRX2 dict_reg_79__0_ ( .D(n35165), .CK(clk), .RN(n42351), .Q(n50662), .QN(
        n33040) );
  DFFRX2 dict_reg_80__0_ ( .D(n35173), .CK(clk), .RN(n42351), .Q(n50663), .QN(
        n33048) );
  DFFRX2 dict_reg_81__0_ ( .D(n35181), .CK(clk), .RN(n42351), .Q(n50664), .QN(
        n33056) );
  DFFRX2 dict_reg_82__0_ ( .D(n35189), .CK(clk), .RN(n42351), .Q(n50665), .QN(
        n33064) );
  DFFRX2 dict_reg_83__0_ ( .D(n35197), .CK(clk), .RN(n42351), .Q(n50666), .QN(
        n33072) );
  DFFRX2 dict_reg_84__0_ ( .D(n35205), .CK(clk), .RN(n42351), .Q(n50667), .QN(
        n33080) );
  DFFRX2 dict_reg_85__0_ ( .D(n35213), .CK(clk), .RN(n42351), .Q(n50668), .QN(
        n33088) );
  DFFRX2 dict_reg_86__0_ ( .D(n35221), .CK(clk), .RN(n42351), .Q(n50669), .QN(
        n33096) );
  DFFRX2 dict_reg_87__0_ ( .D(n35229), .CK(clk), .RN(n42351), .Q(n50670), .QN(
        n33104) );
  DFFRX2 dict_reg_88__0_ ( .D(n35237), .CK(clk), .RN(n42351), .Q(n50671), .QN(
        n33112) );
  DFFRX2 dict_reg_89__0_ ( .D(n35245), .CK(clk), .RN(n42351), .Q(n50672), .QN(
        n33120) );
  DFFRX2 dict_reg_79__2_ ( .D(n35163), .CK(clk), .RN(n42375), .Q(n50876), .QN(
        n33038) );
  DFFRX2 dict_reg_80__2_ ( .D(n35171), .CK(clk), .RN(n42375), .Q(n50877), .QN(
        n33046) );
  DFFRX2 dict_reg_81__2_ ( .D(n35179), .CK(clk), .RN(n42376), .Q(n50878), .QN(
        n33054) );
  DFFRX2 dict_reg_82__2_ ( .D(n35187), .CK(clk), .RN(n42376), .Q(n50879), .QN(
        n33062) );
  DFFRX2 dict_reg_83__2_ ( .D(n35195), .CK(clk), .RN(n42376), .Q(n50880), .QN(
        n33070) );
  DFFRX2 dict_reg_84__2_ ( .D(n35203), .CK(clk), .RN(n42376), .Q(n50881), .QN(
        n33078) );
  DFFRX2 dict_reg_85__2_ ( .D(n35211), .CK(clk), .RN(n42376), .Q(n50882), .QN(
        n33086) );
  DFFRX2 dict_reg_86__2_ ( .D(n35219), .CK(clk), .RN(n42376), .Q(n50883), .QN(
        n33094) );
  DFFRX2 dict_reg_87__2_ ( .D(n35227), .CK(clk), .RN(n42376), .Q(n50884), .QN(
        n33102) );
  DFFRX2 dict_reg_88__2_ ( .D(n35235), .CK(clk), .RN(n42376), .Q(n50885), .QN(
        n33110) );
  DFFRX2 dict_reg_89__2_ ( .D(n35243), .CK(clk), .RN(n42376), .Q(n50886), .QN(
        n33118) );
  DFFRX2 dict_reg_90__2_ ( .D(n35251), .CK(clk), .RN(n42376), .Q(n50887), .QN(
        n33126) );
  DFFRX2 dict_reg_79__3_ ( .D(n35162), .CK(clk), .RN(n42389), .Q(n51090), .QN(
        n33037) );
  DFFRX2 dict_reg_80__3_ ( .D(n35170), .CK(clk), .RN(n42389), .Q(n51091), .QN(
        n33045) );
  DFFRX2 dict_reg_81__3_ ( .D(n35178), .CK(clk), .RN(n42389), .Q(n51092), .QN(
        n33053) );
  DFFRX2 dict_reg_82__3_ ( .D(n35186), .CK(clk), .RN(n42389), .Q(n51093), .QN(
        n33061) );
  DFFRX2 dict_reg_83__3_ ( .D(n35194), .CK(clk), .RN(n42389), .Q(n51094), .QN(
        n33069) );
  DFFRX2 dict_reg_84__3_ ( .D(n35202), .CK(clk), .RN(n42389), .Q(n51095), .QN(
        n33077) );
  DFFRX2 dict_reg_85__3_ ( .D(n35210), .CK(clk), .RN(n42389), .Q(n51096), .QN(
        n33085) );
  DFFRX2 dict_reg_86__3_ ( .D(n35218), .CK(clk), .RN(n42389), .Q(n51097), .QN(
        n33093) );
  DFFRX2 dict_reg_87__3_ ( .D(n35226), .CK(clk), .RN(n42389), .Q(n51098), .QN(
        n33101) );
  DFFRX2 dict_reg_88__3_ ( .D(n35234), .CK(clk), .RN(n42390), .Q(n51099), .QN(
        n33109) );
  DFFRX2 dict_reg_89__3_ ( .D(n35242), .CK(clk), .RN(n42390), .Q(n51100), .QN(
        n33117) );
  DFFRX2 dict_reg_90__3_ ( .D(n35250), .CK(clk), .RN(n42390), .Q(n51101), .QN(
        n33125) );
  DFFRX2 dict_reg_90__0_ ( .D(n35253), .CK(clk), .RN(n42351), .Q(n50673), .QN(
        n33128) );
  DFFRX2 dict_reg_91__0_ ( .D(n35261), .CK(clk), .RN(n42352), .Q(n50674), .QN(
        n33136) );
  DFFRX2 dict_reg_91__2_ ( .D(n35259), .CK(clk), .RN(n42376), .Q(n50888), .QN(
        n33134) );
  DFFRX2 dict_reg_91__3_ ( .D(n35258), .CK(clk), .RN(n42390), .Q(n51102), .QN(
        n33133) );
  DFFRX2 dict_reg_92__0_ ( .D(n35269), .CK(clk), .RN(n42352), .Q(n50675), .QN(
        n33144) );
  DFFRX2 dict_reg_92__2_ ( .D(n35267), .CK(clk), .RN(n42376), .Q(n50889), .QN(
        n33142) );
  DFFRX2 dict_reg_92__3_ ( .D(n35266), .CK(clk), .RN(n42390), .Q(n51103), .QN(
        n33141) );
  DFFRX2 dict_reg_111__7_ ( .D(n35414), .CK(clk), .RN(n42341), .Q(n50482),
        .QN(n33289) );
  DFFRX2 dict_reg_111__0_ ( .D(n35421), .CK(clk), .RN(n42353), .Q(n50694),
        .QN(n33296) );
  DFFRX2 dict_reg_111__2_ ( .D(n35419), .CK(clk), .RN(n42378), .Q(n50908),
        .QN(n33294) );
  DFFRX2 dict_reg_119__0_ ( .D(n35485), .CK(clk), .RN(n42354), .Q(n50702),
        .QN(n33360) );
  DFFRX2 dict_reg_119__2_ ( .D(n35483), .CK(clk), .RN(n42379), .Q(n50916),
        .QN(n33358) );
  DFFRX2 dict_reg_119__3_ ( .D(n35482), .CK(clk), .RN(n42391), .Q(n51130),
        .QN(n33357) );
  DFFRX2 dict_reg_129__7_ ( .D(n35558), .CK(clk), .RN(n42342), .Q(n50498),
        .QN(n33433) );
  DFFRX2 dict_reg_130__7_ ( .D(n35566), .CK(clk), .RN(n42342), .Q(n50499),
        .QN(n33441) );
  DFFRX2 dict_reg_135__7_ ( .D(n35606), .CK(clk), .RN(n42343), .Q(n50504),
        .QN(n33481) );
  DFFRX2 dict_reg_129__0_ ( .D(n35565), .CK(clk), .RN(n42355), .Q(n50712),
        .QN(n33440) );
  DFFRX2 dict_reg_133__0_ ( .D(n35597), .CK(clk), .RN(n42355), .Q(n50716),
        .QN(n33472) );
  DFFRX2 dict_reg_138__0_ ( .D(n35637), .CK(clk), .RN(n42355), .Q(n50721),
        .QN(n33512) );
  DFFRX2 dict_reg_140__0_ ( .D(n35653), .CK(clk), .RN(n42356), .Q(n50723),
        .QN(n33528) );
  DFFRX2 dict_reg_172__0_ ( .D(n35909), .CK(clk), .RN(n42358), .Q(n50755),
        .QN(n33784) );
  DFFRX2 dict_reg_182__0_ ( .D(n35989), .CK(clk), .RN(n42359), .Q(n50765),
        .QN(n33864) );
  DFFRX2 dict_reg_194__0_ ( .D(n36085), .CK(clk), .RN(n42360), .Q(n50777),
        .QN(n33960) );
  DFFRX2 dict_reg_196__0_ ( .D(n36101), .CK(clk), .RN(n42360), .Q(n50779),
        .QN(n33976) );
  DFFRX2 dict_reg_135__2_ ( .D(n35611), .CK(clk), .RN(n42380), .Q(n50932),
        .QN(n33486) );
  DFFRX2 dict_reg_140__2_ ( .D(n35651), .CK(clk), .RN(n42380), .Q(n50937),
        .QN(n33526) );
  DFFRX2 dict_reg_194__2_ ( .D(n36083), .CK(clk), .RN(n42385), .Q(n50991),
        .QN(n33958) );
  DFFRX2 dict_reg_135__3_ ( .D(n35610), .CK(clk), .RN(n42392), .Q(n51146),
        .QN(n33485) );
  DFFRX2 dict_reg_140__3_ ( .D(n35650), .CK(clk), .RN(n42393), .Q(n51151),
        .QN(n33525) );
  DFFRX2 dict_reg_172__3_ ( .D(n35906), .CK(clk), .RN(n42396), .Q(n51183),
        .QN(n33781) );
  DFFRX2 dict_reg_194__3_ ( .D(n36082), .CK(clk), .RN(n42397), .Q(n51205),
        .QN(n33957) );
  DFFRX2 dict_reg_132__7_ ( .D(n35582), .CK(clk), .RN(n42343), .Q(n50501),
        .QN(n33457) );
  DFFRX2 dict_reg_133__7_ ( .D(n35590), .CK(clk), .RN(n42343), .Q(n50502),
        .QN(n33465) );
  DFFRX2 dict_reg_134__7_ ( .D(n35598), .CK(clk), .RN(n42343), .Q(n50503),
        .QN(n33473) );
  DFFRX2 dict_reg_136__7_ ( .D(n35614), .CK(clk), .RN(n42343), .Q(n50505),
        .QN(n33489) );
  DFFRX2 dict_reg_138__7_ ( .D(n35630), .CK(clk), .RN(n42343), .Q(n50507),
        .QN(n33505) );
  DFFRX2 dict_reg_137__0_ ( .D(n35629), .CK(clk), .RN(n42355), .Q(n50720),
        .QN(n33504) );
  DFFRX2 dict_reg_133__2_ ( .D(n35595), .CK(clk), .RN(n42380), .Q(n50930),
        .QN(n33470) );
  DFFRX2 dict_reg_138__2_ ( .D(n35635), .CK(clk), .RN(n42380), .Q(n50935),
        .QN(n33510) );
  DFFRX2 dict_reg_133__3_ ( .D(n35594), .CK(clk), .RN(n42392), .Q(n51144),
        .QN(n33469) );
  DFFRX2 dict_reg_138__3_ ( .D(n35634), .CK(clk), .RN(n42393), .Q(n51149),
        .QN(n33509) );
  DFFRX2 dict_reg_213__2_ ( .D(n36235), .CK(clk), .RN(n42387), .Q(n51010),
        .QN(n34110) );
  DFFRX2 dict_reg_146__7_ ( .D(n35694), .CK(clk), .RN(n42344), .Q(n50515),
        .QN(n33569) );
  DFFRX2 dict_reg_165__7_ ( .D(n35846), .CK(clk), .RN(n42345), .Q(n50534),
        .QN(n33721) );
  DFFRX2 dict_reg_192__7_ ( .D(n36062), .CK(clk), .RN(n42347), .Q(n50561),
        .QN(n33937) );
  DFFRX2 dict_reg_193__7_ ( .D(n36070), .CK(clk), .RN(n42347), .Q(n50562),
        .QN(n33945) );
  DFFRX2 dict_reg_153__0_ ( .D(n35757), .CK(clk), .RN(n42357), .Q(n50736),
        .QN(n33632) );
  DFFRX2 dict_reg_154__0_ ( .D(n35765), .CK(clk), .RN(n42357), .Q(n50737),
        .QN(n33640) );
  DFFRX2 dict_reg_155__0_ ( .D(n35773), .CK(clk), .RN(n42357), .Q(n50738),
        .QN(n33648) );
  DFFRX2 dict_reg_158__0_ ( .D(n35797), .CK(clk), .RN(n42357), .Q(n50741),
        .QN(n33672) );
  DFFRX2 dict_reg_159__0_ ( .D(n35805), .CK(clk), .RN(n42357), .Q(n50742),
        .QN(n33680) );
  DFFRX2 dict_reg_160__0_ ( .D(n35813), .CK(clk), .RN(n42357), .Q(n50743),
        .QN(n33688) );
  DFFRX2 dict_reg_161__0_ ( .D(n35821), .CK(clk), .RN(n42357), .Q(n50744),
        .QN(n33696) );
  DFFRX2 dict_reg_162__0_ ( .D(n35829), .CK(clk), .RN(n42357), .Q(n50745),
        .QN(n33704) );
  DFFRX2 dict_reg_168__0_ ( .D(n35877), .CK(clk), .RN(n42358), .Q(n50751),
        .QN(n33752) );
  DFFRX2 dict_reg_171__0_ ( .D(n35901), .CK(clk), .RN(n42358), .Q(n50754),
        .QN(n33776) );
  DFFRX2 dict_reg_175__0_ ( .D(n35933), .CK(clk), .RN(n42359), .Q(n50758),
        .QN(n33808) );
  DFFRX2 dict_reg_183__0_ ( .D(n35997), .CK(clk), .RN(n42359), .Q(n50766),
        .QN(n33872) );
  DFFRX2 dict_reg_208__0_ ( .D(n36197), .CK(clk), .RN(n42361), .Q(n50791),
        .QN(n34072) );
  DFFRX2 dict_reg_209__0_ ( .D(n36205), .CK(clk), .RN(n42361), .Q(n50792),
        .QN(n34080) );
  DFFRX2 dict_reg_146__2_ ( .D(n35699), .CK(clk), .RN(n42381), .Q(n50943),
        .QN(n33574) );
  DFFRX2 dict_reg_154__2_ ( .D(n35763), .CK(clk), .RN(n42382), .Q(n50951),
        .QN(n33638) );
  DFFRX2 dict_reg_158__2_ ( .D(n35795), .CK(clk), .RN(n42382), .Q(n50955),
        .QN(n33670) );
  DFFRX2 dict_reg_159__2_ ( .D(n35803), .CK(clk), .RN(n42382), .Q(n50956),
        .QN(n33678) );
  DFFRX2 dict_reg_160__2_ ( .D(n35811), .CK(clk), .RN(n42382), .Q(n50957),
        .QN(n33686) );
  DFFRX2 dict_reg_161__2_ ( .D(n35819), .CK(clk), .RN(n42382), .Q(n50958),
        .QN(n33694) );
  DFFRX2 dict_reg_162__2_ ( .D(n35827), .CK(clk), .RN(n42382), .Q(n50959),
        .QN(n33702) );
  DFFRX2 dict_reg_166__2_ ( .D(n35859), .CK(clk), .RN(n42383), .Q(n50963),
        .QN(n33734) );
  DFFRX2 dict_reg_168__2_ ( .D(n35875), .CK(clk), .RN(n42383), .Q(n50965),
        .QN(n33750) );
  DFFRX2 dict_reg_179__2_ ( .D(n35963), .CK(clk), .RN(n42384), .Q(n50976),
        .QN(n33838) );
  DFFRX2 dict_reg_183__2_ ( .D(n35995), .CK(clk), .RN(n42384), .Q(n50980),
        .QN(n33870) );
  DFFRX2 dict_reg_184__2_ ( .D(n36003), .CK(clk), .RN(n42384), .Q(n50981),
        .QN(n33878) );
  DFFRX2 dict_reg_185__2_ ( .D(n36011), .CK(clk), .RN(n42384), .Q(n50982),
        .QN(n33886) );
  DFFRX2 dict_reg_203__2_ ( .D(n36155), .CK(clk), .RN(n42386), .Q(n51000),
        .QN(n34030) );
  DFFRX2 dict_reg_204__2_ ( .D(n36163), .CK(clk), .RN(n42386), .Q(n51001),
        .QN(n34038) );
  DFFRX2 dict_reg_205__2_ ( .D(n36171), .CK(clk), .RN(n42386), .Q(n51002),
        .QN(n34046) );
  DFFRX2 dict_reg_208__2_ ( .D(n36195), .CK(clk), .RN(n42386), .Q(n51005),
        .QN(n34070) );
  DFFRX2 dict_reg_153__3_ ( .D(n35754), .CK(clk), .RN(n42394), .Q(n51164),
        .QN(n33629) );
  DFFRX2 dict_reg_154__3_ ( .D(n35762), .CK(clk), .RN(n42394), .Q(n51165),
        .QN(n33637) );
  DFFRX2 dict_reg_155__3_ ( .D(n35770), .CK(clk), .RN(n42394), .Q(n51166),
        .QN(n33645) );
  DFFRX2 dict_reg_158__3_ ( .D(n35794), .CK(clk), .RN(n42394), .Q(n51169),
        .QN(n33669) );
  DFFRX2 dict_reg_159__3_ ( .D(n35802), .CK(clk), .RN(n42394), .Q(n51170),
        .QN(n33677) );
  DFFRX2 dict_reg_160__3_ ( .D(n35810), .CK(clk), .RN(n42395), .Q(n51171),
        .QN(n33685) );
  DFFRX2 dict_reg_161__3_ ( .D(n35818), .CK(clk), .RN(n42395), .Q(n51172),
        .QN(n33693) );
  DFFRX2 dict_reg_162__3_ ( .D(n35826), .CK(clk), .RN(n42395), .Q(n51173),
        .QN(n33701) );
  DFFRX2 dict_reg_168__3_ ( .D(n35874), .CK(clk), .RN(n42395), .Q(n51179),
        .QN(n33749) );
  DFFRX2 dict_reg_183__3_ ( .D(n35994), .CK(clk), .RN(n42396), .Q(n51194),
        .QN(n33869) );
  DFFRX2 dict_reg_185__3_ ( .D(n36010), .CK(clk), .RN(n42397), .Q(n51196),
        .QN(n33885) );
  DFFRX2 dict_reg_189__3_ ( .D(n36042), .CK(clk), .RN(n42397), .Q(n51200),
        .QN(n33917) );
  DFFRX2 dict_reg_191__3_ ( .D(n36058), .CK(clk), .RN(n42397), .Q(n51202),
        .QN(n33933) );
  DFFRX2 dict_reg_208__3_ ( .D(n36194), .CK(clk), .RN(n42399), .Q(n51219),
        .QN(n34069) );
  DFFRX2 dict_reg_209__3_ ( .D(n36202), .CK(clk), .RN(n42399), .Q(n51220),
        .QN(n34077) );
  DFFRX2 dict_reg_180__0_ ( .D(n35973), .CK(clk), .RN(n42359), .Q(n50763),
        .QN(n33848) );
  DFFRX2 dict_reg_180__3_ ( .D(n35970), .CK(clk), .RN(n42396), .Q(n51191),
        .QN(n33845) );
  DFFSRX1 dict_reg_253__4_ ( .D(n36553), .CK(clk), .SN(1'b1), .RN(n37601), .Q(
        n48557), .QN(n34428) );
  DFFSRX1 dict_reg_253__7_ ( .D(n36550), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49181), .QN(n34425) );
  DFFSRX1 data_num_reg_3_ ( .D(nxt_data_num[3]), .CK(clk), .SN(1'b1), .RN(
        n37594), .Q(n50148), .QN(n32397) );
  DFFSRX1 data_queue_reg_6__1_ ( .D(n36582), .CK(clk), .SN(1'b1), .RN(n37595),
        .Q(n50164), .QN(n34489) );
  DFFSRX1 data_queue_reg_6__0_ ( .D(n36581), .CK(clk), .SN(1'b1), .RN(n37592),
        .Q(n50150), .QN(n34490) );
  DFFSRX1 data_queue_reg_6__7_ ( .D(n36588), .CK(clk), .SN(1'b1), .RN(n37598),
        .Q(n50152), .QN(n34483) );
  DFFSRX1 data_queue_reg_6__6_ ( .D(n36587), .CK(clk), .SN(1'b1), .RN(n37601),
        .Q(n50154), .QN(n34484) );
  DFFSRX1 data_queue_reg_6__5_ ( .D(n36586), .CK(clk), .SN(1'b1), .RN(n37594),
        .Q(n50156), .QN(n34485) );
  DFFSRX1 data_queue_reg_6__4_ ( .D(n36585), .CK(clk), .SN(1'b1), .RN(n37593),
        .Q(n50158), .QN(n34486) );
  DFFSRX1 data_queue_reg_6__3_ ( .D(n36584), .CK(clk), .SN(1'b1), .RN(n37598),
        .Q(n50160), .QN(n34487) );
  DFFSRX1 data_queue_reg_6__2_ ( .D(n36583), .CK(clk), .SN(1'b1), .RN(n37593),
        .Q(n50162), .QN(n34488) );
  DFFSRX1 dict_reg_254__1_ ( .D(n36564), .CK(clk), .SN(1'b1), .RN(n37592),
        .QN(n9663) );
  DFFSRX1 dict_reg_254__0_ ( .D(n36565), .CK(clk), .SN(1'b1), .RN(n37600),
        .QN(n9661) );
  DFFSRX1 codeword_reg_3_ ( .D(net152412), .CK(clk), .SN(1'b1), .RN(n42412),
        .Q(net258320), .QN(n41198) );
  DFFSRX1 state_reg_0_ ( .D(nxt_state[0]), .CK(clk), .SN(1'b1), .RN(n37596),
        .Q(state[0]), .QN(n50143) );
  DFFRX2 dict_reg_214__4_ ( .D(n36241), .CK(clk), .RN(n42411), .Q(n51438),
        .QN(n34116) );
  DFFSRX1 dict_reg_254__6_ ( .D(n36559), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n41217), .QN(n9657) );
  DFFSRX1 data_queue_reg_8__7_ ( .D(n36566), .CK(clk), .SN(1'b1), .RN(n37596),
        .Q(n50151), .QN(n34499) );
  DFFSRX1 data_queue_reg_8__6_ ( .D(n36567), .CK(clk), .SN(1'b1), .RN(n37592),
        .Q(n50153), .QN(n34500) );
  DFFSRX1 data_queue_reg_8__5_ ( .D(n36568), .CK(clk), .SN(1'b1), .RN(n37600),
        .Q(n50155), .QN(n34501) );
  DFFSRX1 data_queue_reg_8__4_ ( .D(n36569), .CK(clk), .SN(1'b1), .RN(n37592),
        .Q(n50157), .QN(n34502) );
  DFFSRX1 data_queue_reg_8__3_ ( .D(n36570), .CK(clk), .SN(1'b1), .RN(n37595),
        .Q(n50159), .QN(n34503) );
  DFFSRX1 data_queue_reg_8__2_ ( .D(n36571), .CK(clk), .SN(1'b1), .RN(n37598),
        .Q(n50161), .QN(n34504) );
  DFFSRX1 data_queue_reg_8__1_ ( .D(n36572), .CK(clk), .SN(1'b1), .RN(n37601),
        .Q(n50163), .QN(n34505) );
  DFFSRX1 data_queue_reg_8__0_ ( .D(n36637), .CK(clk), .SN(1'b1), .RN(n37593),
        .Q(n49557), .QN(n34506) );
  DFFRX2 dict_reg_152__4_ ( .D(n35745), .CK(clk), .RN(n42406), .Q(n51376),
        .QN(n33620) );
  DFFRX2 dict_reg_190__4_ ( .D(n36049), .CK(clk), .RN(n42409), .Q(n51414),
        .QN(n33924) );
  DFFRX2 dict_reg_181__4_ ( .D(n35977), .CK(clk), .RN(n42409), .Q(n51405),
        .QN(n33852) );
  DFFRX2 dict_reg_147__4_ ( .D(n35705), .CK(clk), .RN(n42406), .Q(n51371),
        .QN(n33580) );
  DFFRX2 dict_reg_167__4_ ( .D(n35865), .CK(clk), .RN(n42408), .Q(n51391),
        .QN(n33740) );
  DFFRX2 dict_reg_148__4_ ( .D(n35713), .CK(clk), .RN(n42406), .Q(n51372),
        .QN(n33588) );
  DFFRX2 dict_reg_151__4_ ( .D(n35737), .CK(clk), .RN(n42406), .Q(n51375),
        .QN(n33612) );
  DFFRX2 dict_reg_206__4_ ( .D(n36177), .CK(clk), .RN(n42411), .Q(n51430),
        .QN(n34052) );
  DFFRX2 dict_reg_156__4_ ( .D(n35777), .CK(clk), .RN(n42407), .Q(n51380),
        .QN(n33652) );
  DFFRX2 dict_reg_94__4_ ( .D(n35281), .CK(clk), .RN(n42402), .Q(n51318), .QN(
        n33156) );
  DFFRX2 dict_reg_119__4_ ( .D(n35481), .CK(clk), .RN(n42404), .Q(n51343),
        .QN(n33356) );
  DFFRX2 dict_reg_118__4_ ( .D(n35473), .CK(clk), .RN(n42403), .Q(n51342),
        .QN(n33348) );
  DFFRX2 dict_reg_121__4_ ( .D(n35497), .CK(clk), .RN(n42404), .Q(n51345),
        .QN(n33372) );
  DFFRX2 dict_reg_124__4_ ( .D(n35521), .CK(clk), .RN(n42404), .Q(n51348),
        .QN(n33396) );
  DFFRX2 dict_reg_149__4_ ( .D(n35721), .CK(clk), .RN(n42406), .Q(n51373),
        .QN(n33596) );
  DFFRX2 dict_reg_153__4_ ( .D(n35753), .CK(clk), .RN(n42406), .Q(n51377),
        .QN(n33628) );
  DFFRX2 dict_reg_158__4_ ( .D(n35793), .CK(clk), .RN(n42407), .Q(n51382),
        .QN(n33668) );
  DFFRX2 dict_reg_169__4_ ( .D(n35881), .CK(clk), .RN(n42408), .Q(n51393),
        .QN(n33756) );
  DFFRX2 dict_reg_179__4_ ( .D(n35961), .CK(clk), .RN(n42409), .Q(n51403),
        .QN(n33836) );
  DFFRX2 dict_reg_182__4_ ( .D(n35985), .CK(clk), .RN(n42409), .Q(n51406),
        .QN(n33860) );
  DFFRX2 dict_reg_202__4_ ( .D(n36145), .CK(clk), .RN(n42410), .Q(n51426),
        .QN(n34020) );
  DFFRX2 dict_reg_210__4_ ( .D(n36209), .CK(clk), .RN(n42411), .Q(n51434),
        .QN(n34084) );
  DFFRX2 dict_reg_154__4_ ( .D(n35761), .CK(clk), .RN(n42406), .Q(n51378),
        .QN(n33636) );
  DFFRX2 dict_reg_142__4_ ( .D(n35665), .CK(clk), .RN(n42405), .Q(n51366),
        .QN(n33540) );
  DFFRX2 dict_reg_204__4_ ( .D(n36161), .CK(clk), .RN(n42411), .Q(n51428),
        .QN(n34036) );
  DFFSRX1 state_reg_1_ ( .D(nxt_state[1]), .CK(clk), .SN(1'b1), .RN(n37590),
        .Q(state[1]), .QN(n50149) );
  DFFRX2 dict_reg_214__2_ ( .D(n36243), .CK(clk), .RN(n42387), .Q(n49514),
        .QN(n34118) );
  DFFRX2 dict_reg_213__4_ ( .D(n36233), .CK(clk), .RN(n42411), .Q(n51437),
        .QN(n34108) );
  DFFRX2 dict_reg_81__7_ ( .D(n35174), .CK(clk), .RN(n42339), .Q(n50455), .QN(
        n33049) );
  DFFRX2 dict_reg_82__4_ ( .D(n35185), .CK(clk), .RN(n42401), .Q(n51306), .QN(
        n33060) );
  DFFRX2 dict_reg_83__4_ ( .D(n35193), .CK(clk), .RN(n42402), .Q(n51307), .QN(
        n33068) );
  DFFRX2 dict_reg_84__4_ ( .D(n35201), .CK(clk), .RN(n42402), .Q(n51308), .QN(
        n33076) );
  DFFRX2 dict_reg_85__4_ ( .D(n35209), .CK(clk), .RN(n42402), .Q(n51309), .QN(
        n33084) );
  DFFRX2 dict_reg_86__4_ ( .D(n35217), .CK(clk), .RN(n42402), .Q(n51310), .QN(
        n33092) );
  DFFRX2 dict_reg_87__4_ ( .D(n35225), .CK(clk), .RN(n42402), .Q(n51311), .QN(
        n33100) );
  DFFRX2 dict_reg_88__4_ ( .D(n35233), .CK(clk), .RN(n42402), .Q(n51312), .QN(
        n33108) );
  DFFRX2 dict_reg_89__4_ ( .D(n35241), .CK(clk), .RN(n42402), .Q(n51313), .QN(
        n33116) );
  DFFRX2 dict_reg_90__4_ ( .D(n35249), .CK(clk), .RN(n42402), .Q(n51314), .QN(
        n33124) );
  DFFRX2 dict_reg_91__4_ ( .D(n35257), .CK(clk), .RN(n42402), .Q(n51315), .QN(
        n33132) );
  DFFRX2 dict_reg_92__4_ ( .D(n35265), .CK(clk), .RN(n42402), .Q(n51316), .QN(
        n33140) );
  DFFRX2 dict_reg_93__4_ ( .D(n35273), .CK(clk), .RN(n42402), .Q(n51317), .QN(
        n33148) );
  DFFRX2 dict_reg_114__4_ ( .D(n35441), .CK(clk), .RN(n42403), .Q(n51338),
        .QN(n33316) );
  DFFRX2 dict_reg_115__4_ ( .D(n35449), .CK(clk), .RN(n42403), .Q(n51339),
        .QN(n33324) );
  DFFRX2 dict_reg_117__4_ ( .D(n35465), .CK(clk), .RN(n42403), .Q(n51341),
        .QN(n33340) );
  DFFRX2 dict_reg_116__4_ ( .D(n35457), .CK(clk), .RN(n42403), .Q(n51340),
        .QN(n33332) );
  DFFRX2 dict_reg_120__4_ ( .D(n35489), .CK(clk), .RN(n42404), .Q(n51344),
        .QN(n33364) );
  DFFRX2 dict_reg_139__4_ ( .D(n35641), .CK(clk), .RN(n42405), .Q(n51363),
        .QN(n33516) );
  DFFRX2 dict_reg_183__4_ ( .D(n35993), .CK(clk), .RN(n42409), .Q(n51407),
        .QN(n33868) );
  DFFRX2 dict_reg_185__4_ ( .D(n36009), .CK(clk), .RN(n42409), .Q(n51409),
        .QN(n33884) );
  DFFRX2 dict_reg_203__4_ ( .D(n36153), .CK(clk), .RN(n42411), .Q(n51427),
        .QN(n34028) );
  DFFRX2 dict_reg_170__4_ ( .D(n35889), .CK(clk), .RN(n42408), .Q(n51394),
        .QN(n33764) );
  DFFRX2 dict_reg_140__4_ ( .D(n35649), .CK(clk), .RN(n42405), .Q(n51364),
        .QN(n33524) );
  DFFRX2 dict_reg_205__4_ ( .D(n36169), .CK(clk), .RN(n42411), .Q(n51429),
        .QN(n34044) );
  DFFRX2 dict_reg_141__4_ ( .D(n35657), .CK(clk), .RN(n42405), .Q(n51365),
        .QN(n33532) );
  DFFRX2 dict_reg_180__4_ ( .D(n35969), .CK(clk), .RN(n42409), .Q(n51404),
        .QN(n33844) );
  DFFSRX1 dict_reg_252__2_ ( .D(n36547), .CK(clk), .SN(1'b1), .RN(n37600), .Q(
        n41345), .QN(n34422) );
  DFFSRX1 dict_reg_252__3_ ( .D(n36546), .CK(clk), .SN(1'b1), .RN(n37599), .Q(
        n41643), .QN(n34421) );
  DFFRX1 data_queue_reg_2__5_ ( .D(n36618), .CK(clk), .RN(n42324), .Q(n36939),
        .QN(n34453) );
  DFFRX1 data_queue_reg_3__1_ ( .D(n36606), .CK(clk), .RN(n42323), .Q(n41308),
        .QN(n34465) );
  DFFRX2 dict_reg_243__1_ ( .D(n36476), .CK(clk), .RN(n42374), .Q(n41348),
        .QN(n34351) );
  DFFRX1 data_queue_reg_3__5_ ( .D(n36610), .CK(clk), .RN(n42324), .Q(n41306),
        .QN(n34461) );
  DFFRX1 data_queue_reg_3__7_ ( .D(n36612), .CK(clk), .RN(n42338), .Q(n41307),
        .QN(n36911) );
  DFFRX1 data_queue_reg_3__2_ ( .D(n36607), .CK(clk), .RN(n42323), .Q(n41288),
        .QN(n36916) );
  DFFRX2 data_queue_reg_3__4_ ( .D(n36609), .CK(clk), .RN(n42324), .Q(n41298),
        .QN(n36918) );
  DFFRX2 data_queue_reg_3__3_ ( .D(n36608), .CK(clk), .RN(n42324), .Q(n41326),
        .QN(n36913) );
  DFFRX1 data_queue_reg_0__5_ ( .D(n36634), .CK(clk), .RN(n42322), .Q(n41335),
        .QN(n34437) );
  DFFSRX1 data_queue_reg_4__6_ ( .D(n36603), .CK(clk), .SN(1'b1), .RN(n37595),
        .Q(n36732), .QN(n34468) );
  DFFRX1 data_queue_reg_1__2_ ( .D(n36623), .CK(clk), .RN(n42324), .Q(n41646),
        .QN(n34448) );
  DFFRX2 data_queue_reg_2__6_ ( .D(n36619), .CK(clk), .RN(n42337), .Q(n41629),
        .QN(n34452) );
  DFFSRX1 data_queue_reg_1__7_ ( .D(n36628), .CK(clk), .SN(1'b1), .RN(n37600),
        .Q(n36922), .QN(n34443) );
  DFFSRX1 data_queue_reg_2__0_ ( .D(n36613), .CK(clk), .SN(1'b1), .RN(n37600),
        .Q(n36920), .QN(n34458) );
  DFFSRX1 data_queue_reg_1__4_ ( .D(n36625), .CK(clk), .SN(1'b1), .RN(n37593),
        .Q(n36912), .QN(n36861) );
  DFFSRX1 dict_reg_252__0_ ( .D(n36549), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n49029), .QN(n34424) );
  DFFSRX1 dict_reg_211__6_ ( .D(n36215), .CK(clk), .SN(1'b1), .RN(n37594), .Q(
        n50376), .QN(n34090) );
  DFFSRX4 data_queue_reg_1__0_ ( .D(n36621), .CK(clk), .SN(1'b1), .RN(n37594),
        .Q(n36921), .QN(n34450) );
  DFFRX4 data_queue_reg_0__2_ ( .D(n36631), .CK(clk), .RN(n37594), .Q(
        net258261), .QN(net258262) );
  DFFSRX4 data_queue_reg_0__6_ ( .D(n36635), .CK(clk), .SN(1'b1), .RN(n37593),
        .Q(n36909), .QN(n34436) );
  DFFRX4 data_queue_reg_1__3_ ( .D(n36624), .CK(clk), .RN(n42324), .Q(n37017),
        .QN(n34447) );
  DFFSRX4 data_queue_reg_1__6_ ( .D(n36627), .CK(clk), .SN(1'b1), .RN(n37595),
        .Q(n36924), .QN(n34444) );
  DFFRX4 data_queue_reg_0__3_ ( .D(n36632), .CK(clk), .RN(n42388), .Q(n41280),
        .QN(n34439) );
  DFFSRX4 data_queue_reg_0__0_ ( .D(n36629), .CK(clk), .SN(1'b1), .RN(n37592),
        .Q(n37015), .QN(n34442) );
  DFFRX4 data_queue_reg_0__7_ ( .D(n36636), .CK(clk), .RN(n42322), .Q(n41648),
        .QN(n34435) );
  DFFSRX4 data_queue_reg_0__1_ ( .D(n36630), .CK(clk), .SN(1'b1), .RN(n37600),
        .Q(n36915), .QN(n34441) );
  DFFSRX4 data_queue_reg_1__5_ ( .D(n36626), .CK(clk), .SN(1'b1), .RN(n37593),
        .Q(n36917), .QN(n34445) );
  DFFRX4 data_queue_reg_2__4_ ( .D(n36617), .CK(clk), .RN(n42324), .Q(n41334),
        .QN(n34454) );
  DFFSRX4 data_queue_reg_2__7_ ( .D(n36620), .CK(clk), .SN(1'b1), .RN(n37596),
        .Q(n36910), .QN(n34451) );
  DFFSRX4 data_queue_reg_0__4_ ( .D(n36633), .CK(clk), .SN(1'b1), .RN(n37596),
        .Q(n36923), .QN(n34438) );
  DFFSRX4 data_queue_reg_2__1_ ( .D(n36614), .CK(clk), .SN(1'b1), .RN(n37596),
        .Q(n36908), .QN(n34457) );
  DFFSRX4 data_queue_reg_2__2_ ( .D(n36615), .CK(clk), .SN(1'b1), .RN(n37590),
        .Q(n36914), .QN(n34456) );
  DFFSRX4 dict_reg_240__7_ ( .D(n36446), .CK(clk), .SN(1'b1), .RN(n37596), .Q(
        n49232), .QN(n34321) );
  CLKAND2X3 U24849 ( .A(n40885), .B(n40886), .Y(n36638) );
  NOR2X4 U24850 ( .A(n36638), .B(n40887), .Y(n40884) );
  OA21X4 U24851 ( .A0(n11384), .A1(n11385), .B0(n11386), .Y(n36639) );
  NAND2X1 U24852 ( .A(n36639), .B(n11387), .Y(n11381) );
  AO21X4 U24853 ( .A0(n11380), .A1(n11381), .B0(net151857), .Y(n41214) );
  OR2X6 U24854 ( .A(n47767), .B(n47766), .Y(n36640) );
  NAND2X2 U24855 ( .A(n36640), .B(n41762), .Y(n47768) );
  NOR2X4 U24856 ( .A(n47765), .B(net210522), .Y(n47767) );
  NAND2X2 U24857 ( .A(n47990), .B(n47979), .Y(n47766) );
  CLKAND2X6 U24858 ( .A(n47989), .B(n47995), .Y(n41762) );
  OAI2BB1X4 U24859 ( .A0N(net234521), .A1N(n47768), .B0(net234523), .Y(n47769)
         );
  NAND3X1 U24860 ( .A(n45307), .B(n45305), .C(n45306), .Y(n36641) );
  NAND2X4 U24861 ( .A(n36642), .B(n45308), .Y(net209631) );
  CLKINVX1 U24862 ( .A(n36641), .Y(n36642) );
  OR2X2 U24863 ( .A(n40539), .B(net171544), .Y(n36643) );
  NAND2X1 U24864 ( .A(n36643), .B(n40719), .Y(n40463) );
  NAND4BBX2 U24865 ( .AN(n40461), .BN(n40462), .C(n40463), .D(n40464), .Y(
        n34515) );
  NAND3X1 U24866 ( .A(n44545), .B(n44543), .C(n44544), .Y(n36644) );
  NAND2X2 U24867 ( .A(n36645), .B(n44546), .Y(n12506) );
  CLKINVX1 U24868 ( .A(n36644), .Y(n36645) );
  AO21X1 U24869 ( .A0(n48276), .A1(n12506), .B0(n49505), .Y(n41664) );
  NAND2X1 U24870 ( .A(net215421), .B(n39457), .Y(n36646) );
  NAND2X4 U24871 ( .A(n36647), .B(net215420), .Y(n10393) );
  INVX3 U24872 ( .A(n36646), .Y(n36647) );
  NOR4X1 U24873 ( .A(n27508), .B(n27509), .C(n27510), .D(n27511), .Y(net215420) );
  NAND3X1 U24874 ( .A(n45911), .B(n45912), .C(n45913), .Y(n36648) );
  NAND2X1 U24875 ( .A(n36649), .B(n45914), .Y(n11057) );
  CLKINVX1 U24876 ( .A(n36648), .Y(n36649) );
  NAND3X1 U24877 ( .A(n44605), .B(n44604), .C(n44603), .Y(n36650) );
  NAND2X2 U24878 ( .A(n36651), .B(n44606), .Y(n11744) );
  CLKINVX1 U24879 ( .A(n36650), .Y(n36651) );
  NAND2X1 U24880 ( .A(n43802), .B(n43801), .Y(n36652) );
  NAND3X2 U24881 ( .A(n43804), .B(n43803), .C(n36653), .Y(n12032) );
  CLKINVX1 U24882 ( .A(n36652), .Y(n36653) );
  XNOR2XL U24883 ( .A(n33546), .B(n42569), .Y(n43803) );
  NOR2X1 U24884 ( .A(n27539), .B(n27540), .Y(n36654) );
  NOR3X2 U24885 ( .A(n27541), .B(n36655), .C(n27538), .Y(net215429) );
  CLKINVX1 U24886 ( .A(n36654), .Y(n36655) );
  XOR2XL U24887 ( .A(n41855), .B(n42609), .Y(n27541) );
  NAND3X1 U24888 ( .A(n47094), .B(n47095), .C(n47096), .Y(n36656) );
  NAND2X1 U24889 ( .A(n36657), .B(n47097), .Y(n11365) );
  CLKINVX1 U24890 ( .A(n36656), .Y(n36657) );
  NAND3X6 U24891 ( .A(n11365), .B(n11366), .C(n11367), .Y(n11362) );
  NAND3X1 U24892 ( .A(n45759), .B(n45760), .C(n45761), .Y(n36658) );
  NAND2X2 U24893 ( .A(n36659), .B(n45762), .Y(n11092) );
  CLKINVX1 U24894 ( .A(n36658), .Y(n36659) );
  OAI211X2 U24895 ( .A0(n11090), .A1(n11091), .B0(n11092), .C0(n40398), .Y(
        n11087) );
  NAND2X1 U24896 ( .A(n10368), .B(n10369), .Y(n36660) );
  NAND2X2 U24897 ( .A(n36661), .B(n11738), .Y(n11735) );
  CLKINVX1 U24898 ( .A(n36660), .Y(n36661) );
  NAND3X1 U24899 ( .A(net215227), .B(n39452), .C(net215228), .Y(n10368) );
  OR2X2 U24900 ( .A(n40608), .B(n40493), .Y(n36662) );
  NAND2X2 U24901 ( .A(n36662), .B(n40610), .Y(n40499) );
  NAND2X1 U24902 ( .A(n42129), .B(n36664), .Y(n36665) );
  NAND2XL U24903 ( .A(n36663), .B(n42653), .Y(n36666) );
  NAND2X1 U24904 ( .A(n36665), .B(n36666), .Y(n29259) );
  CLKINVX1 U24905 ( .A(n42129), .Y(n36663) );
  CLKINVX1 U24906 ( .A(n42653), .Y(n36664) );
  BUFX4 U24907 ( .A(n42668), .Y(n42653) );
  OR2X2 U24908 ( .A(n48148), .B(net258199), .Y(n36667) );
  NAND2X2 U24909 ( .A(n36667), .B(n48146), .Y(n48152) );
  NAND2X2 U24910 ( .A(n48306), .B(n46505), .Y(n48146) );
  AOI21X1 U24911 ( .A0(n48152), .A1(n48151), .B0(n48150), .Y(n48153) );
  NAND2X1 U24912 ( .A(n46319), .B(n46317), .Y(n36668) );
  NAND3X4 U24913 ( .A(n46320), .B(n46318), .C(n36669), .Y(net209325) );
  CLKINVX1 U24914 ( .A(n36668), .Y(n36669) );
  NOR2X1 U24915 ( .A(n46310), .B(net209902), .Y(n46320) );
  NOR2X1 U24916 ( .A(n47314), .B(net209325), .Y(n47324) );
  CLKINVX1 U24917 ( .A(net209325), .Y(net209315) );
  OA21X4 U24918 ( .A0(n11374), .A1(n11375), .B0(n11376), .Y(n36670) );
  NAND2X6 U24919 ( .A(n36670), .B(n11377), .Y(n11373) );
  NOR2X4 U24920 ( .A(n41214), .B(net151860), .Y(n11374) );
  NAND2X2 U24921 ( .A(n11378), .B(n11379), .Y(n11375) );
  NAND4X6 U24922 ( .A(n46909), .B(n46908), .C(n46907), .D(n46906), .Y(n11376)
         );
  NAND4X6 U24923 ( .A(n46914), .B(n46913), .C(n46912), .D(n46911), .Y(n11377)
         );
  NAND3X6 U24924 ( .A(n11371), .B(n11372), .C(n11373), .Y(n11370) );
  OR2X6 U24925 ( .A(n47789), .B(net210537), .Y(n36671) );
  NAND2X6 U24926 ( .A(n36671), .B(net210536), .Y(n47790) );
  NAND2X8 U24927 ( .A(net209284), .B(net209277), .Y(net210537) );
  CLKINVX12 U24928 ( .A(net210561), .Y(net210536) );
  NAND2X2 U24929 ( .A(n41868), .B(n36673), .Y(n36674) );
  NAND2XL U24930 ( .A(n36672), .B(n42600), .Y(n36675) );
  NAND2X4 U24931 ( .A(n36674), .B(n36675), .Y(n29315) );
  INVXL U24932 ( .A(n41868), .Y(n36672) );
  CLKINVX1 U24933 ( .A(n42600), .Y(n36673) );
  CLKBUFX6 U24934 ( .A(n33911), .Y(n41868) );
  CLKAND2X3 U24935 ( .A(n41189), .B(n41054), .Y(n36676) );
  NOR2X2 U24936 ( .A(n36676), .B(n41188), .Y(n40804) );
  NAND2X2 U24937 ( .A(n45214), .B(n45216), .Y(n36677) );
  NAND3X4 U24938 ( .A(n45215), .B(n45213), .C(n36678), .Y(n48301) );
  CLKINVX3 U24939 ( .A(n36677), .Y(n36678) );
  NOR4X2 U24940 ( .A(n45204), .B(n45203), .C(n45202), .D(n45201), .Y(n45215)
         );
  NOR2X4 U24941 ( .A(n45217), .B(n48301), .Y(n45227) );
  OR2X2 U24942 ( .A(n47983), .B(n47982), .Y(n36679) );
  NAND2X2 U24943 ( .A(n36679), .B(n47981), .Y(n47985) );
  NAND3X8 U24944 ( .A(n47707), .B(n47706), .C(n48437), .Y(n47981) );
  AOI21X1 U24945 ( .A0(n47985), .A1(n47984), .B0(net210216), .Y(n47986) );
  NAND2X2 U24946 ( .A(n41854), .B(n36681), .Y(n36682) );
  NAND2XL U24947 ( .A(n36680), .B(n42609), .Y(n36683) );
  NAND2X2 U24948 ( .A(n36682), .B(n36683), .Y(n27511) );
  CLKINVX1 U24949 ( .A(n41854), .Y(n36680) );
  INVX1 U24950 ( .A(n42609), .Y(n36681) );
  OA21X4 U24951 ( .A0(n11145), .A1(n11146), .B0(n11147), .Y(n36684) );
  NAND2X4 U24952 ( .A(n36684), .B(n11148), .Y(n11142) );
  AOI21X4 U24953 ( .A0(net210557), .A1(n47790), .B0(net210559), .Y(n11145) );
  NAND4X8 U24954 ( .A(n46188), .B(n46187), .C(n46186), .D(n46185), .Y(n11148)
         );
  OA21X4 U24955 ( .A0(n11312), .A1(n11313), .B0(n11314), .Y(n36685) );
  NAND2X6 U24956 ( .A(n36685), .B(n11315), .Y(n11309) );
  AOI211X2 U24957 ( .A0(n11318), .A1(n11319), .B0(n36943), .C0(n39626), .Y(
        n11312) );
  NAND2X2 U24958 ( .A(n11316), .B(n11317), .Y(n11313) );
  NAND4X2 U24959 ( .A(n46813), .B(n46812), .C(n46811), .D(n46810), .Y(n11314)
         );
  NAND4X8 U24960 ( .A(n46818), .B(n46817), .C(n46816), .D(n46815), .Y(n11315)
         );
  NOR2X6 U24961 ( .A(n11309), .B(n40829), .Y(n40828) );
  OR2X8 U24962 ( .A(n47715), .B(net210442), .Y(n36686) );
  NAND2X8 U24963 ( .A(n36686), .B(n47714), .Y(n47717) );
  AOI21X4 U24964 ( .A0(net234998), .A1(n47713), .B0(net210698), .Y(n47715) );
  NAND2XL U24965 ( .A(n48156), .B(n48158), .Y(net210442) );
  NAND3X1 U24966 ( .A(n46409), .B(n46408), .C(n46410), .Y(n36687) );
  NAND2X2 U24967 ( .A(n36688), .B(n46411), .Y(net209290) );
  CLKINVX1 U24968 ( .A(n36687), .Y(n36688) );
  NOR2X4 U24969 ( .A(n47413), .B(net209290), .Y(n47423) );
  INVX1 U24970 ( .A(net209290), .Y(net210567) );
  OR2X6 U24971 ( .A(n40489), .B(net151773), .Y(n36689) );
  NAND2X6 U24972 ( .A(n36689), .B(n12596), .Y(n40763) );
  AOI21X4 U24973 ( .A0(n40490), .A1(net271431), .B0(net171259), .Y(n40489) );
  INVX12 U24974 ( .A(n10448), .Y(net151773) );
  NAND2BX4 U24975 ( .AN(n40459), .B(net212567), .Y(n12596) );
  NAND2X6 U24976 ( .A(net260394), .B(n40763), .Y(n40758) );
  NAND3X2 U24977 ( .A(n44279), .B(n44280), .C(n44278), .Y(n36690) );
  NAND2X2 U24978 ( .A(n36691), .B(n44281), .Y(n12584) );
  INVX3 U24979 ( .A(n36690), .Y(n36691) );
  NOR3X1 U24980 ( .A(n26796), .B(n37207), .C(n26795), .Y(n44279) );
  NOR2X4 U24981 ( .A(n12584), .B(n44282), .Y(n44286) );
  NAND4XL U24982 ( .A(n11850), .B(n11849), .C(n12530), .D(n12584), .Y(n10113)
         );
  INVXL U24983 ( .A(n12584), .Y(n49503) );
  OAI21X2 U24984 ( .A0(n49507), .A1(n48285), .B0(n12584), .Y(n48287) );
  OR2X6 U24985 ( .A(net210058), .B(n48105), .Y(n36692) );
  NAND2X6 U24986 ( .A(n36692), .B(n11327), .Y(n48106) );
  INVX3 U24987 ( .A(n11326), .Y(net210058) );
  AOI21X4 U24988 ( .A0(n48104), .A1(n12893), .B0(net151445), .Y(n48105) );
  NAND4X8 U24989 ( .A(n46894), .B(n46893), .C(n46892), .D(n46891), .Y(n11327)
         );
  AOI21X4 U24990 ( .A0(n48106), .A1(n11324), .B0(net210057), .Y(n48107) );
  NAND3X1 U24991 ( .A(n46164), .B(n46165), .C(n46166), .Y(n36693) );
  NAND2X2 U24992 ( .A(n36694), .B(n46167), .Y(n11115) );
  CLKINVX1 U24993 ( .A(n36693), .Y(n36694) );
  NOR2X4 U24994 ( .A(n12064), .B(n46163), .Y(n46167) );
  OAI2BB1XL U24995 ( .A0N(n11115), .A1N(net209234), .B0(n12318), .Y(n48498) );
  INVXL U24996 ( .A(n11115), .Y(n39408) );
  NAND2X4 U24997 ( .A(n41356), .B(n11115), .Y(n11109) );
  NAND2X6 U24998 ( .A(n47738), .B(n47737), .Y(n36695) );
  INVX6 U24999 ( .A(n47736), .Y(n36696) );
  AND2X8 U25000 ( .A(n36695), .B(n36696), .Y(n47741) );
  NOR2BX1 U25001 ( .AN(net209604), .B(net209633), .Y(n47738) );
  OAI2BB1X4 U25002 ( .A0N(n47735), .A1N(n47734), .B0(n47733), .Y(n47737) );
  NAND2XL U25003 ( .A(net209602), .B(net209631), .Y(n47736) );
  NOR3X2 U25004 ( .A(n45029), .B(n45030), .C(n45031), .Y(n36697) );
  NOR2X2 U25005 ( .A(n45032), .B(n36698), .Y(n45043) );
  CLKINVX1 U25006 ( .A(n36697), .Y(n36698) );
  XOR2XL U25007 ( .A(n34423), .B(n42607), .Y(n45032) );
  XOR2XL U25008 ( .A(n34424), .B(n42592), .Y(n45031) );
  NAND2X4 U25009 ( .A(n34321), .B(n36700), .Y(n36701) );
  NAND2XL U25010 ( .A(n36699), .B(n41379), .Y(n36702) );
  NAND2X4 U25011 ( .A(n36701), .B(n36702), .Y(n45424) );
  INVXL U25012 ( .A(n34321), .Y(n36699) );
  INVXL U25013 ( .A(n41379), .Y(n36700) );
  NOR4X4 U25014 ( .A(n45424), .B(n45423), .C(n45422), .D(n45421), .Y(n45435)
         );
  NAND2X6 U25015 ( .A(n41806), .B(n36704), .Y(n36705) );
  NAND2X2 U25016 ( .A(n36703), .B(n42607), .Y(n36706) );
  NAND2X6 U25017 ( .A(n36705), .B(n36706), .Y(n45017) );
  CLKINVX1 U25018 ( .A(n41806), .Y(n36703) );
  INVX2 U25019 ( .A(n42607), .Y(n36704) );
  BUFX8 U25020 ( .A(n34415), .Y(n41806) );
  NOR4X4 U25021 ( .A(n45018), .B(n45017), .C(n45016), .D(n45015), .Y(n45019)
         );
  NOR2X6 U25022 ( .A(n12033), .B(n45833), .Y(n45837) );
  OAI2BB1X4 U25023 ( .A0N(n12032), .A1N(n41689), .B0(n12033), .Y(n48122) );
  NAND4X4 U25024 ( .A(n43813), .B(n43812), .C(n43811), .D(n43810), .Y(n12033)
         );
  CLKINVX8 U25025 ( .A(n42721), .Y(n36707) );
  INVX4 U25026 ( .A(n36707), .Y(n36708) );
  CLKINVX12 U25027 ( .A(n36707), .Y(n36709) );
  NOR4X2 U25028 ( .A(n45420), .B(n45419), .C(n45418), .D(n45417), .Y(n45436)
         );
  XOR2X1 U25029 ( .A(n34326), .B(n42615), .Y(n45419) );
  CLKBUFX3 U25030 ( .A(n42603), .Y(n36710) );
  CLKBUFX3 U25031 ( .A(n42603), .Y(n36711) );
  CLKBUFX2 U25032 ( .A(n42611), .Y(n42603) );
  OAI21X2 U25033 ( .A0(n40890), .A1(n41001), .B0(n41003), .Y(n41195) );
  AOI21X4 U25034 ( .A0(n40891), .A1(n40892), .B0(n40893), .Y(n40890) );
  AND2XL U25035 ( .A(n11082), .B(n11210), .Y(n48510) );
  AND2XL U25036 ( .A(n11210), .B(n11211), .Y(n11076) );
  CLKINVX4 U25037 ( .A(n11210), .Y(net209211) );
  NAND3XL U25038 ( .A(n11210), .B(n12292), .C(n39433), .Y(n10242) );
  NAND4X2 U25039 ( .A(n45832), .B(n45831), .C(n45830), .D(n45829), .Y(n11210)
         );
  NOR2X6 U25040 ( .A(n40830), .B(n40833), .Y(n40832) );
  NOR2X2 U25041 ( .A(n40828), .B(n40831), .Y(n40830) );
  INVX8 U25042 ( .A(n10367), .Y(net171249) );
  NOR2XL U25043 ( .A(n10367), .B(n44277), .Y(net215271) );
  NAND4BX4 U25044 ( .AN(n37304), .B(net215279), .C(net215276), .D(net215277),
        .Y(n10367) );
  CLKINVX1 U25045 ( .A(n36712), .Y(n36713) );
  CLKBUFX6 U25046 ( .A(n36713), .Y(n36714) );
  CLKBUFX6 U25047 ( .A(n36713), .Y(n36715) );
  CLKBUFX6 U25048 ( .A(n36713), .Y(n36716) );
  CLKBUFX6 U25049 ( .A(n36713), .Y(n36717) );
  CLKBUFX6 U25050 ( .A(n36713), .Y(n36718) );
  CLKINVX1 U25051 ( .A(n34471), .Y(n36719) );
  INVX6 U25052 ( .A(n36719), .Y(n36720) );
  INVX6 U25053 ( .A(n36719), .Y(n36721) );
  INVX6 U25054 ( .A(n36719), .Y(n36722) );
  NAND2X1 U25055 ( .A(net209341), .B(net209301), .Y(net210544) );
  NAND4X4 U25056 ( .A(n46444), .B(n46443), .C(n46442), .D(n46441), .Y(
        net209301) );
  NOR2X6 U25057 ( .A(n45853), .B(net209800), .Y(n45857) );
  INVX1 U25058 ( .A(net209800), .Y(net171210) );
  NAND4X4 U25059 ( .A(n43759), .B(n43758), .C(n43757), .D(n43756), .Y(
        net209800) );
  CLKXOR2X2 U25060 ( .A(n34377), .B(n42680), .Y(n44917) );
  AOI21X2 U25061 ( .A0(n48240), .A1(n48239), .B0(n48238), .Y(n48247) );
  OAI21X1 U25062 ( .A0(n48233), .A1(n48232), .B0(n48231), .Y(n48239) );
  INVX3 U25063 ( .A(n42566), .Y(n36723) );
  CLKINVX1 U25064 ( .A(n36723), .Y(n36724) );
  INVX2 U25065 ( .A(n36723), .Y(n36725) );
  INVX3 U25066 ( .A(n36723), .Y(n36726) );
  AO21X2 U25067 ( .A0(n48092), .A1(n48091), .B0(n48090), .Y(n41702) );
  OAI21X1 U25068 ( .A0(n48083), .A1(n48082), .B0(n48081), .Y(n48091) );
  INVX6 U25069 ( .A(n42682), .Y(n36727) );
  CLKINVX16 U25070 ( .A(n36727), .Y(n36728) );
  INVX4 U25071 ( .A(net209623), .Y(net212262) );
  NAND4X4 U25072 ( .A(n45044), .B(n45043), .C(n45042), .D(n45041), .Y(
        net209623) );
  NAND3X8 U25073 ( .A(net215352), .B(net215353), .C(n39317), .Y(n10566) );
  NOR2X6 U25074 ( .A(n12542), .B(n44228), .Y(net215352) );
  NAND4X4 U25075 ( .A(n46122), .B(n46121), .C(n46120), .D(n46119), .Y(
        net209249) );
  NOR2X1 U25076 ( .A(n12736), .B(n46118), .Y(n46122) );
  AOI21X2 U25077 ( .A0(n48297), .A1(n11777), .B0(net209638), .Y(n48347) );
  NOR2X8 U25078 ( .A(n11777), .B(n44182), .Y(n44186) );
  NAND3XL U25079 ( .A(n11777), .B(n12582), .C(n39464), .Y(n10419) );
  NAND4X4 U25080 ( .A(n44181), .B(n44180), .C(n44179), .D(n44178), .Y(n11777)
         );
  NOR4X4 U25081 ( .A(n28290), .B(n28291), .C(n28292), .D(n28293), .Y(n43754)
         );
  CLKXOR2X1 U25082 ( .A(n41923), .B(n42600), .Y(n28293) );
  OAI31X2 U25083 ( .A0(n11424), .A1(net171555), .A2(net171554), .B0(n10715),
        .Y(n11419) );
  NOR2X2 U25084 ( .A(n41226), .B(net151600), .Y(n11424) );
  NAND4X4 U25085 ( .A(n45436), .B(n45435), .C(n45434), .D(n45433), .Y(
        net209635) );
  NOR2X6 U25086 ( .A(n10870), .B(n47892), .Y(n47896) );
  AND2XL U25087 ( .A(n10872), .B(n10870), .Y(n11133) );
  INVXL U25088 ( .A(n10870), .Y(net209255) );
  NAND2BX4 U25089 ( .AN(n39424), .B(net213347), .Y(n10870) );
  CLKBUFX2 U25090 ( .A(n42677), .Y(n42678) );
  CLKINVX20 U25091 ( .A(n42500), .Y(n36729) );
  CLKINVX20 U25092 ( .A(n36729), .Y(n36730) );
  CLKINVX20 U25093 ( .A(n36729), .Y(n36731) );
  NAND3X8 U25094 ( .A(n39419), .B(net212466), .C(net212463), .Y(net209343) );
  NOR2X6 U25095 ( .A(n46383), .B(n48159), .Y(net212463) );
  NAND4X6 U25096 ( .A(n46107), .B(n46106), .C(n46105), .D(n46104), .Y(n12384)
         );
  NOR2X6 U25097 ( .A(n12145), .B(n46103), .Y(n46107) );
  NAND2X4 U25098 ( .A(net210222), .B(net210207), .Y(net210522) );
  NAND4X4 U25099 ( .A(n47589), .B(n47588), .C(n47587), .D(n47586), .Y(
        net210222) );
  INVX12 U25100 ( .A(n36732), .Y(n36733) );
  INVX12 U25101 ( .A(n36732), .Y(n36734) );
  BUFX12 U25102 ( .A(n34468), .Y(n36735) );
  BUFX12 U25103 ( .A(n34468), .Y(n36736) );
  AOI211X2 U25104 ( .A0(n11406), .A1(n11407), .B0(net151753), .C0(net151750),
        .Y(n11404) );
  NOR2BXL U25105 ( .AN(n12940), .B(n37253), .Y(n48068) );
  AND4X4 U25106 ( .A(n47158), .B(n47157), .C(n47156), .D(n47155), .Y(n37253)
         );
  XNOR2X4 U25107 ( .A(n50987), .B(n41284), .Y(n29162) );
  CLKINVX6 U25108 ( .A(n42622), .Y(n41284) );
  BUFX20 U25109 ( .A(n42507), .Y(n36737) );
  NOR4X2 U25110 ( .A(n44140), .B(n44139), .C(n44138), .D(n44137), .Y(n44151)
         );
  CLKXOR2X1 U25111 ( .A(n34193), .B(n36903), .Y(n44140) );
  NAND4X4 U25112 ( .A(n44121), .B(n44120), .C(n44119), .D(n44118), .Y(
        net209595) );
  NOR4X4 U25113 ( .A(n44109), .B(n44108), .C(n44107), .D(n44106), .Y(n44120)
         );
  BUFX2 U25114 ( .A(n36921), .Y(n42593) );
  INVX20 U25115 ( .A(n36862), .Y(n36863) );
  INVX12 U25116 ( .A(n42593), .Y(n42591) );
  NAND3X6 U25117 ( .A(n47673), .B(n47672), .C(net210749), .Y(n47982) );
  NOR4X2 U25118 ( .A(n47667), .B(n47666), .C(n47665), .D(n47664), .Y(n47673)
         );
  INVX8 U25119 ( .A(n42645), .Y(n42637) );
  CLKINVX20 U25120 ( .A(n36866), .Y(n36867) );
  OAI21X4 U25121 ( .A0(n40858), .A1(n41022), .B0(n41024), .Y(n41193) );
  NOR2X8 U25122 ( .A(n11627), .B(n40859), .Y(n40858) );
  OAI21X2 U25123 ( .A0(n11972), .A1(n40945), .B0(n40972), .Y(n41194) );
  OAI211X2 U25124 ( .A0(n11974), .A1(n11975), .B0(n11976), .C0(n11977), .Y(
        n11972) );
  CLKBUFX12 U25125 ( .A(n36873), .Y(n41323) );
  NAND2XL U25126 ( .A(n12741), .B(n12744), .Y(n10572) );
  NOR2X8 U25127 ( .A(n12741), .B(n47036), .Y(n47040) );
  NAND4X8 U25128 ( .A(n44216), .B(n44215), .C(n44214), .D(n44213), .Y(n12741)
         );
  NAND4X6 U25129 ( .A(n45726), .B(n45725), .C(n45724), .D(n45723), .Y(n11209)
         );
  NOR2X6 U25130 ( .A(n12708), .B(n45722), .Y(n45726) );
  XNOR2X4 U25131 ( .A(n50773), .B(n42586), .Y(n29164) );
  CLKINVX4 U25132 ( .A(n42594), .Y(n42586) );
  INVX20 U25133 ( .A(net219480), .Y(net219442) );
  CLKBUFX6 U25134 ( .A(net219472), .Y(net219480) );
  AND4XL U25135 ( .A(n10382), .B(n10384), .C(n10383), .D(n10381), .Y(n24717)
         );
  AOI21X2 U25136 ( .A0(n48351), .A1(n10381), .B0(net209543), .Y(n48353) );
  NOR2X6 U25137 ( .A(n10381), .B(n44229), .Y(n44233) );
  NAND3X4 U25138 ( .A(net215348), .B(net215349), .C(n39456), .Y(n10381) );
  AOI211X2 U25139 ( .A0(n11352), .A1(n11353), .B0(n39631), .C0(n36942), .Y(
        n11346) );
  NOR4X4 U25140 ( .A(n44649), .B(n44648), .C(n44647), .D(n44646), .Y(n44660)
         );
  CLKXOR2X1 U25141 ( .A(n34217), .B(n36903), .Y(n44649) );
  CLKINVX3 U25142 ( .A(n36914), .Y(n42544) );
  CLKINVX8 U25143 ( .A(n36914), .Y(n42533) );
  INVX12 U25144 ( .A(n36914), .Y(n42534) );
  CLKINVX6 U25145 ( .A(n36914), .Y(n42542) );
  CLKINVX3 U25146 ( .A(n36914), .Y(n42536) );
  NAND2BX4 U25147 ( .AN(n39416), .B(net212385), .Y(net209344) );
  NOR2X6 U25148 ( .A(n46456), .B(n48160), .Y(net212385) );
  NAND3XL U25149 ( .A(net210615), .B(net210209), .C(net210213), .Y(net210525)
         );
  CLKINVX8 U25150 ( .A(net210209), .Y(net210617) );
  NAND4X6 U25151 ( .A(n47633), .B(n47632), .C(n47631), .D(n47630), .Y(
        net210209) );
  CLKINVX16 U25152 ( .A(net219356), .Y(net219310) );
  NAND2X4 U25153 ( .A(n47984), .B(n47981), .Y(n47761) );
  BUFX20 U25154 ( .A(n42679), .Y(n42677) );
  INVX3 U25155 ( .A(n36738), .Y(n36739) );
  BUFX4 U25156 ( .A(n36739), .Y(n36740) );
  BUFX4 U25157 ( .A(n36739), .Y(n36741) );
  BUFX4 U25158 ( .A(n36739), .Y(n36742) );
  BUFX4 U25159 ( .A(n36739), .Y(n36743) );
  BUFX4 U25160 ( .A(n36739), .Y(n36744) );
  CLKBUFX3 U25161 ( .A(n34470), .Y(n36745) );
  CLKBUFX8 U25162 ( .A(n36745), .Y(n36746) );
  CLKBUFX8 U25163 ( .A(n36745), .Y(n36747) );
  CLKBUFX6 U25164 ( .A(n36745), .Y(n36748) );
  CLKBUFX6 U25165 ( .A(n36745), .Y(n36749) );
  BUFX4 U25166 ( .A(n36745), .Y(n36750) );
  INVX8 U25167 ( .A(net213678), .Y(net209617) );
  AND2XL U25168 ( .A(net213678), .B(net213679), .Y(n41752) );
  NAND4XL U25169 ( .A(net213678), .B(net210477), .C(net209615), .D(net213679),
        .Y(n39707) );
  NAND4BX4 U25170 ( .AN(n41709), .B(n45079), .C(n45078), .D(n45077), .Y(
        net213678) );
  INVX3 U25171 ( .A(n36751), .Y(n36752) );
  CLKBUFX6 U25172 ( .A(n36752), .Y(n36753) );
  CLKBUFX6 U25173 ( .A(n36752), .Y(n36754) );
  CLKBUFX6 U25174 ( .A(n36752), .Y(n36755) );
  CLKBUFX6 U25175 ( .A(n36752), .Y(n36756) );
  CLKBUFX6 U25176 ( .A(n36752), .Y(n36757) );
  INVX1 U25177 ( .A(n34473), .Y(n36758) );
  INVX6 U25178 ( .A(n36758), .Y(n36759) );
  INVX6 U25179 ( .A(n36758), .Y(n36760) );
  INVX6 U25180 ( .A(n36758), .Y(n36761) );
  CLKBUFX2 U25181 ( .A(n34457), .Y(n42514) );
  BUFX8 U25182 ( .A(n34457), .Y(n42513) );
  INVX3 U25183 ( .A(n36762), .Y(n36763) );
  BUFX4 U25184 ( .A(n36763), .Y(n36764) );
  BUFX4 U25185 ( .A(n36763), .Y(n36765) );
  BUFX4 U25186 ( .A(n36763), .Y(n36766) );
  BUFX4 U25187 ( .A(n36763), .Y(n36767) );
  CLKBUFX6 U25188 ( .A(n36763), .Y(n36768) );
  CLKBUFX3 U25189 ( .A(n34467), .Y(n36769) );
  BUFX4 U25190 ( .A(n36769), .Y(n36770) );
  BUFX4 U25191 ( .A(n36769), .Y(n36771) );
  BUFX4 U25192 ( .A(n36769), .Y(n36772) );
  BUFX4 U25193 ( .A(n36769), .Y(n36773) );
  BUFX4 U25194 ( .A(n36769), .Y(n36774) );
  INVX1 U25195 ( .A(net219480), .Y(net219444) );
  NOR2BXL U25196 ( .AN(net209636), .B(net209634), .Y(n47733) );
  NOR2X4 U25197 ( .A(n45485), .B(net209636), .Y(net213731) );
  NAND4BX4 U25198 ( .AN(n41683), .B(n45484), .C(n45483), .D(n45482), .Y(
        net209636) );
  CLKBUFX3 U25199 ( .A(n36911), .Y(n36775) );
  CLKBUFX6 U25200 ( .A(n36775), .Y(n36776) );
  CLKBUFX6 U25201 ( .A(n36775), .Y(n36777) );
  CLKBUFX6 U25202 ( .A(n36775), .Y(n36778) );
  CLKBUFX6 U25203 ( .A(n36775), .Y(n36779) );
  BUFX4 U25204 ( .A(n36775), .Y(n36780) );
  INVX6 U25205 ( .A(n41307), .Y(n36781) );
  BUFX16 U25206 ( .A(n36781), .Y(n36782) );
  BUFX12 U25207 ( .A(n36781), .Y(n36783) );
  BUFX8 U25208 ( .A(n36781), .Y(n36784) );
  BUFX8 U25209 ( .A(n36781), .Y(n36785) );
  BUFX4 U25210 ( .A(n36781), .Y(n36786) );
  CLKBUFX4 U25211 ( .A(n42610), .Y(n42600) );
  AOI21X4 U25212 ( .A0(n40487), .A1(n11885), .B0(n40488), .Y(n40486) );
  OAI21X2 U25213 ( .A0(net151786), .A1(n40485), .B0(n12602), .Y(n40487) );
  BUFX3 U25214 ( .A(n34438), .Y(n42692) );
  CLKINVX6 U25215 ( .A(n42677), .Y(n42672) );
  OAI21X2 U25216 ( .A0(n40866), .A1(n41045), .B0(n41046), .Y(n40872) );
  AOI21X4 U25217 ( .A0(n40867), .A1(n40868), .B0(n40869), .Y(n40866) );
  NOR2X6 U25218 ( .A(n47424), .B(net209312), .Y(n47434) );
  AND2XL U25219 ( .A(net209312), .B(net209343), .Y(n41764) );
  NAND2XL U25220 ( .A(net209312), .B(net209343), .Y(n39945) );
  NAND2X4 U25221 ( .A(n39418), .B(net212474), .Y(net209312) );
  NOR4X2 U25222 ( .A(n45111), .B(n45110), .C(n45109), .D(n45108), .Y(n45125)
         );
  CLKBUFX12 U25223 ( .A(n41288), .Y(n41289) );
  INVX3 U25224 ( .A(n36787), .Y(n36788) );
  BUFX4 U25225 ( .A(n36788), .Y(n36789) );
  BUFX4 U25226 ( .A(n36788), .Y(n36790) );
  BUFX4 U25227 ( .A(n36788), .Y(n36791) );
  BUFX4 U25228 ( .A(n36788), .Y(n36792) );
  BUFX4 U25229 ( .A(n36788), .Y(n36793) );
  CLKBUFX3 U25230 ( .A(n34472), .Y(n36794) );
  BUFX4 U25231 ( .A(n36794), .Y(n36795) );
  BUFX4 U25232 ( .A(n36794), .Y(n36796) );
  BUFX4 U25233 ( .A(n36794), .Y(n36797) );
  BUFX4 U25234 ( .A(n36794), .Y(n36798) );
  BUFX4 U25235 ( .A(n36794), .Y(n36799) );
  INVX12 U25236 ( .A(n42594), .Y(n42592) );
  INVX12 U25237 ( .A(net209615), .Y(net210479) );
  NAND4X4 U25238 ( .A(n44899), .B(n44898), .C(n44897), .D(n44896), .Y(
        net209615) );
  NAND4X4 U25239 ( .A(n45156), .B(n45155), .C(n45154), .D(n45153), .Y(n48312)
         );
  NOR4X2 U25240 ( .A(n45144), .B(n45143), .C(n45142), .D(n45141), .Y(n45155)
         );
  CLKINVX16 U25241 ( .A(n36864), .Y(n36865) );
  CLKINVX8 U25242 ( .A(n42593), .Y(n42590) );
  CLKBUFX2 U25243 ( .A(n42598), .Y(n42596) );
  CLKBUFX20 U25244 ( .A(n42611), .Y(n42605) );
  BUFX8 U25245 ( .A(n42611), .Y(n42604) );
  NOR2X6 U25246 ( .A(n44984), .B(n48307), .Y(n44994) );
  NAND2X2 U25247 ( .A(n48308), .B(n48307), .Y(n48311) );
  NAND4BX4 U25248 ( .AN(n41697), .B(n44983), .C(n44982), .D(n44981), .Y(n48307) );
  CLKINVX4 U25249 ( .A(n37017), .Y(n42629) );
  CLKINVX6 U25250 ( .A(n37017), .Y(n42628) );
  CLKINVX20 U25251 ( .A(n42634), .Y(n42633) );
  NAND4X4 U25252 ( .A(n45777), .B(n45776), .C(n45775), .D(n45774), .Y(n11084)
         );
  NOR2X1 U25253 ( .A(n12702), .B(n45773), .Y(n45777) );
  BUFX12 U25254 ( .A(n34435), .Y(n42717) );
  BUFX16 U25255 ( .A(n36924), .Y(n42679) );
  CLKINVX12 U25256 ( .A(n42678), .Y(n42671) );
  NAND4X4 U25257 ( .A(n46375), .B(n46374), .C(n46373), .D(n46372), .Y(
        net209311) );
  NOR2X2 U25258 ( .A(n46365), .B(n48137), .Y(n46375) );
  OAI2BB1X4 U25259 ( .A0N(n12073), .A1N(n41704), .B0(n12147), .Y(n48127) );
  NAND2X2 U25260 ( .A(n10559), .B(n12073), .Y(n48207) );
  NOR2X6 U25261 ( .A(n12073), .B(n46143), .Y(n46147) );
  NAND4X4 U25262 ( .A(n43577), .B(n43576), .C(n43575), .D(n43574), .Y(n12073)
         );
  AOI21X1 U25263 ( .A0(n48055), .A1(n10727), .B0(n37199), .Y(n48056) );
  NAND2XL U25264 ( .A(n10727), .B(n39892), .Y(n39646) );
  NAND2BX4 U25265 ( .AN(n39363), .B(net211473), .Y(n10727) );
  CLKINVX6 U25266 ( .A(n42556), .Y(n42548) );
  CLKBUFX20 U25267 ( .A(n42548), .Y(n36832) );
  CLKINVX20 U25268 ( .A(n42555), .Y(n42552) );
  BUFX12 U25269 ( .A(n34455), .Y(n42546) );
  NOR2X8 U25270 ( .A(n47325), .B(net209317), .Y(n47335) );
  NAND2XL U25271 ( .A(net209314), .B(net209317), .Y(n47780) );
  NAND4X6 U25272 ( .A(n46331), .B(n46330), .C(n46329), .D(n46328), .Y(
        net209317) );
  INVX12 U25273 ( .A(n41325), .Y(n36800) );
  CLKINVX20 U25274 ( .A(n36800), .Y(n36801) );
  INVX8 U25275 ( .A(n42626), .Y(n36802) );
  INVX1 U25276 ( .A(n42630), .Y(n36803) );
  INVXL U25277 ( .A(n42628), .Y(n36804) );
  INVXL U25278 ( .A(n42628), .Y(n36805) );
  INVX4 U25279 ( .A(n42635), .Y(n42626) );
  CLKINVX3 U25280 ( .A(n42635), .Y(n42625) );
  CLKINVX16 U25281 ( .A(n42634), .Y(n42632) );
  CLKINVX16 U25282 ( .A(n42634), .Y(n42630) );
  CLKINVX16 U25283 ( .A(n42634), .Y(n42631) );
  INVX3 U25284 ( .A(n42624), .Y(n42636) );
  NOR2X6 U25285 ( .A(n45733), .B(n48225), .Y(n45737) );
  OAI21X4 U25286 ( .A0(n49501), .A1(n48118), .B0(n48225), .Y(n48119) );
  NAND4X4 U25287 ( .A(n44525), .B(n44524), .C(n44523), .D(n44522), .Y(n48225)
         );
  NAND4X4 U25288 ( .A(n43558), .B(n43557), .C(n43556), .D(n43555), .Y(n11751)
         );
  NOR4X4 U25289 ( .A(n29432), .B(n29433), .C(n29434), .D(n29435), .Y(n43558)
         );
  NOR4X2 U25290 ( .A(n29436), .B(n29437), .C(n29438), .D(n29439), .Y(n43557)
         );
  INVX6 U25291 ( .A(n41306), .Y(n36806) );
  CLKBUFX8 U25292 ( .A(n36806), .Y(n36807) );
  BUFX16 U25293 ( .A(n36806), .Y(n36808) );
  BUFX16 U25294 ( .A(n36806), .Y(n36809) );
  BUFX12 U25295 ( .A(n36806), .Y(n36810) );
  BUFX12 U25296 ( .A(n36806), .Y(n36811) );
  BUFX4 U25297 ( .A(n34461), .Y(n36812) );
  BUFX8 U25298 ( .A(n36812), .Y(n36813) );
  CLKBUFX8 U25299 ( .A(n36812), .Y(n36814) );
  CLKBUFX8 U25300 ( .A(n36812), .Y(n36815) );
  CLKBUFX6 U25301 ( .A(n36812), .Y(n36816) );
  CLKBUFX6 U25302 ( .A(n36812), .Y(n36817) );
  CLKBUFX20 U25303 ( .A(n42700), .Y(n42696) );
  AND4XL U25304 ( .A(net209325), .B(net209317), .C(net209314), .D(net209316),
        .Y(n37468) );
  NAND2X4 U25305 ( .A(n37204), .B(n46342), .Y(net209314) );
  BUFX20 U25306 ( .A(n36910), .Y(n42585) );
  CLKINVX6 U25307 ( .A(n36910), .Y(n42576) );
  CLKINVX3 U25308 ( .A(n36910), .Y(n42583) );
  CLKINVX3 U25309 ( .A(n36910), .Y(n42580) );
  CLKINVX8 U25310 ( .A(n42604), .Y(n36818) );
  INVX20 U25311 ( .A(n36818), .Y(n36819) );
  BUFX8 U25312 ( .A(n41646), .Y(n42621) );
  INVX16 U25313 ( .A(n42622), .Y(n42615) );
  CLKINVX4 U25314 ( .A(n42726), .Y(n42723) );
  NOR2X6 U25315 ( .A(n44307), .B(net209519), .Y(net215231) );
  INVXL U25316 ( .A(net209519), .Y(net171255) );
  NAND2XL U25317 ( .A(n10369), .B(net209519), .Y(n39849) );
  AOI21XL U25318 ( .A0(net209519), .A1(net209520), .B0(net171249), .Y(n48367)
         );
  NAND4X4 U25319 ( .A(n44306), .B(n44305), .C(n44304), .D(n44303), .Y(
        net209519) );
  CLKINVX8 U25320 ( .A(net258261), .Y(net219330) );
  XOR2X1 U25321 ( .A(n41817), .B(n42610), .Y(n45438) );
  CLKBUFX12 U25322 ( .A(n42595), .Y(n42610) );
  NOR2X6 U25323 ( .A(n12798), .B(n45843), .Y(n45847) );
  NAND2XL U25324 ( .A(n12798), .B(n12017), .Y(n48235) );
  AOI21X2 U25325 ( .A0(n48242), .A1(n12798), .B0(net209791), .Y(n48243) );
  NAND3XL U25326 ( .A(n12692), .B(n12798), .C(n39291), .Y(n10532) );
  NAND4X4 U25327 ( .A(n43722), .B(n43721), .C(n43720), .D(n43719), .Y(n12798)
         );
  AOI21X4 U25328 ( .A0(n40902), .A1(n40903), .B0(n40904), .Y(n40901) );
  OAI21X2 U25329 ( .A0(n40898), .A1(n41007), .B0(n41009), .Y(n40903) );
  NAND2XL U25330 ( .A(n12915), .B(n11359), .Y(n48089) );
  NAND3XL U25331 ( .A(n11359), .B(n11358), .C(n11352), .Y(n10024) );
  NAND4X2 U25332 ( .A(n47072), .B(n47071), .C(n47070), .D(n47069), .Y(n11359)
         );
  CLKBUFX3 U25333 ( .A(n36920), .Y(n42509) );
  INVX6 U25334 ( .A(n42510), .Y(n42501) );
  AOI21X4 U25335 ( .A0(n40875), .A1(n40876), .B0(n40877), .Y(n40874) );
  OAI21X2 U25336 ( .A0(n40870), .A1(n41047), .B0(n41048), .Y(n40876) );
  INVX12 U25337 ( .A(n34454), .Y(n36820) );
  CLKINVX12 U25338 ( .A(n36820), .Y(n36821) );
  CLKINVX12 U25339 ( .A(n36820), .Y(n36822) );
  CLKINVX12 U25340 ( .A(n36820), .Y(n36823) );
  CLKINVX12 U25341 ( .A(n36820), .Y(n36824) );
  CLKINVX12 U25342 ( .A(n36820), .Y(n36825) );
  CLKINVX8 U25343 ( .A(n41334), .Y(n36826) );
  CLKBUFX20 U25344 ( .A(n36826), .Y(n36827) );
  CLKBUFX4 U25345 ( .A(n36826), .Y(n36828) );
  CLKBUFX4 U25346 ( .A(n36826), .Y(n36829) );
  CLKBUFX4 U25347 ( .A(n36826), .Y(n36830) );
  BUFX12 U25348 ( .A(n36826), .Y(n36831) );
  NOR4BBX4 U25349 ( .AN(n41732), .BN(n41733), .C(n45450), .D(n45449), .Y(
        n45451) );
  XOR2X1 U25350 ( .A(n34324), .B(n42690), .Y(n45449) );
  INVX8 U25351 ( .A(n42683), .Y(n36833) );
  CLKINVX16 U25352 ( .A(n36833), .Y(n36834) );
  NAND2XL U25353 ( .A(n48301), .B(n48309), .Y(net210660) );
  NOR2X4 U25354 ( .A(n45126), .B(n48309), .Y(n45136) );
  NAND4X4 U25355 ( .A(n45125), .B(n45124), .C(n45123), .D(n45122), .Y(n48309)
         );
  AOI21X2 U25356 ( .A0(n48124), .A1(n12144), .B0(net171191), .Y(n48125) );
  NOR2X6 U25357 ( .A(n12144), .B(n46123), .Y(n46127) );
  NAND3XL U25358 ( .A(n12145), .B(n12144), .C(n39300), .Y(n10564) );
  NAND4BBX4 U25359 ( .AN(n43624), .BN(n43623), .C(n43622), .D(n43621), .Y(
        n12144) );
  XNOR2X2 U25360 ( .A(n50559), .B(n42723), .Y(n29145) );
  OAI2BB1XL U25361 ( .A0N(n12746), .A1N(n41783), .B0(n12742), .Y(n48203) );
  NAND2X2 U25362 ( .A(n12085), .B(n12742), .Y(n48195) );
  NAND2XL U25363 ( .A(n12746), .B(n12742), .Y(n10570) );
  NOR2X4 U25364 ( .A(n12742), .B(n45694), .Y(net213342) );
  NAND4X4 U25365 ( .A(n44211), .B(n44210), .C(n44209), .D(n44208), .Y(n12742)
         );
  XNOR2X1 U25366 ( .A(n50772), .B(n36863), .Y(n29134) );
  OAI21X4 U25367 ( .A0(net171105), .A1(n48262), .B0(n40388), .Y(n48263) );
  AOI21X4 U25368 ( .A0(n48261), .A1(n11976), .B0(n39289), .Y(n48262) );
  BUFX6 U25369 ( .A(n42556), .Y(n42555) );
  XNOR2X1 U25370 ( .A(n51200), .B(n42629), .Y(n29133) );
  AOI21X4 U25371 ( .A0(n40879), .A1(n40880), .B0(n40881), .Y(n40878) );
  OAI21X2 U25372 ( .A0(n40874), .A1(n41049), .B0(n41050), .Y(n40880) );
  OAI21X4 U25373 ( .A0(n40888), .A1(n40991), .B0(n40997), .Y(n40891) );
  NOR2X2 U25374 ( .A(n40884), .B(n40889), .Y(n40888) );
  AOI21X4 U25375 ( .A0(n40839), .A1(n40840), .B0(n40841), .Y(n40838) );
  OAI21X2 U25376 ( .A0(n40834), .A1(n37517), .B0(n41100), .Y(n40840) );
  NOR4XL U25377 ( .A(n29135), .B(n29133), .C(n29132), .D(n29134), .Y(n44597)
         );
  XOR2X2 U25378 ( .A(n41867), .B(n42601), .Y(n29135) );
  OAI21X4 U25379 ( .A0(n40760), .A1(n40486), .B0(n11884), .Y(n40490) );
  OAI21X2 U25380 ( .A0(n40878), .A1(n41051), .B0(n41052), .Y(n41189) );
  AOI21X4 U25381 ( .A0(n40851), .A1(n40852), .B0(n40853), .Y(n40850) );
  OAI21X2 U25382 ( .A0(n40848), .A1(n41109), .B0(n41110), .Y(n40852) );
  INVX4 U25383 ( .A(n36835), .Y(n36836) );
  BUFX8 U25384 ( .A(n36836), .Y(n36837) );
  BUFX20 U25385 ( .A(n36836), .Y(n36838) );
  BUFX16 U25386 ( .A(n36836), .Y(n36839) );
  BUFX12 U25387 ( .A(n36836), .Y(n36840) );
  BUFX12 U25388 ( .A(n36836), .Y(n36841) );
  BUFX12 U25389 ( .A(n34460), .Y(n36842) );
  CLKBUFX16 U25390 ( .A(n36842), .Y(n36843) );
  CLKBUFX16 U25391 ( .A(n36842), .Y(n36844) );
  CLKBUFX16 U25392 ( .A(n36842), .Y(n36845) );
  CLKBUFX16 U25393 ( .A(n36842), .Y(n36846) );
  CLKBUFX16 U25394 ( .A(n36842), .Y(n36847) );
  INVX4 U25395 ( .A(n36848), .Y(n36849) );
  CLKBUFX12 U25396 ( .A(n36849), .Y(n36850) );
  CLKBUFX12 U25397 ( .A(n36849), .Y(n36851) );
  BUFX20 U25398 ( .A(n36849), .Y(n36852) );
  BUFX20 U25399 ( .A(n36849), .Y(n36853) );
  CLKBUFX12 U25400 ( .A(n36849), .Y(n36854) );
  BUFX8 U25401 ( .A(n34466), .Y(n36855) );
  BUFX20 U25402 ( .A(n36855), .Y(n36856) );
  BUFX20 U25403 ( .A(n36855), .Y(n36857) );
  BUFX20 U25404 ( .A(n36855), .Y(n36858) );
  BUFX20 U25405 ( .A(n36855), .Y(n36859) );
  BUFX20 U25406 ( .A(n36855), .Y(n36860) );
  NOR2XL U25407 ( .A(net210205), .B(net210216), .Y(n47663) );
  NOR2X6 U25408 ( .A(net210211), .B(net210216), .Y(n47760) );
  NOR3X4 U25409 ( .A(net209335), .B(n47662), .C(n47661), .Y(net210216) );
  OAI211X2 U25410 ( .A0(net209659), .A1(n11750), .B0(n11751), .C0(n11752), .Y(
        n11746) );
  NAND2X6 U25411 ( .A(n41366), .B(n11756), .Y(n11750) );
  OAI31X2 U25412 ( .A0(n12083), .A1(net171236), .A2(net209844), .B0(net151723),
        .Y(n12081) );
  NAND4X2 U25413 ( .A(net209333), .B(n47696), .C(n47695), .D(n47694), .Y(
        n47984) );
  CLKINVX12 U25414 ( .A(n42715), .Y(n41641) );
  CLKBUFX4 U25415 ( .A(n42716), .Y(n42715) );
  AOI21X2 U25416 ( .A0(n48298), .A1(net209604), .B0(net209633), .Y(n48299) );
  NAND4XL U25417 ( .A(net209604), .B(net209606), .C(net209636), .D(net210669),
        .Y(net210469) );
  NAND4X4 U25418 ( .A(n45511), .B(n45510), .C(n45509), .D(n45508), .Y(
        net209604) );
  CLKINVX8 U25419 ( .A(n42591), .Y(n36862) );
  NAND4X4 U25420 ( .A(n46433), .B(n46432), .C(n46431), .D(n46430), .Y(
        net209300) );
  NOR2X2 U25421 ( .A(n46423), .B(net209884), .Y(n46433) );
  INVX4 U25422 ( .A(n34448), .Y(n42623) );
  INVX8 U25423 ( .A(n41646), .Y(n41647) );
  NOR2X4 U25424 ( .A(n44873), .B(net209628), .Y(net214389) );
  NAND2XL U25425 ( .A(net209628), .B(net209603), .Y(n47740) );
  AND3XL U25426 ( .A(net209602), .B(net209631), .C(net209628), .Y(n37126) );
  NAND2X8 U25427 ( .A(n37197), .B(n44871), .Y(net209628) );
  INVX3 U25428 ( .A(n42635), .Y(n42627) );
  AOI21X4 U25429 ( .A0(n48252), .A1(n10157), .B0(net171136), .Y(n48253) );
  OAI21X4 U25430 ( .A0(net171132), .A1(n48251), .B0(n10525), .Y(n48252) );
  CLKBUFX4 U25431 ( .A(n42691), .Y(n42701) );
  CLKINVX8 U25432 ( .A(n42590), .Y(n36864) );
  INVX4 U25433 ( .A(n34443), .Y(n42688) );
  CLKINVX8 U25434 ( .A(n42685), .Y(n42684) );
  CLKBUFX2 U25435 ( .A(n34445), .Y(n42650) );
  BUFX12 U25436 ( .A(n34445), .Y(n42649) );
  CLKINVX12 U25437 ( .A(n36915), .Y(n36890) );
  NAND2X1 U25438 ( .A(n41876), .B(n36915), .Y(n41268) );
  INVX3 U25439 ( .A(n42640), .Y(n36866) );
  INVXL U25440 ( .A(n42645), .Y(n42640) );
  INVX1 U25441 ( .A(n41648), .Y(n41649) );
  BUFX16 U25442 ( .A(n41648), .Y(n42726) );
  INVX1 U25443 ( .A(n41648), .Y(n42718) );
  CLKINVX3 U25444 ( .A(n41648), .Y(n42719) );
  BUFX20 U25445 ( .A(n42511), .Y(n42529) );
  CLKBUFX2 U25446 ( .A(n42513), .Y(n42530) );
  CLKBUFX20 U25447 ( .A(n42529), .Y(n42519) );
  NOR4X2 U25448 ( .A(n45115), .B(n45114), .C(n45113), .D(n45112), .Y(n45124)
         );
  XOR2X1 U25449 ( .A(n34346), .B(n36907), .Y(n45114) );
  CLKBUFX20 U25450 ( .A(n42519), .Y(n42518) );
  CLKBUFX20 U25451 ( .A(n36877), .Y(n41322) );
  BUFX12 U25452 ( .A(n42596), .Y(n42611) );
  CLKINVX8 U25453 ( .A(n36909), .Y(n42707) );
  BUFX20 U25454 ( .A(n41647), .Y(n36868) );
  NAND3X4 U25455 ( .A(n36941), .B(n37238), .C(n39463), .Y(net210477) );
  NOR4X2 U25456 ( .A(n45085), .B(n45084), .C(n45083), .D(n45082), .Y(n37238)
         );
  CLKXOR2X1 U25457 ( .A(n34388), .B(n42637), .Y(n44884) );
  INVX4 U25458 ( .A(net219322), .Y(n36869) );
  CLKINVX12 U25459 ( .A(n36869), .Y(n36870) );
  INVX1 U25460 ( .A(net258261), .Y(net219322) );
  NOR2X6 U25461 ( .A(n10376), .B(n43564), .Y(n43568) );
  INVXL U25462 ( .A(n10376), .Y(net171185) );
  NAND3X6 U25463 ( .A(net216137), .B(n39455), .C(net216138), .Y(n10376) );
  OAI2BB1X4 U25464 ( .A0N(n48186), .A1N(n41781), .B0(n48132), .Y(n48135) );
  NAND3X2 U25465 ( .A(n48186), .B(net209862), .C(n48185), .Y(n48190) );
  CLKAND2X3 U25466 ( .A(n48186), .B(n48130), .Y(n36947) );
  NOR2X4 U25467 ( .A(n46200), .B(n48186), .Y(n46204) );
  NAND4X4 U25468 ( .A(n43885), .B(n43884), .C(n43883), .D(n43882), .Y(n48186)
         );
  BUFX20 U25469 ( .A(n41384), .Y(n36871) );
  BUFX20 U25470 ( .A(n42689), .Y(n42693) );
  CLKBUFX4 U25471 ( .A(n42692), .Y(n42689) );
  CLKBUFX2 U25472 ( .A(net258261), .Y(net219346) );
  CLKBUFX20 U25473 ( .A(net219330), .Y(n40039) );
  INVX8 U25474 ( .A(n41320), .Y(n36872) );
  CLKINVX20 U25475 ( .A(n36872), .Y(n36873) );
  CLKBUFX2 U25476 ( .A(n34453), .Y(n41320) );
  NOR2X6 U25477 ( .A(n10565), .B(n46113), .Y(n46117) );
  OAI21X1 U25478 ( .A0(net171188), .A1(n48125), .B0(n10565), .Y(n48126) );
  NAND2XL U25479 ( .A(n12736), .B(n10565), .Y(n39801) );
  NAND2BX4 U25480 ( .AN(n39299), .B(net216047), .Y(n10565) );
  CLKBUFX2 U25481 ( .A(n42688), .Y(n42686) );
  INVX12 U25482 ( .A(n36922), .Y(n41380) );
  INVX3 U25483 ( .A(n34442), .Y(net219492) );
  BUFX4 U25484 ( .A(n34442), .Y(net219494) );
  CLKBUFX2 U25485 ( .A(n42688), .Y(n42685) );
  INVXL U25486 ( .A(n10377), .Y(net151308) );
  NOR2X6 U25487 ( .A(n10377), .B(n43630), .Y(n43634) );
  AO21X4 U25488 ( .A0(n10377), .A1(net171189), .B0(net209661), .Y(n41381) );
  NAND4X4 U25489 ( .A(net216043), .B(net216044), .C(net216045), .D(net216046),
        .Y(n10377) );
  CLKBUFX2 U25490 ( .A(net219472), .Y(net219478) );
  XNOR2X1 U25491 ( .A(n41811), .B(n42526), .Y(n44936) );
  XNOR2X1 U25492 ( .A(n41809), .B(n42526), .Y(n45104) );
  CLKBUFX20 U25493 ( .A(n42526), .Y(n42515) );
  XOR2X1 U25494 ( .A(n41843), .B(n42526), .Y(n27712) );
  XOR2X1 U25495 ( .A(n42526), .B(n41840), .Y(n44029) );
  BUFX20 U25496 ( .A(n42527), .Y(n42526) );
  INVX8 U25497 ( .A(net219494), .Y(net219484) );
  INVX16 U25498 ( .A(net219472), .Y(net219468) );
  CLKINVX20 U25499 ( .A(net219484), .Y(net219434) );
  BUFX6 U25500 ( .A(n36920), .Y(n42510) );
  CLKBUFX4 U25501 ( .A(n42598), .Y(n42597) );
  BUFX4 U25502 ( .A(n34449), .Y(n42599) );
  CLKXOR2X2 U25503 ( .A(n41866), .B(n42601), .Y(n29165) );
  CLKBUFX4 U25504 ( .A(n42612), .Y(n42601) );
  INVX3 U25505 ( .A(n41649), .Y(n36874) );
  CLKINVX12 U25506 ( .A(n36874), .Y(n36875) );
  CLKBUFX20 U25507 ( .A(n34439), .Y(n41283) );
  CLKBUFX16 U25508 ( .A(n34439), .Y(n41281) );
  CLKBUFX12 U25509 ( .A(n34439), .Y(n41282) );
  BUFX20 U25510 ( .A(n34444), .Y(n42669) );
  XOR2X1 U25511 ( .A(n34386), .B(n34444), .Y(n44886) );
  XOR2X1 U25512 ( .A(n34146), .B(n34444), .Y(n43985) );
  XOR2X1 U25513 ( .A(n34290), .B(n34444), .Y(n45384) );
  XOR2X1 U25514 ( .A(n34210), .B(n34444), .Y(n44739) );
  NAND2X1 U25515 ( .A(n41217), .B(n34444), .Y(n41220) );
  CLKBUFX6 U25516 ( .A(n42623), .Y(n42622) );
  BUFX20 U25517 ( .A(n42636), .Y(n42634) );
  BUFX16 U25518 ( .A(n37017), .Y(n42635) );
  BUFX20 U25519 ( .A(n34447), .Y(n42624) );
  CLKBUFX20 U25520 ( .A(n42664), .Y(n42652) );
  BUFX12 U25521 ( .A(n42646), .Y(n42664) );
  OAI21X4 U25522 ( .A0(n47718), .A1(net210688), .B0(net234529), .Y(n47720) );
  AOI21X4 U25523 ( .A0(net210690), .A1(n47717), .B0(n47716), .Y(n47718) );
  XOR2X1 U25524 ( .A(n34400), .B(net219434), .Y(n44888) );
  BUFX8 U25525 ( .A(n36921), .Y(n42594) );
  CLKBUFX20 U25526 ( .A(n41385), .Y(n42697) );
  CLKBUFX12 U25527 ( .A(n34456), .Y(n42532) );
  INVX20 U25528 ( .A(n42532), .Y(n42545) );
  BUFX20 U25529 ( .A(n42703), .Y(n41385) );
  CLKBUFX20 U25530 ( .A(n42699), .Y(n42698) );
  CLKBUFX6 U25531 ( .A(n42689), .Y(n42699) );
  NAND4X6 U25532 ( .A(n44039), .B(n44038), .C(n44037), .D(n44036), .Y(
        net209862) );
  NOR2X6 U25533 ( .A(n44029), .B(n48336), .Y(n44039) );
  CLKINVX3 U25534 ( .A(n41629), .Y(n41630) );
  CLKBUFX2 U25535 ( .A(n41629), .Y(n42573) );
  XNOR2X2 U25536 ( .A(n50355), .B(n42671), .Y(n29166) );
  AOI211X2 U25537 ( .A0(net151479), .A1(n11336), .B0(net151481), .C0(n39908),
        .Y(n11332) );
  OAI31X2 U25538 ( .A0(n11339), .A1(net151467), .A2(net151465), .B0(n10015),
        .Y(n11336) );
  INVX6 U25539 ( .A(n41324), .Y(n36876) );
  CLKINVX20 U25540 ( .A(n36876), .Y(n36877) );
  CLKBUFX2 U25541 ( .A(n34453), .Y(n41324) );
  BUFX20 U25542 ( .A(n41380), .Y(n41319) );
  XNOR2XL U25543 ( .A(n50394), .B(n41380), .Y(n26218) );
  XNOR2XL U25544 ( .A(n50385), .B(n41380), .Y(n26429) );
  CLKBUFX12 U25545 ( .A(n42523), .Y(n42524) );
  CLKBUFX4 U25546 ( .A(n42512), .Y(n42523) );
  CLKBUFX2 U25547 ( .A(n34438), .Y(n42703) );
  CLKBUFX20 U25548 ( .A(n42607), .Y(n42608) );
  CLKINVX12 U25549 ( .A(n42545), .Y(n42537) );
  CLKBUFX20 U25550 ( .A(n42530), .Y(n42522) );
  XOR2X1 U25551 ( .A(n41818), .B(n42609), .Y(n45467) );
  CLKBUFX6 U25552 ( .A(n42595), .Y(n42609) );
  CLKINVX8 U25553 ( .A(n41335), .Y(n36878) );
  BUFX20 U25554 ( .A(n36878), .Y(n36879) );
  BUFX20 U25555 ( .A(n36878), .Y(n36880) );
  BUFX20 U25556 ( .A(n36878), .Y(n36881) );
  BUFX20 U25557 ( .A(n36878), .Y(n36882) );
  BUFX20 U25558 ( .A(n36878), .Y(n36883) );
  INVX6 U25559 ( .A(n34437), .Y(n36884) );
  INVX12 U25560 ( .A(n36884), .Y(n36885) );
  CLKINVX12 U25561 ( .A(n36884), .Y(n36886) );
  CLKINVX8 U25562 ( .A(n36884), .Y(n36887) );
  CLKINVX8 U25563 ( .A(n36884), .Y(n36888) );
  CLKINVX8 U25564 ( .A(n36884), .Y(n36889) );
  BUFX12 U25565 ( .A(n36909), .Y(n42714) );
  BUFX6 U25566 ( .A(n36909), .Y(n42713) );
  BUFX8 U25567 ( .A(net219492), .Y(net219472) );
  INVX8 U25568 ( .A(net210524), .Y(net210210) );
  NAND2X2 U25569 ( .A(net210526), .B(net210524), .Y(n47762) );
  NAND4X6 U25570 ( .A(n47644), .B(n47643), .C(n47642), .D(n47641), .Y(
        net210524) );
  NOR2X4 U25571 ( .A(n12086), .B(n45680), .Y(n45684) );
  INVX8 U25572 ( .A(n12086), .Y(net209846) );
  NAND4BXL U25573 ( .AN(net171234), .B(n12087), .C(n12089), .D(n12086), .Y(
        n39315) );
  AOI31X2 U25574 ( .A0(n12086), .A1(n12087), .A2(n12088), .B0(n10577), .Y(
        n12083) );
  NAND3X6 U25575 ( .A(n45679), .B(n45678), .C(net209638), .Y(n12086) );
  BUFX20 U25576 ( .A(n42605), .Y(n42602) );
  BUFX16 U25577 ( .A(n36890), .Y(n36891) );
  BUFX20 U25578 ( .A(n36890), .Y(n36892) );
  BUFX16 U25579 ( .A(n36890), .Y(n36893) );
  CLKBUFX12 U25580 ( .A(n36890), .Y(n36894) );
  BUFX12 U25581 ( .A(n36890), .Y(n36895) );
  BUFX12 U25582 ( .A(n34441), .Y(n36896) );
  CLKBUFX16 U25583 ( .A(n36896), .Y(n36897) );
  CLKBUFX16 U25584 ( .A(n36896), .Y(n36898) );
  CLKBUFX16 U25585 ( .A(n36896), .Y(n36899) );
  CLKBUFX16 U25586 ( .A(n36896), .Y(n36900) );
  CLKBUFX16 U25587 ( .A(n36896), .Y(n36901) );
  CLKBUFX12 U25588 ( .A(n42690), .Y(n42700) );
  INVX12 U25589 ( .A(n42546), .Y(n42556) );
  INVX12 U25590 ( .A(net258262), .Y(net219356) );
  XOR2X1 U25591 ( .A(n34334), .B(net258262), .Y(n45427) );
  XNOR2X2 U25592 ( .A(n50970), .B(net258262), .Y(n26853) );
  XNOR2X2 U25593 ( .A(n50984), .B(net258262), .Y(n29260) );
  XNOR2X4 U25594 ( .A(n50943), .B(net258262), .Y(n24810) );
  BUFX12 U25595 ( .A(n41286), .Y(n42656) );
  CLKINVX8 U25596 ( .A(n41285), .Y(n41286) );
  INVX8 U25597 ( .A(n42684), .Y(n36902) );
  CLKINVX20 U25598 ( .A(n36902), .Y(n36903) );
  NOR2X6 U25599 ( .A(n10368), .B(n44308), .Y(net215222) );
  BUFX20 U25600 ( .A(n42665), .Y(n42655) );
  CLKBUFX6 U25601 ( .A(n42646), .Y(n42665) );
  CLKINVX8 U25602 ( .A(n42645), .Y(n42638) );
  CLKINVX3 U25603 ( .A(n42645), .Y(n42642) );
  CLKINVX3 U25604 ( .A(n42645), .Y(n42644) );
  BUFX12 U25605 ( .A(n36912), .Y(n42645) );
  CLKXOR2X2 U25606 ( .A(n34385), .B(n41380), .Y(n44887) );
  INVX12 U25607 ( .A(n42681), .Y(n36904) );
  CLKINVX20 U25608 ( .A(n36904), .Y(n36905) );
  NAND2XL U25609 ( .A(net210677), .B(net209862), .Y(n39306) );
  NOR2BXL U25610 ( .AN(net209862), .B(net209944), .Y(n47725) );
  NOR2XL U25611 ( .A(n46210), .B(net209862), .Y(n46220) );
  AO21X4 U25612 ( .A0(net209944), .A1(net209862), .B0(n48131), .Y(n41781) );
  INVX6 U25613 ( .A(n42676), .Y(n36906) );
  CLKINVX16 U25614 ( .A(n36906), .Y(n36907) );
  NAND2XL U25615 ( .A(n33800), .B(n36921), .Y(n41263) );
  BUFX8 U25616 ( .A(n42597), .Y(n42612) );
  BUFX16 U25617 ( .A(n42664), .Y(n42661) );
  BUFX20 U25618 ( .A(n42610), .Y(n42607) );
  OAI21XL U25619 ( .A0(n11762), .A1(net209537), .B0(n12538), .Y(n48358) );
  NAND2BX4 U25620 ( .AN(n11762), .B(n41682), .Y(n12079) );
  NAND4BX2 U25621 ( .AN(n41669), .B(n43589), .C(n43588), .D(n43587), .Y(n11762) );
  CLKINVX3 U25622 ( .A(net219356), .Y(net219308) );
  INVX1 U25623 ( .A(n36868), .Y(n41656) );
  INVX1 U25624 ( .A(n42623), .Y(n42614) );
  BUFX20 U25625 ( .A(n42702), .Y(n42695) );
  CLKBUFX8 U25626 ( .A(n42691), .Y(n42702) );
  OAI21X4 U25627 ( .A0(n40854), .A1(n41117), .B0(n41120), .Y(n41190) );
  AOI21X4 U25628 ( .A0(n40855), .A1(n40856), .B0(n40857), .Y(n40854) );
  CLKINVX12 U25629 ( .A(n42687), .Y(n41379) );
  CLKBUFX2 U25630 ( .A(n42688), .Y(n42687) );
  INVX1 U25631 ( .A(net209635), .Y(net210667) );
  NOR2X2 U25632 ( .A(n41375), .B(net171188), .Y(n12070) );
  OAI21XL U25633 ( .A0(net210205), .A1(n47988), .B0(net210207), .Y(n47993) );
  OAI211X1 U25634 ( .A0(n11719), .A1(n11720), .B0(n11721), .C0(n11722), .Y(
        n11714) );
  NOR3X1 U25635 ( .A(n41031), .B(n40919), .C(n40917), .Y(n40861) );
  NAND4X1 U25636 ( .A(n40418), .B(n40422), .C(n41032), .D(n41033), .Y(n40863)
         );
  NAND2X1 U25637 ( .A(n41030), .B(n41193), .Y(n40862) );
  NAND2X1 U25638 ( .A(n11524), .B(n11525), .Y(n41102) );
  NOR4X1 U25639 ( .A(net171528), .B(n_cell_303546_net277636), .C(net151562),
        .D(n39929), .Y(n41103) );
  NAND2X1 U25640 ( .A(net260299), .B(net260295), .Y(n40897) );
  NOR2X1 U25641 ( .A(n_cell_301249_net269596), .B(n39835), .Y(n40895) );
  NAND2X1 U25642 ( .A(n41004), .B(n41195), .Y(n40896) );
  AOI21X1 U25643 ( .A0(n39833), .A1(net271996), .B0(n40736), .Y(n40737) );
  NAND3BX1 U25644 ( .AN(net171180), .B(n12168), .C(n40735), .Y(n40734) );
  NOR2X1 U25645 ( .A(n40470), .B(n40475), .Y(n40474) );
  NAND2XL U25646 ( .A(net209320), .B(net209323), .Y(n47778) );
  NOR2X6 U25647 ( .A(n47777), .B(net210579), .Y(n47779) );
  AND2X2 U25648 ( .A(n41633), .B(n41373), .Y(n47777) );
  NOR2X4 U25649 ( .A(net209584), .B(net209592), .Y(n47743) );
  OAI2BB1XL U25650 ( .A0N(n10378), .A1N(n41381), .B0(n10376), .Y(n48282) );
  INVXL U25651 ( .A(n10378), .Y(net171192) );
  AOI211X1 U25652 ( .A0(net151733), .A1(n12081), .B0(net171242), .C0(net171240), .Y(n12076) );
  NAND2XL U25653 ( .A(n12064), .B(n12065), .Y(n12061) );
  INVXL U25654 ( .A(n48032), .Y(n48033) );
  NAND2X1 U25655 ( .A(net209903), .B(net209902), .Y(net210492) );
  AOI211X1 U25656 ( .A0(n11701), .A1(n11702), .B0(net151333), .C0(net151330),
        .Y(n11695) );
  NOR2X4 U25657 ( .A(n10257), .B(n47281), .Y(n47285) );
  NOR2X4 U25658 ( .A(n47623), .B(n48435), .Y(n47633) );
  NOR2X4 U25659 ( .A(n47579), .B(n48449), .Y(n47589) );
  NOR2XL U25660 ( .A(n10585), .B(n47007), .Y(n47011) );
  OAI211X1 U25661 ( .A0(net171524), .A1(n11281), .B0(n12858), .C0(n12856), .Y(
        n40694) );
  NOR2X1 U25662 ( .A(n40696), .B(net151539), .Y(n40697) );
  CLKBUFX3 U25663 ( .A(n42498), .Y(n42494) );
  CLKINVX4 U25664 ( .A(net212214), .Y(net209923) );
  NAND2X1 U25665 ( .A(n10966), .B(n10965), .Y(n41163) );
  NOR2X1 U25666 ( .A(net171406), .B(net171408), .Y(n41164) );
  NAND4X1 U25667 ( .A(n11585), .B(net259626), .C(net261422), .D(n11586), .Y(
        n41037) );
  AOI211X1 U25668 ( .A0(n41038), .A1(n11584), .B0(n41039), .C0(
        n_cell_301249_net269638), .Y(n41040) );
  NOR2X4 U25669 ( .A(n40865), .B(n40860), .Y(n40864) );
  BUFX3 U25670 ( .A(n42477), .Y(n42498) );
  NAND3X1 U25671 ( .A(n41106), .B(net260461), .C(n39341), .Y(n40847) );
  NOR2X1 U25672 ( .A(net151790), .B(n_cell_301249_net269740), .Y(n41106) );
  NOR2X1 U25673 ( .A(n40744), .B(n40480), .Y(n40745) );
  NAND2X1 U25674 ( .A(net272583), .B(n40742), .Y(n40743) );
  NOR3BXL U25675 ( .AN(n40668), .B(n_cell_301249_net269836), .C(n39481), .Y(
        n40667) );
  NAND2X1 U25676 ( .A(n_cell_303546_net278017), .B(n10947), .Y(n40668) );
  NAND2X1 U25677 ( .A(n11894), .B(n11893), .Y(n41012) );
  NOR2X1 U25678 ( .A(net171272), .B(net171274), .Y(n41013) );
  AOI21X1 U25679 ( .A0(n40711), .A1(n12834), .B0(n40712), .Y(n40533) );
  OAI21XL U25680 ( .A0(n_cell_303546_net277814), .A1(n10635), .B0(n40715), .Y(
        n40534) );
  NAND3XL U25681 ( .A(net210580), .B(net209335), .C(net210581), .Y(n41633) );
  INVX3 U25682 ( .A(net210213), .Y(net210616) );
  INVX1 U25683 ( .A(net210660), .Y(net210659) );
  INVX1 U25684 ( .A(n11442), .Y(net151708) );
  INVX1 U25685 ( .A(net209296), .Y(net209289) );
  NAND2X2 U25686 ( .A(n41386), .B(n11139), .Y(n11134) );
  NAND2XL U25687 ( .A(n11140), .B(n10879), .Y(n11137) );
  NOR2X2 U25688 ( .A(n41203), .B(n48157), .Y(n48165) );
  NOR2X2 U25689 ( .A(n37221), .B(n41202), .Y(n41203) );
  NAND2X2 U25690 ( .A(n12087), .B(net209846), .Y(n48201) );
  AOI21X1 U25691 ( .A0(n48481), .A1(n11138), .B0(net209258), .Y(n48482) );
  AOI21X1 U25692 ( .A0(n48429), .A1(n48467), .B0(net209350), .Y(n48430) );
  INVXL U25693 ( .A(n11149), .Y(net209347) );
  INVXL U25694 ( .A(n10257), .Y(net209350) );
  AOI21XL U25695 ( .A0(n48415), .A1(n11094), .B0(net171447), .Y(n48416) );
  AOI21X1 U25696 ( .A0(n48413), .A1(n12303), .B0(net171445), .Y(n48414) );
  OAI21X1 U25697 ( .A0(n10843), .A1(net209372), .B0(n12306), .Y(n48413) );
  NAND2XL U25698 ( .A(n11116), .B(n11117), .Y(n11113) );
  INVX1 U25699 ( .A(n12717), .Y(n48223) );
  AOI21X1 U25700 ( .A0(n48497), .A1(n48496), .B0(n48495), .Y(n48509) );
  NAND2XL U25701 ( .A(n41210), .B(n11072), .Y(n48519) );
  OAI211X1 U25702 ( .A0(n11100), .A1(n11101), .B0(n10843), .C0(n10846), .Y(
        n11097) );
  NOR2X1 U25703 ( .A(n48026), .B(n48025), .Y(n48045) );
  OAI211X1 U25704 ( .A0(n11707), .A1(n11708), .B0(n11709), .C0(n11710), .Y(
        n11702) );
  NAND2X1 U25705 ( .A(n48062), .B(n11410), .Y(n47968) );
  CLKINVX1 U25706 ( .A(n10231), .Y(net209185) );
  OAI211X1 U25707 ( .A0(n11080), .A1(n11081), .B0(n11082), .C0(n11083), .Y(
        n11077) );
  NAND3X4 U25708 ( .A(n40394), .B(n11369), .C(n11370), .Y(n11367) );
  AOI21X2 U25709 ( .A0(n48265), .A1(n11967), .B0(net209749), .Y(n48266) );
  CLKINVX1 U25710 ( .A(n12453), .Y(net209455) );
  NAND2X1 U25711 ( .A(n11639), .B(n11640), .Y(n11636) );
  NOR4X1 U25712 ( .A(n44657), .B(n44656), .C(n44655), .D(n44654), .Y(n44658)
         );
  NAND2X1 U25713 ( .A(n41205), .B(n42530), .Y(n41207) );
  XOR2X1 U25714 ( .A(n42059), .B(n42575), .Y(n45049) );
  XOR2X1 U25715 ( .A(n41806), .B(n42522), .Y(n45046) );
  NAND2X2 U25716 ( .A(n41277), .B(n41278), .Y(n41710) );
  NAND2XL U25717 ( .A(n37201), .B(n41322), .Y(n41278) );
  XOR2X1 U25718 ( .A(n41803), .B(n42533), .Y(n45047) );
  NOR2X2 U25719 ( .A(n46401), .B(n48175), .Y(n46411) );
  NOR3BXL U25720 ( .AN(n41085), .B(n_cell_301249_net269701), .C(
        n_cell_303546_net277772), .Y(n41087) );
  NAND2X1 U25721 ( .A(n10662), .B(n41080), .Y(n41081) );
  CLKINVX3 U25722 ( .A(net209316), .Y(net210583) );
  NOR2X2 U25723 ( .A(n47358), .B(net209343), .Y(n47368) );
  AOI21X1 U25724 ( .A0(n39605), .A1(n_cell_303546_net275967), .B0(n40727), .Y(
        n40728) );
  OAI21XL U25725 ( .A0(n12640), .A1(n_cell_301249_net269568), .B0(n40724), .Y(
        n40725) );
  NOR2X4 U25726 ( .A(net209732), .B(n40468), .Y(n40467) );
  NAND2X1 U25727 ( .A(n_cell_303546_net275956), .B(n12867), .Y(n40687) );
  NOR2X1 U25728 ( .A(n40689), .B(n40517), .Y(n40690) );
  NOR2X2 U25729 ( .A(n47590), .B(net209323), .Y(n47600) );
  CLKINVX3 U25730 ( .A(net213680), .Y(net209622) );
  NAND4X2 U25731 ( .A(n44994), .B(n44993), .C(n44992), .D(n44991), .Y(n48149)
         );
  NOR4X1 U25732 ( .A(n43982), .B(n43981), .C(n43980), .D(n43979), .Y(n43998)
         );
  NAND4X2 U25733 ( .A(n46505), .B(n46504), .C(n46503), .D(n46502), .Y(n46510)
         );
  NAND4X4 U25734 ( .A(n46521), .B(n46520), .C(n46519), .D(n46518), .Y(n48449)
         );
  NAND4X2 U25735 ( .A(n46532), .B(n46531), .C(n46530), .D(n46529), .Y(n48446)
         );
  INVX4 U25736 ( .A(n46595), .Y(n48142) );
  NOR2X2 U25737 ( .A(n39304), .B(n46997), .Y(n47001) );
  XOR2XL U25738 ( .A(n9668), .B(n41281), .Y(n45247) );
  NOR3X1 U25739 ( .A(n40625), .B(net151374), .C(n40580), .Y(n40626) );
  NOR2BX1 U25740 ( .AN(n_cell_303546_net276365), .B(net259665), .Y(n40580) );
  NAND3X1 U25741 ( .A(net212131), .B(net212130), .C(net212132), .Y(
        n_cell_301249_net267409) );
  CLKBUFX3 U25742 ( .A(n12851), .Y(net260474) );
  NOR2X1 U25743 ( .A(n37378), .B(n41097), .Y(n40797) );
  NAND2X1 U25744 ( .A(net212126), .B(net212125), .Y(n41097) );
  NAND2X6 U25745 ( .A(n37208), .B(n43841), .Y(n48187) );
  NOR2X1 U25746 ( .A(n28014), .B(n28013), .Y(n43822) );
  NAND4X4 U25747 ( .A(n43833), .B(n43832), .C(n43831), .D(n43830), .Y(n48133)
         );
  NOR4X1 U25748 ( .A(n26838), .B(n26837), .C(n26836), .D(n26835), .Y(net215216) );
  NOR2X2 U25749 ( .A(n36984), .B(n37261), .Y(n39468) );
  NAND2X1 U25750 ( .A(n39808), .B(net214882), .Y(n39293) );
  NOR2X2 U25751 ( .A(n37106), .B(n37309), .Y(n39808) );
  NOR2X1 U25752 ( .A(n36981), .B(n37215), .Y(n39458) );
  NOR4X1 U25753 ( .A(n29226), .B(n29227), .C(n29228), .D(n29229), .Y(n43580)
         );
  NOR4X2 U25754 ( .A(n28114), .B(n28115), .C(n28116), .D(n28117), .Y(n43807)
         );
  NOR4X2 U25755 ( .A(n28452), .B(n28453), .C(n28454), .D(n28455), .Y(n43714)
         );
  XOR2X1 U25756 ( .A(n41879), .B(n36892), .Y(n26796) );
  NAND2BX1 U25757 ( .AN(n40412), .B(n_cell_301249_net267429), .Y(n11601) );
  NAND2X1 U25758 ( .A(net216300), .B(net216299), .Y(n40412) );
  NOR2X1 U25759 ( .A(n36992), .B(n37296), .Y(n_cell_301249_net267429) );
  CLKINVX4 U25760 ( .A(net210553), .Y(net210749) );
  NAND4X2 U25761 ( .A(n43263), .B(n43262), .C(n43261), .D(n43260), .Y(n12005)
         );
  NOR2X2 U25762 ( .A(n11849), .B(n43664), .Y(n43668) );
  NOR2X2 U25763 ( .A(n11700), .B(n43773), .Y(n43777) );
  NAND2BX1 U25764 ( .AN(n_cell_301249_net267526), .B(net216211), .Y(
        n_cell_303546_net276178) );
  NAND2X1 U25765 ( .A(n40962), .B(net216212), .Y(n_cell_301249_net267526) );
  NAND2BX1 U25766 ( .AN(n_cell_301249_net267451), .B(net216301), .Y(n11935) );
  NAND3X1 U25767 ( .A(net216303), .B(net216302), .C(net216304), .Y(
        n_cell_301249_net267451) );
  NAND3X1 U25768 ( .A(net216434), .B(net216435), .C(n40793), .Y(n11614) );
  NOR2X1 U25769 ( .A(n36972), .B(n37281), .Y(n40793) );
  NAND3X1 U25770 ( .A(n12840), .B(n39342), .C(n40706), .Y(n40705) );
  NOR2X1 U25771 ( .A(n40707), .B(n40578), .Y(n40708) );
  NAND2BX1 U25772 ( .AN(n40441), .B(net213587), .Y(n12194) );
  NAND2X1 U25773 ( .A(n40636), .B(net213590), .Y(n40441) );
  NOR2X1 U25774 ( .A(n37166), .B(n37499), .Y(n40636) );
  NAND4X2 U25775 ( .A(n43572), .B(n43571), .C(n43570), .D(n43569), .Y(n11756)
         );
  CLKINVX1 U25776 ( .A(n11335), .Y(net151444) );
  NAND2BX1 U25777 ( .AN(n_cell_303546_net275906), .B(n_cell_301249_net267089),
        .Y(n39444) );
  NAND2X1 U25778 ( .A(net216397), .B(net216396), .Y(n_cell_303546_net275906)
         );
  NOR2X1 U25779 ( .A(n36965), .B(n37274), .Y(n_cell_301249_net267089) );
  NAND2X1 U25780 ( .A(n37341), .B(net215069), .Y(n11907) );
  NAND2X1 U25781 ( .A(n41173), .B(net213616), .Y(n_cell_301249_net267828) );
  NAND2X1 U25782 ( .A(n41129), .B(net213490), .Y(n_cell_301249_net267628) );
  NOR2X1 U25783 ( .A(n37025), .B(n37464), .Y(n41129) );
  NAND2BX1 U25784 ( .AN(n40426), .B(net213502), .Y(n12207) );
  NAND2X1 U25785 ( .A(n40663), .B(net213505), .Y(n40426) );
  NAND2X1 U25786 ( .A(n40595), .B(net213480), .Y(n40417) );
  NOR2X1 U25787 ( .A(n37039), .B(n37449), .Y(n40595) );
  NAND2BX1 U25788 ( .AN(n_cell_301249_net267754), .B(net216175), .Y(n11916) );
  NAND2X1 U25789 ( .A(n40957), .B(net216176), .Y(n_cell_301249_net267754) );
  NAND2X1 U25790 ( .A(net260277), .B(n39598), .Y(n39597) );
  NOR2X1 U25791 ( .A(n39823), .B(n39596), .Y(n39598) );
  CLKINVX1 U25792 ( .A(n11967), .Y(n39596) );
  NAND2X1 U25793 ( .A(n11969), .B(n11968), .Y(n39823) );
  CLKBUFX3 U25794 ( .A(net214677), .Y(net261422) );
  NAND2BX1 U25795 ( .AN(n_cell_301249_net267613), .B(net216229), .Y(n11925) );
  NAND2X1 U25796 ( .A(n40960), .B(net216230), .Y(n_cell_301249_net267613) );
  NAND2BX1 U25797 ( .AN(n_cell_301249_net267466), .B(net213467), .Y(n10960) );
  NAND2X1 U25798 ( .A(n41130), .B(net213469), .Y(n_cell_301249_net267466) );
  NAND2BX1 U25799 ( .AN(n_cell_301249_net267556), .B(net213472), .Y(n10958) );
  NAND2BX1 U25800 ( .AN(n41166), .B(net213475), .Y(n_cell_301249_net267556) );
  NAND2X1 U25801 ( .A(net213474), .B(net213473), .Y(n41166) );
  NAND2X1 U25802 ( .A(n41165), .B(net213464), .Y(n_cell_301249_net267562) );
  CLKBUFX3 U25803 ( .A(net211568), .Y(net261069) );
  CLKINVX1 U25804 ( .A(n11555), .Y(n_cell_303546_net277496) );
  CLKINVX1 U25805 ( .A(n11558), .Y(n_cell_303546_net277494) );
  NAND2BX1 U25806 ( .AN(n40458), .B(net213317), .Y(net209087) );
  NAND2X1 U25807 ( .A(n40598), .B(net213320), .Y(n40458) );
  CLKBUFX3 U25808 ( .A(n12183), .Y(net260302) );
  NAND3X1 U25809 ( .A(n11241), .B(n11242), .C(n39340), .Y(n10621) );
  NOR2X1 U25810 ( .A(n39619), .B(n39620), .Y(n39340) );
  CLKINVX1 U25811 ( .A(n12821), .Y(n39620) );
  CLKBUFX3 U25812 ( .A(n12403), .Y(net260346) );
  NAND2BX1 U25813 ( .AN(n_cell_301249_net268272), .B(net215141), .Y(n11883) );
  NAND2X1 U25814 ( .A(n41014), .B(net215144), .Y(n_cell_301249_net268272) );
  NOR2BX1 U25815 ( .AN(net215143), .B(n37362), .Y(n41014) );
  NAND2X1 U25816 ( .A(n12611), .B(n12614), .Y(n11904) );
  NAND3X1 U25817 ( .A(n39282), .B(n11907), .C(net260403), .Y(n10456) );
  NOR2X1 U25818 ( .A(n_cell_303546_net277854), .B(n39550), .Y(n39282) );
  NAND2BX1 U25819 ( .AN(n40444), .B(net214952), .Y(n11896) );
  NAND2X1 U25820 ( .A(net214955), .B(n_cell_301249_net268065), .Y(n40444) );
  NOR2X1 U25821 ( .A(n37127), .B(n37424), .Y(n_cell_301249_net268065) );
  NAND3X1 U25822 ( .A(net214973), .B(n_cell_301249_net268136), .C(net214970),
        .Y(n11894) );
  NOR2X1 U25823 ( .A(n37021), .B(n37423), .Y(n_cell_301249_net268136) );
  NAND3X1 U25824 ( .A(net214964), .B(n_cell_301249_net268071), .C(net214961),
        .Y(n11895) );
  AND2X2 U25825 ( .A(net214963), .B(net214962), .Y(n_cell_301249_net268071) );
  CLKBUFX3 U25826 ( .A(net211584), .Y(net272417) );
  NAND2X1 U25827 ( .A(n41174), .B(net213606), .Y(n_cell_301249_net267822) );
  NOR2X1 U25828 ( .A(n37086), .B(n37502), .Y(n41174) );
  NAND2X1 U25829 ( .A(n_cell_301249_net267763), .B(net213597), .Y(n10941) );
  NOR2X1 U25830 ( .A(n37377), .B(n41125), .Y(n_cell_301249_net267763) );
  NAND2X1 U25831 ( .A(net213599), .B(net213598), .Y(n41125) );
  CLKINVX1 U25832 ( .A(n12602), .Y(net151788) );
  NAND2X1 U25833 ( .A(n40951), .B(net212555), .Y(n_cell_301249_net268336) );
  AND2X2 U25834 ( .A(net212554), .B(net212553), .Y(n40951) );
  NOR2X1 U25835 ( .A(n_cell_301249_net269755), .B(n39935), .Y(n41116) );
  NAND2X1 U25836 ( .A(n11241), .B(n11242), .Y(n41115) );
  CLKBUFX3 U25837 ( .A(n12592), .Y(net260384) );
  CLKINVX3 U25838 ( .A(n41752), .Y(n41364) );
  NAND2X1 U25839 ( .A(net209300), .B(net209298), .Y(n47786) );
  OR2X6 U25840 ( .A(n47775), .B(n47774), .Y(n41357) );
  CLKINVX3 U25841 ( .A(net210598), .Y(net210597) );
  CLKINVX1 U25842 ( .A(n47772), .Y(n47773) );
  CLKINVX2 U25843 ( .A(net210650), .Y(net209591) );
  INVX1 U25844 ( .A(net210670), .Y(net209584) );
  INVXL U25845 ( .A(net209628), .Y(net209627) );
  AOI21X1 U25846 ( .A0(net209582), .A1(net209583), .B0(net209584), .Y(n48330)
         );
  AOI21X1 U25847 ( .A0(n48292), .A1(n48335), .B0(n48291), .Y(n48294) );
  NAND2X1 U25848 ( .A(n41374), .B(n48288), .Y(n48292) );
  OR2X4 U25849 ( .A(n48290), .B(n48289), .Y(n41374) );
  CLKINVX1 U25850 ( .A(n48336), .Y(n48290) );
  OR2X2 U25851 ( .A(net209547), .B(n48348), .Y(n41216) );
  AOI21X2 U25852 ( .A0(n48371), .A1(n48370), .B0(n49502), .Y(n48372) );
  NAND2XL U25853 ( .A(n41344), .B(n11732), .Y(n48371) );
  OAI2BB1X1 U25854 ( .A0N(n11706), .A1N(n41664), .B0(n11705), .Y(n48277) );
  CLKINVX3 U25855 ( .A(net210615), .Y(net210211) );
  INVXL U25856 ( .A(n12326), .Y(n48423) );
  NAND2X1 U25857 ( .A(n41352), .B(n12292), .Y(n48517) );
  OR2X1 U25858 ( .A(n11211), .B(net209211), .Y(n41352) );
  OAI21XL U25859 ( .A0(net171440), .A1(n48418), .B0(n11084), .Y(n48420) );
  OAI2BB1X1 U25860 ( .A0N(n41659), .A1N(n41660), .B0(n12493), .Y(n48388) );
  INVXL U25861 ( .A(n11057), .Y(net209197) );
  AO21X2 U25862 ( .A0(n48052), .A1(n48051), .B0(n48050), .Y(n41700) );
  NAND2X1 U25863 ( .A(net209311), .B(net209308), .Y(net210548) );
  CLKINVX1 U25864 ( .A(n11035), .Y(net209179) );
  OAI211X1 U25865 ( .A0(n11070), .A1(n11071), .B0(n11072), .C0(n11073), .Y(
        n11068) );
  AOI21X1 U25866 ( .A0(n48540), .A1(n12255), .B0(net151494), .Y(n48541) );
  CLKINVX1 U25867 ( .A(n11639), .Y(net209463) );
  NAND3X2 U25868 ( .A(n11035), .B(n10820), .C(n11036), .Y(n11033) );
  CLKINVX1 U25869 ( .A(net259645), .Y(net171146) );
  NAND2X6 U25870 ( .A(n41372), .B(n10808), .Y(n48550) );
  NAND2X1 U25871 ( .A(n10806), .B(n37012), .Y(n41372) );
  NAND2X4 U25872 ( .A(n41215), .B(net151251), .Y(n11627) );
  CLKINVX1 U25873 ( .A(n40404), .Y(net151251) );
  XOR2XL U25874 ( .A(n41833), .B(n36901), .Y(n44080) );
  NOR2X2 U25875 ( .A(n46195), .B(n48132), .Y(n46199) );
  NOR4X1 U25876 ( .A(n44653), .B(n44652), .C(n44651), .D(n44650), .Y(n44659)
         );
  NOR4X1 U25877 ( .A(n44645), .B(n44644), .C(n44643), .D(n44642), .Y(n44661)
         );
  NOR2X4 U25878 ( .A(n47336), .B(net209314), .Y(n47346) );
  NOR2X2 U25879 ( .A(n47369), .B(net209311), .Y(n47379) );
  NOR2X1 U25880 ( .A(n12065), .B(n47189), .Y(n47193) );
  NOR2XL U25881 ( .A(n12078), .B(n46093), .Y(n46097) );
  XOR2XL U25882 ( .A(n42494), .B(n42069), .Y(n47615) );
  NOR2XL U25883 ( .A(n12152), .B(n45738), .Y(n45742) );
  NAND2X2 U25884 ( .A(n41256), .B(n41257), .Y(n29322) );
  NAND2XL U25885 ( .A(n33920), .B(n37015), .Y(n41257) );
  NOR4X1 U25886 ( .A(n44864), .B(n44863), .C(n44862), .D(n44861), .Y(n44870)
         );
  XOR2X1 U25887 ( .A(n41824), .B(n42602), .Y(n44854) );
  NOR4X1 U25888 ( .A(n44136), .B(n44135), .C(n44134), .D(n44133), .Y(n44152)
         );
  NOR4X1 U25889 ( .A(n44144), .B(n44143), .C(n44142), .D(n44141), .Y(n44150)
         );
  NOR4X1 U25890 ( .A(n44113), .B(n44112), .C(n44111), .D(n44110), .Y(n44119)
         );
  NOR2X4 U25891 ( .A(n46321), .B(net209903), .Y(n46331) );
  NOR2X4 U25892 ( .A(n46412), .B(n48173), .Y(n46422) );
  NAND4X2 U25893 ( .A(n46499), .B(n46498), .C(n46497), .D(n46496), .Y(n48443)
         );
  NOR2X6 U25894 ( .A(n46533), .B(n48158), .Y(n46543) );
  NAND4X2 U25895 ( .A(n46564), .B(n46563), .C(n36934), .D(net212262), .Y(
        n47705) );
  NOR4X1 U25896 ( .A(n46558), .B(n46557), .C(n46556), .D(n46555), .Y(n46564)
         );
  NOR4X1 U25897 ( .A(n46562), .B(n46561), .C(n46560), .D(n46559), .Y(n46563)
         );
  NOR2X2 U25898 ( .A(n44060), .B(net209589), .Y(n44070) );
  NOR2X2 U25899 ( .A(n36985), .B(n37228), .Y(n39780) );
  NAND4X4 U25900 ( .A(n44732), .B(n44731), .C(n44730), .D(n44729), .Y(n48171)
         );
  INVX1 U25901 ( .A(net209873), .Y(net210702) );
  NOR2X1 U25902 ( .A(n46282), .B(net210677), .Y(n46292) );
  NAND4X6 U25903 ( .A(n46204), .B(n46203), .C(n46202), .D(n46201), .Y(n48426)
         );
  NOR4X1 U25904 ( .A(n25196), .B(n25197), .C(n25198), .D(n25199), .Y(n44425)
         );
  CLKINVX3 U25905 ( .A(n46573), .Y(n46574) );
  NAND2X1 U25906 ( .A(net210771), .B(net210770), .Y(n39370) );
  NAND4X2 U25907 ( .A(n44533), .B(n44532), .C(n44531), .D(n44530), .Y(n45727)
         );
  NAND4X6 U25908 ( .A(n45377), .B(n45376), .C(n45375), .D(n45374), .Y(n48159)
         );
  NAND4X2 U25909 ( .A(n45346), .B(n45345), .C(n45344), .D(n45343), .Y(n48160)
         );
  NAND4X4 U25910 ( .A(n45319), .B(n45318), .C(n45317), .D(n45316), .Y(n48138)
         );
  NOR2X4 U25911 ( .A(n45309), .B(net209631), .Y(n45319) );
  NOR2X1 U25912 ( .A(n37373), .B(n37044), .Y(n41070) );
  NOR2X1 U25913 ( .A(n37374), .B(n37045), .Y(n41069) );
  NAND2XL U25914 ( .A(n12957), .B(n12954), .Y(n39648) );
  INVX1 U25915 ( .A(n12962), .Y(net151600) );
  NOR2X1 U25916 ( .A(n37165), .B(n37411), .Y(n39903) );
  NAND3X1 U25917 ( .A(net212136), .B(net212135), .C(net212137), .Y(
        n_cell_301249_net267415) );
  CLKBUFX3 U25918 ( .A(n12847), .Y(net260470) );
  NAND2X1 U25919 ( .A(net212196), .B(net212195), .Y(n40695) );
  NAND2X1 U25920 ( .A(net212190), .B(net212192), .Y(n40686) );
  NAND4X4 U25921 ( .A(n45136), .B(n45135), .C(n45134), .D(n45133), .Y(n48156)
         );
  NOR4X1 U25922 ( .A(n45132), .B(n45131), .C(n45130), .D(n45129), .Y(n45133)
         );
  NAND3X4 U25923 ( .A(n45024), .B(n45023), .C(net209624), .Y(n46595) );
  NOR4X1 U25924 ( .A(n44998), .B(n44997), .C(n44996), .D(n44995), .Y(n45024)
         );
  NAND4X6 U25925 ( .A(n44825), .B(n44824), .C(n44823), .D(n44822), .Y(
        net209893) );
  NOR4X1 U25926 ( .A(n43974), .B(n43973), .C(n43972), .D(n43971), .Y(n43975)
         );
  NOR4X1 U25927 ( .A(n43928), .B(n43927), .C(n43926), .D(n43925), .Y(n43934)
         );
  NOR4X1 U25928 ( .A(n43924), .B(n43923), .C(n43922), .D(n43921), .Y(n43935)
         );
  NOR4X1 U25929 ( .A(n27576), .B(n27577), .C(n27578), .D(n27579), .Y(n44170)
         );
  NAND4X1 U25930 ( .A(n43176), .B(n43175), .C(n43174), .D(n43173), .Y(n11661)
         );
  NAND4X1 U25931 ( .A(n43167), .B(n43166), .C(n43165), .D(n43164), .Y(
        net209476) );
  NAND2X1 U25932 ( .A(n40968), .B(net216502), .Y(n40789) );
  NOR2X1 U25933 ( .A(n37390), .B(n37115), .Y(n40968) );
  NAND2X4 U25934 ( .A(n48443), .B(n48435), .Y(net210579) );
  NAND4X2 U25935 ( .A(n46473), .B(n46472), .C(n46471), .D(n46470), .Y(n46478)
         );
  NAND4X6 U25936 ( .A(n47001), .B(n47000), .C(n46999), .D(n46998), .Y(n12344)
         );
  NAND4X4 U25937 ( .A(n45674), .B(n45673), .C(n45672), .D(n45671), .Y(
        net209267) );
  NAND2X1 U25938 ( .A(n39949), .B(net212694), .Y(n39413) );
  NOR2X1 U25939 ( .A(n10184), .B(n46194), .Y(net212691) );
  AND2X2 U25940 ( .A(net216366), .B(net216367), .Y(n40966) );
  AND2X4 U25941 ( .A(n47996), .B(n48000), .Y(net234521) );
  AND2X2 U25942 ( .A(n47974), .B(n47997), .Y(net234523) );
  OAI21XL U25943 ( .A0(n39343), .A1(n11264), .B0(n40703), .Y(n40528) );
  NOR2BX1 U25944 ( .AN(n40702), .B(n40701), .Y(n40527) );
  NAND2BX1 U25945 ( .AN(n40431), .B(net213633), .Y(net209111) );
  NAND2X1 U25946 ( .A(n40596), .B(net213636), .Y(n40431) );
  NAND2X1 U25947 ( .A(net211631), .B(net211630), .Y(n40585) );
  NAND2X1 U25948 ( .A(n40588), .B(net211626), .Y(n40440) );
  NOR2X2 U25949 ( .A(n37058), .B(n37408), .Y(n39966) );
  NOR2X1 U25950 ( .A(n37077), .B(n37437), .Y(n39968) );
  INVXL U25951 ( .A(n12316), .Y(net151751) );
  NOR2XL U25952 ( .A(n12032), .B(n45828), .Y(n45832) );
  NAND2BX2 U25953 ( .AN(n39435), .B(net213125), .Y(n10827) );
  NAND2X1 U25954 ( .A(n39943), .B(net213126), .Y(n39435) );
  NOR2X1 U25955 ( .A(n37057), .B(n37412), .Y(n39943) );
  NOR2XL U25956 ( .A(net209513), .B(n39704), .Y(n39731) );
  INVXL U25957 ( .A(n11732), .Y(n39704) );
  NOR4X1 U25958 ( .A(n26879), .B(n26880), .C(n26881), .D(n26882), .Y(net215228) );
  NOR2X2 U25959 ( .A(n36983), .B(n37332), .Y(n39452) );
  NAND4BX1 U25960 ( .AN(n37110), .B(net216363), .C(net216360), .D(net216361),
        .Y(n11607) );
  NAND3X1 U25961 ( .A(net214787), .B(net214786), .C(n40410), .Y(n11605) );
  NOR2X1 U25962 ( .A(n36955), .B(n37267), .Y(n40410) );
  NAND2X2 U25963 ( .A(n48034), .B(n48029), .Y(n47774) );
  NAND2X2 U25964 ( .A(n48032), .B(n48027), .Y(n47772) );
  NAND2X4 U25965 ( .A(n48038), .B(n48036), .Y(net210620) );
  NAND2X2 U25966 ( .A(n48040), .B(n48037), .Y(net210587) );
  NOR2X1 U25967 ( .A(n20106), .B(n20105), .Y(net211475) );
  NOR2X2 U25968 ( .A(n37026), .B(n37329), .Y(n39886) );
  NOR2X1 U25969 ( .A(n37074), .B(n37327), .Y(n39884) );
  NAND4X1 U25970 ( .A(n45684), .B(n45683), .C(n45682), .D(n45681), .Y(
        net209268) );
  NOR2X2 U25971 ( .A(n37031), .B(n37330), .Y(n39887) );
  NOR2X1 U25972 ( .A(n37081), .B(n37328), .Y(n39885) );
  BUFX2 U25973 ( .A(n11093), .Y(n40398) );
  CLKINVX2 U25974 ( .A(net209225), .Y(net171443) );
  NOR2X2 U25975 ( .A(n12479), .B(n43321), .Y(n43325) );
  NOR4X1 U25976 ( .A(n29264), .B(n29265), .C(n29266), .D(n29267), .Y(n43625)
         );
  AND2X4 U25977 ( .A(net213702), .B(net213701), .Y(n39308) );
  CLKAND2X4 U25978 ( .A(n48138), .B(n48160), .Y(net234529) );
  NAND3X2 U25979 ( .A(net215905), .B(net215906), .C(net215904), .Y(n39327) );
  NOR2X1 U25980 ( .A(n37370), .B(n37146), .Y(n41088) );
  NAND2BX1 U25981 ( .AN(n40406), .B(n_cell_301249_net267239), .Y(
        n_cell_303546_net275934) );
  NAND2X1 U25982 ( .A(net216426), .B(net216425), .Y(n40406) );
  NOR2X1 U25983 ( .A(n36970), .B(n37273), .Y(n_cell_301249_net267239) );
  NOR2X1 U25984 ( .A(n37160), .B(n37458), .Y(n41159) );
  NOR2X1 U25985 ( .A(n37094), .B(n37435), .Y(n41161) );
  NOR2X1 U25986 ( .A(n37092), .B(n37457), .Y(n41128) );
  NOR2X1 U25987 ( .A(n37151), .B(n37492), .Y(n40946) );
  NOR2X1 U25988 ( .A(n19700), .B(n19699), .Y(net211263) );
  CLKINVX4 U25989 ( .A(n39648), .Y(n10715) );
  OR4XL U25990 ( .A(net151600), .B(net151601), .C(n37199), .D(n36948), .Y(
        n39647) );
  NOR2X1 U25991 ( .A(n19962), .B(n19961), .Y(n47075) );
  NOR2X1 U25992 ( .A(n20014), .B(n20012), .Y(n47065) );
  NAND2BX1 U25993 ( .AN(n39348), .B(net210507), .Y(n10672) );
  NAND2X1 U25994 ( .A(n39909), .B(net210510), .Y(n39348) );
  NAND4X1 U25995 ( .A(n47941), .B(n47940), .C(n47939), .D(n47938), .Y(n12878)
         );
  CLKINVX1 U25996 ( .A(net260474), .Y(net151554) );
  CLKINVX1 U25997 ( .A(net260470), .Y(net151555) );
  NAND2BX1 U25998 ( .AN(n_cell_301249_net267201), .B(net212184), .Y(
        n_cell_303546_net276009) );
  NAND3X1 U25999 ( .A(net212186), .B(net212185), .C(net212187), .Y(
        n_cell_301249_net267201) );
  NAND3X1 U26000 ( .A(net216345), .B(net216344), .C(n40409), .Y(n11606) );
  NOR2X1 U26001 ( .A(n36956), .B(n37268), .Y(n40409) );
  NOR2X1 U26002 ( .A(n37061), .B(n37322), .Y(n40965) );
  NAND3X1 U26003 ( .A(net216327), .B(net216326), .C(n40408), .Y(n11600) );
  NOR2X1 U26004 ( .A(n36952), .B(n37266), .Y(n40408) );
  NOR2X1 U26005 ( .A(n37060), .B(n37427), .Y(n40963) );
  NAND4BX1 U26006 ( .AN(n37002), .B(net216336), .C(net216333), .D(net216334),
        .Y(n10319) );
  NOR2X1 U26007 ( .A(n37062), .B(n37426), .Y(n40964) );
  NAND3X1 U26008 ( .A(net216285), .B(net216284), .C(net216286), .Y(
        n_cell_301249_net267373) );
  NAND3X4 U26009 ( .A(n45256), .B(n45255), .C(net210475), .Y(net212214) );
  NAND4X2 U26010 ( .A(n45227), .B(n45226), .C(n45225), .D(n45224), .Y(
        net210695) );
  NAND4X4 U26011 ( .A(n45196), .B(n45195), .C(n45194), .D(n45193), .Y(
        net209900) );
  NOR2X4 U26012 ( .A(n45186), .B(net209605), .Y(n45196) );
  NAND2X2 U26013 ( .A(n46595), .B(n48143), .Y(net210699) );
  NAND2XL U26014 ( .A(net214515), .B(net234527), .Y(n39571) );
  INVXL U26015 ( .A(net210682), .Y(net214515) );
  NOR2X1 U26016 ( .A(n36975), .B(n37222), .Y(n39302) );
  NOR2X2 U26017 ( .A(n37301), .B(n37008), .Y(n39790) );
  NAND2X1 U26018 ( .A(n39786), .B(net215292), .Y(n39325) );
  NOR2X2 U26019 ( .A(n37103), .B(n37316), .Y(n39786) );
  NAND2X2 U26020 ( .A(n39785), .B(net215301), .Y(n39324) );
  NOR2X1 U26021 ( .A(n37104), .B(n37320), .Y(n39785) );
  OR3X2 U26022 ( .A(net171245), .B(net171247), .C(n12047), .Y(n39580) );
  NOR2X1 U26023 ( .A(n37051), .B(n37461), .Y(n40961) );
  CLKBUFX3 U26024 ( .A(n11970), .Y(net260277) );
  NAND3X1 U26025 ( .A(n40783), .B(net216520), .C(net216517), .Y(n11960) );
  NOR2X1 U26026 ( .A(n37389), .B(n37117), .Y(n40783) );
  NAND2X1 U26027 ( .A(n40969), .B(net216511), .Y(n40782) );
  NOR2X1 U26028 ( .A(n37391), .B(n37118), .Y(n40969) );
  NAND4X2 U26029 ( .A(n44929), .B(n44928), .C(n44927), .D(n44926), .Y(n47727)
         );
  NOR4X1 U26030 ( .A(n44921), .B(n44920), .C(n44919), .D(n44918), .Y(n44927)
         );
  NOR4X1 U26031 ( .A(n44913), .B(n44912), .C(n44911), .D(n44910), .Y(n44929)
         );
  NAND4BBX2 U26032 ( .AN(n44949), .BN(n44948), .C(n41653), .D(n41654), .Y(
        n41652) );
  NOR4X1 U26033 ( .A(n45428), .B(n45427), .C(n45426), .D(n45425), .Y(n45434)
         );
  NOR4X1 U26034 ( .A(n45432), .B(n45431), .C(n45430), .D(n45429), .Y(n45433)
         );
  NOR2X2 U26035 ( .A(n36937), .B(n37214), .Y(n39457) );
  NOR2X4 U26036 ( .A(n37010), .B(n37232), .Y(n39465) );
  NOR2X2 U26037 ( .A(n36938), .B(n37213), .Y(n39456) );
  CLKBUFX3 U26038 ( .A(n11761), .Y(n40393) );
  NAND4X2 U26039 ( .A(n43258), .B(n43257), .C(n43256), .D(n43255), .Y(n11672)
         );
  CLKBUFX3 U26040 ( .A(n11130), .Y(n40397) );
  INVX1 U26041 ( .A(n12344), .Y(net151673) );
  CLKINVX1 U26042 ( .A(net209267), .Y(net171425) );
  INVXL U26043 ( .A(net209268), .Y(net171427) );
  NAND4X4 U26044 ( .A(n45669), .B(n45668), .C(n45667), .D(n45666), .Y(n11138)
         );
  NAND4X4 U26045 ( .A(n45659), .B(n45658), .C(n45657), .D(n45656), .Y(n11139)
         );
  NAND4X4 U26046 ( .A(n45664), .B(n45663), .C(n45662), .D(n45661), .Y(n11140)
         );
  NAND2X2 U26047 ( .A(net210919), .B(net209303), .Y(net210539) );
  NAND2X1 U26048 ( .A(n48461), .B(n48464), .Y(net210561) );
  NAND4X2 U26049 ( .A(n46183), .B(n46182), .C(n46181), .D(n46180), .Y(n10257)
         );
  NAND2BX1 U26050 ( .AN(n40407), .B(net213537), .Y(net209136) );
  NAND2X1 U26051 ( .A(n40594), .B(net213540), .Y(n40407) );
  NOR2X1 U26052 ( .A(n37095), .B(n37450), .Y(n40594) );
  NAND2X1 U26053 ( .A(n41151), .B(net213545), .Y(n40790) );
  NOR2X1 U26054 ( .A(n37090), .B(n37459), .Y(n41151) );
  CLKBUFX3 U26055 ( .A(n12228), .Y(net260332) );
  NAND2X1 U26056 ( .A(n40640), .B(net212025), .Y(n40420) );
  AND2X2 U26057 ( .A(net212024), .B(net212023), .Y(n40640) );
  NAND2BX1 U26058 ( .AN(n40949), .B(net211597), .Y(n_cell_301249_net269874) );
  NAND2X1 U26059 ( .A(n40948), .B(net211600), .Y(n40949) );
  NAND2X1 U26060 ( .A(n40684), .B(net210371), .Y(n40446) );
  NAND2X1 U26061 ( .A(n40682), .B(net211466), .Y(n40454) );
  NOR2X1 U26062 ( .A(n37481), .B(n37176), .Y(n41118) );
  NAND2X2 U26063 ( .A(n39962), .B(net213405), .Y(n39404) );
  NOR2X1 U26064 ( .A(n37036), .B(n37467), .Y(n39962) );
  NAND2X2 U26065 ( .A(n39959), .B(net212729), .Y(n39407) );
  OR4XL U26066 ( .A(net171421), .B(net171423), .C(net151612), .D(net151751),
        .Y(n39510) );
  NOR2X1 U26067 ( .A(n22331), .B(n22330), .Y(n46160) );
  NAND4X2 U26068 ( .A(n46152), .B(n46151), .C(n46150), .D(n46149), .Y(n11114)
         );
  NOR2X1 U26069 ( .A(n22351), .B(n22350), .Y(n46150) );
  NOR4X1 U26070 ( .A(n24772), .B(n24773), .C(n24774), .D(n24775), .Y(n44555)
         );
  NOR4X1 U26071 ( .A(n24926), .B(n24927), .C(n24928), .D(n24929), .Y(n44510)
         );
  CLKINVX1 U26072 ( .A(n10319), .Y(net171169) );
  CLKBUFX3 U26073 ( .A(net209441), .Y(net260900) );
  NAND4X1 U26074 ( .A(n11605), .B(n11600), .C(n11601), .D(n11606), .Y(n10311)
         );
  NAND2X2 U26075 ( .A(n39879), .B(net211150), .Y(n39371) );
  NAND2X2 U26076 ( .A(n39880), .B(net211155), .Y(n39372) );
  INVXL U26077 ( .A(n12931), .Y(net151860) );
  INVXL U26078 ( .A(n40398), .Y(net171447) );
  NAND3XL U26079 ( .A(n11095), .B(n11094), .C(n11092), .Y(n10839) );
  OR4XL U26080 ( .A(net151848), .B(net171445), .C(net171443), .D(net151738),
        .Y(n39511) );
  NAND2X1 U26081 ( .A(n39800), .B(net216023), .Y(n39318) );
  NOR2X2 U26082 ( .A(n37108), .B(n37311), .Y(n39800) );
  NAND3X1 U26083 ( .A(net216407), .B(net216408), .C(n40794), .Y(n11613) );
  NOR2X1 U26084 ( .A(n36971), .B(n37280), .Y(n40794) );
  CLKBUFX3 U26085 ( .A(net209960), .Y(n40386) );
  NAND4X1 U26086 ( .A(n46864), .B(n46863), .C(n46862), .D(n46861), .Y(n11324)
         );
  NAND2BX1 U26087 ( .AN(n_cell_301249_net267063), .B(net211793), .Y(n12867) );
  NAND3X1 U26088 ( .A(net211795), .B(net211796), .C(net211794), .Y(
        n_cell_301249_net267063) );
  NOR2X1 U26089 ( .A(n37372), .B(n37149), .Y(n41068) );
  NOR2X1 U26090 ( .A(n36990), .B(n37293), .Y(n_cell_301249_net267595) );
  CLKBUFX3 U26091 ( .A(n10429), .Y(net259653) );
  CLKBUFX3 U26092 ( .A(n10428), .Y(net259649) );
  NOR2X1 U26093 ( .A(n36966), .B(n37275), .Y(n_cell_301249_net267233) );
  CLKBUFX3 U26094 ( .A(n12445), .Y(net260367) );
  CLKINVX1 U26095 ( .A(n11614), .Y(net171151) );
  NAND2X1 U26096 ( .A(net215041), .B(net215040), .Y(n40434) );
  NOR2X1 U26097 ( .A(n36988), .B(n37291), .Y(n_cell_301249_net267903) );
  NAND2BX1 U26098 ( .AN(n40438), .B(n_cell_301249_net267932), .Y(n11566) );
  NAND2X1 U26099 ( .A(net215014), .B(net215013), .Y(n40438) );
  NOR2X1 U26100 ( .A(n36986), .B(n37284), .Y(n_cell_301249_net267932) );
  NAND2BX1 U26101 ( .AN(n40437), .B(n_cell_301249_net267909), .Y(n11567) );
  NAND2X1 U26102 ( .A(net215050), .B(net215049), .Y(n40437) );
  NOR2X1 U26103 ( .A(n36987), .B(n37290), .Y(n_cell_301249_net267909) );
  NAND4BBX1 U26104 ( .AN(n37394), .BN(n37003), .C(net215059), .D(net215057),
        .Y(n11565) );
  NAND4X1 U26105 ( .A(n43334), .B(n43333), .C(n43332), .D(n43331), .Y(n10157)
         );
  NOR2X1 U26106 ( .A(n31174), .B(n31173), .Y(n43332) );
  NAND2BX1 U26107 ( .AN(n_cell_301249_net267325), .B(net213522), .Y(n10968) );
  NAND2X1 U26108 ( .A(n41160), .B(net213525), .Y(n_cell_301249_net267325) );
  NOR2X1 U26109 ( .A(n37076), .B(n37504), .Y(n41160) );
  NAND2X1 U26110 ( .A(n41126), .B(net213611), .Y(n_cell_301249_net267769) );
  NOR2X1 U26111 ( .A(n37088), .B(n37455), .Y(n41126) );
  NAND2X1 U26112 ( .A(n41127), .B(net213626), .Y(n_cell_301249_net267700) );
  NAND2X1 U26113 ( .A(n40655), .B(net212051), .Y(n40416) );
  AND2X2 U26114 ( .A(net212050), .B(net212049), .Y(n40655) );
  NOR2X1 U26115 ( .A(n37157), .B(n37387), .Y(n41062) );
  NOR2X1 U26116 ( .A(n37155), .B(n37486), .Y(n40587) );
  NOR2X1 U26117 ( .A(n37072), .B(n37386), .Y(n41061) );
  NAND2BX1 U26118 ( .AN(n40428), .B(net213497), .Y(n12210) );
  NAND2X1 U26119 ( .A(n40638), .B(net213500), .Y(n40428) );
  NOR2X1 U26120 ( .A(n37071), .B(n37385), .Y(n41104) );
  CLKINVX1 U26121 ( .A(net209992), .Y(net171542) );
  NAND2X1 U26122 ( .A(n40589), .B(net211606), .Y(n40445) );
  CLKINVX1 U26123 ( .A(n_cell_301249_net269874), .Y(net238789) );
  NAND2BX1 U26124 ( .AN(n40447), .B(net210363), .Y(n12824) );
  NAND2X1 U26125 ( .A(n40683), .B(net210366), .Y(n40447) );
  NAND3XL U26126 ( .A(n11397), .B(n11396), .C(n11399), .Y(n10702) );
  OR4XL U26127 ( .A(net151746), .B(net151744), .C(n37253), .D(net171550), .Y(
        n39653) );
  NAND3XL U26128 ( .A(n11371), .B(n11372), .C(n39353), .Y(n10028) );
  NOR2X1 U26129 ( .A(n39632), .B(n39633), .Y(n39353) );
  INVXL U26130 ( .A(n40394), .Y(n39633) );
  INVXL U26131 ( .A(n11369), .Y(n39632) );
  NOR2X1 U26132 ( .A(n37134), .B(n37403), .Y(n41072) );
  NAND2X1 U26133 ( .A(n39913), .B(net210499), .Y(n39346) );
  NAND2BX1 U26134 ( .AN(n40780), .B(net211982), .Y(n12873) );
  NAND2X1 U26135 ( .A(n41073), .B(net211984), .Y(n40780) );
  NOR2X1 U26136 ( .A(n37150), .B(n37384), .Y(n41073) );
  CLKINVX1 U26137 ( .A(n12878), .Y(net151426) );
  AND4X1 U26138 ( .A(n46838), .B(n46837), .C(n46836), .D(n46835), .Y(net238947) );
  NOR2X1 U26139 ( .A(n37490), .B(n37175), .Y(n41065) );
  NAND2BX1 U26140 ( .AN(n_cell_301249_net267331), .B(net213507), .Y(n10966) );
  NAND2X1 U26141 ( .A(n41162), .B(net213510), .Y(n_cell_301249_net267331) );
  CLKBUFX3 U26142 ( .A(n12634), .Y(net260412) );
  NAND2X1 U26143 ( .A(n41005), .B(net216158), .Y(n_cell_301249_net267810) );
  NAND2BX1 U26144 ( .AN(n_cell_301249_net267670), .B(net216184), .Y(n12806) );
  NAND2X1 U26145 ( .A(n41002), .B(net216185), .Y(n_cell_301249_net267670) );
  NAND2X4 U26146 ( .A(n12747), .B(n12751), .Y(n10577) );
  NAND2X6 U26147 ( .A(n37217), .B(net171314), .Y(n12087) );
  XOR2XL U26148 ( .A(n42207), .B(n41323), .Y(n31834) );
  NAND4X1 U26149 ( .A(n44585), .B(n44584), .C(n44583), .D(n44582), .Y(n11662)
         );
  NAND4X1 U26150 ( .A(n44639), .B(n44638), .C(n44637), .D(n44636), .Y(n12474)
         );
  NOR2X1 U26151 ( .A(n37392), .B(n37007), .Y(n39817) );
  CLKBUFX3 U26152 ( .A(n12629), .Y(net271999) );
  NAND2X1 U26153 ( .A(n39821), .B(net216808), .Y(n39336) );
  NOR2X1 U26154 ( .A(n37388), .B(n37114), .Y(n39821) );
  CLKBUFX3 U26155 ( .A(n12801), .Y(n40388) );
  NAND2X1 U26156 ( .A(n40976), .B(net216871), .Y(n_cell_301249_net266916) );
  CLKBUFX3 U26157 ( .A(n10493), .Y(net259747) );
  NAND3X1 U26158 ( .A(n11960), .B(n11961), .C(n39286), .Y(n10492) );
  NOR2X1 U26159 ( .A(n39555), .B(n39556), .Y(n39286) );
  CLKBUFX3 U26160 ( .A(net214757), .Y(net272625) );
  NOR2X1 U26161 ( .A(n36969), .B(n37276), .Y(n_cell_301249_net267786) );
  CLKINVX1 U26162 ( .A(n10086), .Y(net151265) );
  CLKINVX1 U26163 ( .A(n39741), .Y(n10091) );
  NAND4BXL U26164 ( .AN(net151258), .B(net214730), .C(n12493), .D(net214729),
        .Y(n39741) );
  NAND4X2 U26165 ( .A(n43311), .B(n43310), .C(n43309), .D(n43308), .Y(n10089)
         );
  NAND3XL U26166 ( .A(n11669), .B(n11672), .C(n39450), .Y(n10085) );
  NOR2BXL U26167 ( .AN(n11673), .B(net209479), .Y(n39450) );
  NAND2X1 U26168 ( .A(n12482), .B(n12486), .Y(n10093) );
  NAND2X1 U26169 ( .A(n40721), .B(net213223), .Y(n40453) );
  CLKBUFX3 U26170 ( .A(n12651), .Y(net260427) );
  CLKBUFX3 U26171 ( .A(n11955), .Y(net260251) );
  NOR2X1 U26172 ( .A(n37257), .B(n40967), .Y(n40788) );
  NAND2X1 U26173 ( .A(net216492), .B(net216491), .Y(n40967) );
  NAND2X2 U26174 ( .A(n39950), .B(net213345), .Y(n39425) );
  NOR2X1 U26175 ( .A(n36997), .B(n37315), .Y(n39950) );
  NAND3X1 U26176 ( .A(net213354), .B(net213355), .C(net213353), .Y(n39411) );
  NOR2X1 U26177 ( .A(n12085), .B(n45692), .Y(net213352) );
  NOR2X1 U26178 ( .A(n23758), .B(n23757), .Y(net213354) );
  INVXL U26179 ( .A(n40397), .Y(net171435) );
  NAND3XL U26180 ( .A(n11140), .B(n11139), .C(n11138), .Y(n10877) );
  NOR2X1 U26181 ( .A(n22978), .B(n22977), .Y(n45907) );
  NAND2BX1 U26182 ( .AN(n_cell_301249_net267263), .B(net213572), .Y(n10973) );
  NAND2X1 U26183 ( .A(n41133), .B(net213575), .Y(n_cell_301249_net267263) );
  NOR2X1 U26184 ( .A(n37161), .B(n37505), .Y(n41133) );
  NAND2BX2 U26185 ( .AN(n_cell_301249_net267189), .B(net213567), .Y(
        n_cell_303546_net275998) );
  NAND2X1 U26186 ( .A(n41135), .B(net213570), .Y(n_cell_301249_net267189) );
  NOR2X1 U26187 ( .A(n37169), .B(n37507), .Y(n41135) );
  NAND2X1 U26188 ( .A(n41136), .B(net213555), .Y(n_cell_301249_net267117) );
  NOR2X1 U26189 ( .A(n37083), .B(n37453), .Y(n41136) );
  CLKBUFX3 U26190 ( .A(n12230), .Y(net271956) );
  NAND2X1 U26191 ( .A(n37472), .B(net213532), .Y(n10983) );
  NOR2X1 U26192 ( .A(n37087), .B(n37460), .Y(n41149) );
  NAND2X1 U26193 ( .A(n41137), .B(net213530), .Y(n_cell_301249_net267123) );
  NOR2X1 U26194 ( .A(n37084), .B(n37454), .Y(n41137) );
  CLKINVX1 U26195 ( .A(net209136), .Y(net171401) );
  CLKBUFX3 U26196 ( .A(n10793), .Y(net259873) );
  CLKINVX1 U26197 ( .A(n10982), .Y(net171398) );
  CLKINVX1 U26198 ( .A(net260332), .Y(net151536) );
  CLKINVX1 U26199 ( .A(net212037), .Y(net171406) );
  NAND3X1 U26200 ( .A(n39287), .B(net216880), .C(net216877), .Y(n10503) );
  AND2X2 U26201 ( .A(net216879), .B(net216878), .Y(n39287) );
  NAND3X2 U26202 ( .A(n40776), .B(net216907), .C(net216904), .Y(n11968) );
  NOR2X1 U26203 ( .A(n37099), .B(n37425), .Y(n40776) );
  NAND2BX1 U26204 ( .AN(n39285), .B(net216427), .Y(n10484) );
  NAND2X1 U26205 ( .A(n39829), .B(net216428), .Y(n39285) );
  NOR2X1 U26206 ( .A(n37041), .B(n37429), .Y(n41139) );
  NAND2BX1 U26207 ( .AN(n40773), .B(net212856), .Y(n10992) );
  NAND2X1 U26208 ( .A(n41140), .B(net212859), .Y(n40773) );
  NOR2X1 U26209 ( .A(n37033), .B(n37433), .Y(n41140) );
  NAND2BX1 U26210 ( .AN(n40778), .B(net212851), .Y(n10990) );
  NAND2X1 U26211 ( .A(n41144), .B(net212854), .Y(n40778) );
  BUFX4 U26212 ( .A(n34469), .Y(n42482) );
  NAND2X1 U26213 ( .A(n12196), .B(n12194), .Y(n10926) );
  NOR2BX1 U26214 ( .AN(net215134), .B(n37363), .Y(n41015) );
  NAND2BX1 U26215 ( .AN(n_cell_301249_net268056), .B(net211468), .Y(n12821) );
  NAND3X1 U26216 ( .A(net211470), .B(net211469), .C(net211471), .Y(
        n_cell_301249_net268056) );
  NAND2BX1 U26217 ( .AN(n40456), .B(net215186), .Y(n12594) );
  NAND2X1 U26218 ( .A(n40634), .B(net215189), .Y(n40456) );
  NOR2X1 U26219 ( .A(n37128), .B(n37421), .Y(n40634) );
  NOR2X1 U26220 ( .A(n36982), .B(n37381), .Y(n40449) );
  CLKINVX1 U26221 ( .A(net261069), .Y(net171437) );
  CLKINVX1 U26222 ( .A(net209087), .Y(net171439) );
  OR2X1 U26223 ( .A(net238790), .B(n40710), .Y(n_cell_301249_net269872) );
  CLKINVX1 U26224 ( .A(n40713), .Y(net238790) );
  NAND2BX1 U26225 ( .AN(n40800), .B(net211182), .Y(n10612) );
  NAND2X1 U26226 ( .A(n41119), .B(net211184), .Y(n40800) );
  NAND4XL U26227 ( .A(n11717), .B(n11711), .C(n11712), .D(n11718), .Y(n10105)
         );
  CLKBUFX3 U26228 ( .A(n10106), .Y(n40403) );
  CLKBUFX3 U26229 ( .A(n10176), .Y(n40401) );
  NAND3XL U26230 ( .A(n12147), .B(n12146), .C(n39298), .Y(n10177) );
  NOR2XL U26231 ( .A(n39564), .B(net209953), .Y(n39298) );
  INVXL U26232 ( .A(n12073), .Y(n39564) );
  OR2X1 U26233 ( .A(n37337), .B(n_cell_301249_net267171), .Y(n10485) );
  NAND2X1 U26234 ( .A(n40984), .B(net216394), .Y(n_cell_301249_net267171) );
  NOR2X1 U26235 ( .A(n37023), .B(n37323), .Y(n40984) );
  CLKBUFX3 U26236 ( .A(n10165), .Y(n40402) );
  NAND3XL U26237 ( .A(n12026), .B(n12025), .C(n12797), .Y(n10166) );
  NAND4X1 U26238 ( .A(n11326), .B(n11327), .C(n12893), .D(n13019), .Y(n39670)
         );
  NAND3X1 U26239 ( .A(n11324), .B(n11325), .C(n39350), .Y(n10679) );
  NOR2X1 U26240 ( .A(n39627), .B(n39628), .Y(n39350) );
  CLKINVX1 U26241 ( .A(n11515), .Y(n39627) );
  NAND2X1 U26242 ( .A(n39878), .B(net212000), .Y(n39383) );
  NAND2BX1 U26243 ( .AN(n39380), .B(net212002), .Y(n10754) );
  NAND2X1 U26244 ( .A(n39876), .B(net212005), .Y(n39380) );
  NAND2BX1 U26245 ( .AN(n39381), .B(net211987), .Y(n10757) );
  NAND2X1 U26246 ( .A(n39877), .B(net211990), .Y(n39381) );
  NAND3X1 U26247 ( .A(net211994), .B(net211993), .C(net211995), .Y(n39382) );
  OR4X1 U26248 ( .A(net151443), .B(net151444), .C(net151453), .D(net151451),
        .Y(n39666) );
  NAND2X1 U26249 ( .A(n41089), .B(net211780), .Y(n_cell_301249_net267225) );
  NAND2X1 U26250 ( .A(n41067), .B(net211775), .Y(n_cell_301249_net267207) );
  NAND2X1 U26251 ( .A(n41058), .B(net211450), .Y(n_cell_301249_net268172) );
  NAND3X1 U26252 ( .A(net214782), .B(n39765), .C(n39766), .Y(n39764) );
  CLKINVX1 U26253 ( .A(net171278), .Y(n39765) );
  NOR2X1 U26254 ( .A(net151373), .B(net151374), .Y(n39766) );
  CLKINVX1 U26255 ( .A(net214783), .Y(net171278) );
  NAND3X1 U26256 ( .A(n11565), .B(n11567), .C(n11566), .Y(n10295) );
  NAND2BX1 U26257 ( .AN(n_cell_301249_net268190), .B(net215114), .Y(n11886) );
  NAND2X1 U26258 ( .A(n40952), .B(net215117), .Y(n_cell_301249_net268190) );
  CLKINVX1 U26259 ( .A(n40900), .Y(n11897) );
  NAND2X1 U26260 ( .A(n40639), .B(net212081), .Y(n40423) );
  CLKINVX1 U26261 ( .A(n10940), .Y(n39481) );
  NAND2BX1 U26262 ( .AN(n_cell_301249_net267640), .B(net212068), .Y(n11263) );
  NAND3X1 U26263 ( .A(net212070), .B(net212069), .C(net212071), .Y(
        n_cell_301249_net267640) );
  NAND3X1 U26264 ( .A(net211619), .B(net211621), .C(net211620), .Y(
        n_cell_301249_net267855) );
  NAND2X1 U26265 ( .A(n41060), .B(net211611), .Y(n_cell_301249_net267966) );
  CLKINVX1 U26266 ( .A(n_cell_301249_net269872), .Y(n10632) );
  NAND2BX1 U26267 ( .AN(n_cell_301249_net267960), .B(net211613), .Y(n10635) );
  NAND3X1 U26268 ( .A(net211614), .B(net211616), .C(net211615), .Y(
        n_cell_301249_net267960) );
  OR2X1 U26269 ( .A(net238801), .B(n37351), .Y(n39689) );
  CLKINVX1 U26270 ( .A(n_cell_301249_net269738), .Y(net238801) );
  CLKINVX1 U26271 ( .A(net260461), .Y(net151793) );
  NAND2X1 U26272 ( .A(n40597), .B(net213585), .Y(n40442) );
  NOR2X1 U26273 ( .A(n37162), .B(n37500), .Y(n40597) );
  NAND2BX1 U26274 ( .AN(n40791), .B(net211957), .Y(n11299) );
  NAND2X1 U26275 ( .A(n41071), .B(net211959), .Y(n40791) );
  NOR2X1 U26276 ( .A(n37375), .B(n37144), .Y(n41071) );
  NAND2X1 U26277 ( .A(n41112), .B(net211594), .Y(n_cell_301249_net268103) );
  NOR2X1 U26278 ( .A(n37480), .B(n37178), .Y(n41112) );
  NAND2BX1 U26279 ( .AN(n_cell_301249_net268038), .B(net211585), .Y(n10630) );
  NAND2X1 U26280 ( .A(n41059), .B(net211588), .Y(n_cell_301249_net268038) );
  CLKINVX1 U26281 ( .A(net213230), .Y(net171272) );
  NAND2X1 U26282 ( .A(net271999), .B(n39339), .Y(n10611) );
  NOR2X1 U26283 ( .A(n39551), .B(n39781), .Y(n39339) );
  NAND2X1 U26284 ( .A(n11924), .B(n11925), .Y(n39781) );
  NAND2X1 U26285 ( .A(n41000), .B(net214675), .Y(n_cell_301249_net267676) );
  AND2X2 U26286 ( .A(net214674), .B(net214673), .Y(n41000) );
  NAND2X1 U26287 ( .A(n40959), .B(net214681), .Y(n_cell_301249_net267694) );
  NOR2BX1 U26288 ( .AN(net214680), .B(n37360), .Y(n40959) );
  NAND2BX1 U26289 ( .AN(n_cell_301249_net267688), .B(net216202), .Y(n12168) );
  NAND2X1 U26290 ( .A(n40958), .B(net216203), .Y(n_cell_301249_net267688) );
  NAND2BX1 U26291 ( .AN(n_cell_301249_net267682), .B(net214683), .Y(n10471) );
  NAND2X1 U26292 ( .A(n40999), .B(net214686), .Y(n_cell_301249_net267682) );
  NOR2BX1 U26293 ( .AN(net214685), .B(n37356), .Y(n40999) );
  CLKBUFX3 U26294 ( .A(net210704), .Y(net261020) );
  CLKBUFX3 U26295 ( .A(net214755), .Y(net272620) );
  NOR2X1 U26296 ( .A(n37367), .B(n36994), .Y(n_cell_301249_net267980) );
  OR2X1 U26297 ( .A(n37353), .B(n_cell_303546_net276554), .Y(n10434) );
  NAND2X1 U26298 ( .A(net215005), .B(net215004), .Y(n_cell_303546_net276554)
         );
  CLKBUFX3 U26299 ( .A(n10435), .Y(net259677) );
  NAND4X1 U26300 ( .A(net215020), .B(net215021), .C(net215022), .D(net215023),
        .Y(n10436) );
  CLKINVX1 U26301 ( .A(net272625), .Y(net171297) );
  CLKINVX1 U26302 ( .A(net214756), .Y(net171270) );
  NAND3X1 U26303 ( .A(n_cell_303546_net276365), .B(n11575), .C(n39443), .Y(
        n10301) );
  NOR2X1 U26304 ( .A(n39700), .B(n39701), .Y(n39443) );
  CLKINVX1 U26305 ( .A(n11578), .Y(n39700) );
  CLKINVX1 U26306 ( .A(net261422), .Y(net171318) );
  CLKBUFX3 U26307 ( .A(n10303), .Y(net259626) );
  NAND3X1 U26308 ( .A(n_cell_301249_net267607), .B(net216246), .C(net216243),
        .Y(n10302) );
  NOR2X1 U26309 ( .A(n37068), .B(n37286), .Y(n_cell_301249_net267607) );
  NAND2BX1 U26310 ( .AN(net171315), .B(n39763), .Y(n39762) );
  NOR2X1 U26311 ( .A(n_cell_301249_net269635), .B(n11584), .Y(n39763) );
  NAND3X1 U26312 ( .A(net213227), .B(net213226), .C(net213228), .Y(
        n_cell_301249_net268023) );
  NAND2BX1 U26313 ( .AN(n40450), .B(net213205), .Y(n12602) );
  NAND2X1 U26314 ( .A(n40750), .B(net213208), .Y(n40450) );
  NAND2BX1 U26315 ( .AN(n_cell_301249_net268196), .B(net215123), .Y(n11885) );
  NAND2X1 U26316 ( .A(n40953), .B(net215126), .Y(n_cell_301249_net268196) );
  NAND2X1 U26317 ( .A(n40592), .B(net215099), .Y(n40451) );
  NAND4BX2 U26318 ( .AN(n39394), .B(n11029), .C(n11030), .D(n11031), .Y(n10814) );
  CLKINVX1 U26319 ( .A(n40399), .Y(n39394) );
  NAND2X1 U26320 ( .A(net209101), .B(net272417), .Y(n41175) );
  NOR2X1 U26321 ( .A(net171394), .B(n41177), .Y(n41178) );
  NAND2X1 U26322 ( .A(n41124), .B(net212565), .Y(n_cell_301249_net268386) );
  NOR2X1 U26323 ( .A(n37141), .B(n37495), .Y(n41124) );
  NAND2X1 U26324 ( .A(n11884), .B(n11883), .Y(n41016) );
  NOR2X1 U26325 ( .A(net171262), .B(net171259), .Y(n41017) );
  NAND2X1 U26326 ( .A(n40751), .B(net212570), .Y(n40459) );
  NOR2BX1 U26327 ( .AN(net212569), .B(n37358), .Y(n40751) );
  CLKINVX1 U26328 ( .A(n11538), .Y(n39548) );
  NAND2BX1 U26329 ( .AN(n40448), .B(net210348), .Y(n12813) );
  NAND2X1 U26330 ( .A(n40720), .B(net210350), .Y(n40448) );
  CLKINVX1 U26331 ( .A(net260346), .Y(n_cell_303546_net277497) );
  NAND2BXL U26332 ( .AN(n9747), .B(n40593), .Y(n40457) );
  NOR2X1 U26333 ( .A(net260384), .B(n39549), .Y(n40593) );
  NAND2X1 U26334 ( .A(n41057), .B(net211435), .Y(n_cell_301249_net268166) );
  NAND2BX1 U26335 ( .AN(n_cell_301249_net268097), .B(net211453), .Y(n11242) );
  NAND2X1 U26336 ( .A(n41113), .B(net211456), .Y(n_cell_301249_net268097) );
  OAI21XL U26337 ( .A0(net151767), .A1(net209087), .B0(net260302), .Y(n40681)
         );
  CLKINVX1 U26338 ( .A(n10097), .Y(net151325) );
  CLKINVX1 U26339 ( .A(n10113), .Y(net168850) );
  CLKBUFX3 U26340 ( .A(n9768), .Y(net260527) );
  NAND4X1 U26341 ( .A(n43485), .B(n43484), .C(n43483), .D(n43482), .Y(n9768)
         );
  CLKINVX1 U26342 ( .A(n40387), .Y(net151789) );
  CLKINVX1 U26343 ( .A(net260925), .Y(net171283) );
  CLKINVX1 U26344 ( .A(net272583), .Y(net171288) );
  NAND2X1 U26345 ( .A(n12190), .B(n12188), .Y(n11228) );
  CLKINVX1 U26346 ( .A(n9716), .Y(net171380) );
  CLKBUFX3 U26347 ( .A(net218256), .Y(net218152) );
  CLKBUFX3 U26348 ( .A(net218258), .Y(net218148) );
  BUFX2 U26349 ( .A(net217116), .Y(n40315) );
  CLKBUFX3 U26350 ( .A(net218258), .Y(net218146) );
  CLKBUFX3 U26351 ( .A(net218254), .Y(net218156) );
  CLKBUFX3 U26352 ( .A(n9739), .Y(n41199) );
  CLKBUFX3 U26353 ( .A(net218580), .Y(net218294) );
  NOR2X1 U26354 ( .A(net210479), .B(net209620), .Y(n47730) );
  CLKAND2X3 U26355 ( .A(n48439), .B(n48441), .Y(n41373) );
  NOR2X1 U26356 ( .A(net209315), .B(net210583), .Y(n47782) );
  AOI21X1 U26357 ( .A0(net210599), .A1(n47769), .B0(net210601), .Y(n47770) );
  CLKINVX1 U26358 ( .A(net210618), .Y(net210599) );
  AND2X2 U26359 ( .A(net209930), .B(net209893), .Y(n47721) );
  CLKINVX1 U26360 ( .A(net209606), .Y(net209634) );
  NAND2X1 U26361 ( .A(net209923), .B(net209924), .Y(n48144) );
  NOR2X1 U26362 ( .A(net151712), .B(net151673), .Y(n11141) );
  OAI211X1 U26363 ( .A0(n11443), .A1(n10040), .B0(n10044), .C0(n10045), .Y(
        n11438) );
  AOI21X1 U26364 ( .A0(net210585), .A1(n47776), .B0(net210587), .Y(n11443) );
  NAND2X1 U26365 ( .A(n41357), .B(n47773), .Y(n47776) );
  CLKINVX1 U26366 ( .A(n11441), .Y(net151711) );
  AOI21X1 U26367 ( .A0(n47752), .A1(n47751), .B0(n47750), .Y(n11775) );
  NAND2X1 U26368 ( .A(n41365), .B(n47748), .Y(n47751) );
  NOR2BX1 U26369 ( .AN(n48335), .B(n48291), .Y(n47748) );
  NAND2X1 U26370 ( .A(n37233), .B(net258903), .Y(n41276) );
  AOI21X1 U26371 ( .A0(n10394), .A1(net171231), .B0(net209549), .Y(n48348) );
  OAI21XL U26372 ( .A0(net209333), .A1(n48438), .B0(net209335), .Y(n48442) );
  CLKINVX1 U26373 ( .A(n48137), .Y(n48140) );
  OR2X1 U26374 ( .A(net209513), .B(n48369), .Y(n41344) );
  AOI21X1 U26375 ( .A0(n48368), .A1(n11733), .B0(net209516), .Y(n48369) );
  OAI21XL U26376 ( .A0(net209517), .A1(n48367), .B0(n10423), .Y(n48368) );
  AO21X1 U26377 ( .A0(n48324), .A1(n48323), .B0(n48322), .Y(n41673) );
  OAI21XL U26378 ( .A0(n48318), .A1(n48317), .B0(n48316), .Y(n48323) );
  OA21XL U26379 ( .A0(net209570), .A1(n48333), .B0(net209572), .Y(n41674) );
  CLKINVX1 U26380 ( .A(net210460), .Y(net209642) );
  OAI21XL U26381 ( .A0(n48428), .A1(n48427), .B0(n48426), .Y(n48429) );
  OAI211X1 U26382 ( .A0(n11128), .A1(n11129), .B0(n40397), .C0(n11131), .Y(
        n11125) );
  NOR2X1 U26383 ( .A(n36948), .B(n37199), .Y(n11425) );
  CLKINVX1 U26384 ( .A(n12749), .Y(net171236) );
  CLKINVX1 U26385 ( .A(n12793), .Y(net171242) );
  CLKINVX1 U26386 ( .A(n11733), .Y(net171248) );
  OA21XL U26387 ( .A0(n48354), .A1(n48353), .B0(n48352), .Y(n41663) );
  CLKINVX1 U26388 ( .A(n13015), .Y(net171555) );
  AO21X1 U26389 ( .A0(n11425), .A1(n11426), .B0(net151601), .Y(n41226) );
  CLKINVX1 U26390 ( .A(n12794), .Y(net171188) );
  CLKINVX1 U26391 ( .A(n12736), .Y(net171191) );
  OAI2BB1X1 U26392 ( .A0N(n10606), .A1N(n41708), .B0(n10607), .Y(n48222) );
  AO21X1 U26393 ( .A0(n48221), .A1(n10553), .B0(net209821), .Y(n41708) );
  OAI21XL U26394 ( .A0(n39806), .A1(n48220), .B0(n10556), .Y(n48221) );
  OAI21XL U26395 ( .A0(net171423), .A1(n48499), .B0(n10854), .Y(n48500) );
  AOI21X1 U26396 ( .A0(n48498), .A1(n12316), .B0(net171421), .Y(n48499) );
  AOI21X1 U26397 ( .A0(n48483), .A1(net209253), .B0(net209254), .Y(n48484) );
  NAND2X1 U26398 ( .A(n41371), .B(n10869), .Y(n48483) );
  OR2X1 U26399 ( .A(net209255), .B(n48482), .Y(n41371) );
  OAI21XL U26400 ( .A0(n48473), .A1(n48472), .B0(n48471), .Y(n48479) );
  NAND4BBXL U26401 ( .AN(n48477), .BN(n48476), .C(n48475), .D(n48474), .Y(
        n48478) );
  AND2X2 U26402 ( .A(net209242), .B(n12316), .Y(n48491) );
  AOI21X1 U26403 ( .A0(n41776), .A1(n48123), .B0(net209958), .Y(n48240) );
  CLKINVX1 U26404 ( .A(n12960), .Y(net171554) );
  NAND4BBXL U26405 ( .AN(n48513), .BN(n48512), .C(n48511), .D(n48510), .Y(
        n48514) );
  AOI21X1 U26406 ( .A0(n48420), .A1(n11085), .B0(n48419), .Y(n48516) );
  OAI21XL U26407 ( .A0(n48509), .A1(n48508), .B0(n48507), .Y(n48515) );
  OAI211X1 U26408 ( .A0(n12054), .A1(n12055), .B0(n10608), .C0(n10606), .Y(
        n12051) );
  AOI211X1 U26409 ( .A0(n12056), .A1(n12057), .B0(net171257), .C0(n39806), .Y(
        n12054) );
  CLKINVX1 U26410 ( .A(n12150), .Y(net151741) );
  NOR2X1 U26411 ( .A(n39566), .B(net210494), .Y(n39567) );
  NOR2X1 U26412 ( .A(net210441), .B(n37509), .Y(n39566) );
  NOR3BXL U26413 ( .AN(net209894), .B(net210492), .C(n39792), .Y(n39791) );
  CLKINVX1 U26414 ( .A(net209898), .Y(n39792) );
  NOR2X1 U26415 ( .A(net210476), .B(net210475), .Y(n39705) );
  CLKINVX1 U26416 ( .A(n12297), .Y(net171441) );
  AOI21X1 U26417 ( .A0(n48250), .A1(net209778), .B0(net171124), .Y(n48251) );
  OAI21X1 U26418 ( .A0(net171125), .A1(n48249), .B0(n12005), .Y(n48250) );
  NOR2X1 U26419 ( .A(n39311), .B(n39570), .Y(n39569) );
  NAND2X1 U26420 ( .A(net209930), .B(n37469), .Y(n39570) );
  NOR2X1 U26421 ( .A(net210490), .B(n37511), .Y(n39311) );
  OAI21XL U26422 ( .A0(net210392), .A1(n39706), .B0(n40011), .Y(n39709) );
  NOR2X1 U26423 ( .A(n39707), .B(n39705), .Y(n39706) );
  CLKINVX1 U26424 ( .A(net210390), .Y(n40011) );
  NAND2X1 U26425 ( .A(n37126), .B(net209603), .Y(n39711) );
  CLKINVX1 U26426 ( .A(net210469), .Y(n39710) );
  NOR2X1 U26427 ( .A(net210550), .B(n39496), .Y(n39497) );
  NOR2X1 U26428 ( .A(net210553), .B(net210554), .Y(n39496) );
  NAND2X1 U26429 ( .A(net209344), .B(net209313), .Y(n39946) );
  NOR2X1 U26430 ( .A(n39641), .B(n39642), .Y(n39643) );
  NOR2X1 U26431 ( .A(n39640), .B(net211102), .Y(n39641) );
  NOR4X1 U26432 ( .A(net210522), .B(net210210), .C(net210205), .D(n39639), .Y(
        n39640) );
  NOR2X1 U26433 ( .A(net210525), .B(net210216), .Y(n39639) );
  NOR2X1 U26434 ( .A(net171538), .B(net171537), .Y(n11380) );
  AOI21X1 U26435 ( .A0(n48072), .A1(n48071), .B0(n48070), .Y(n48083) );
  OAI21XL U26436 ( .A0(net210100), .A1(n48077), .B0(n11387), .Y(n48082) );
  NAND2X1 U26437 ( .A(n10184), .B(n39304), .Y(n39793) );
  NAND2X1 U26438 ( .A(n40010), .B(n40024), .Y(n39572) );
  CLKINVX1 U26439 ( .A(net210444), .Y(n40010) );
  OAI21XL U26440 ( .A0(n39569), .A1(n39571), .B0(n40009), .Y(n40024) );
  CLKINVX1 U26441 ( .A(net210445), .Y(n40009) );
  AOI21X1 U26442 ( .A0(n39715), .A1(n37125), .B0(net210426), .Y(n39714) );
  OAI21XL U26443 ( .A0(n39708), .A1(n39840), .B0(net235251), .Y(n39715) );
  NAND4X1 U26444 ( .A(net209583), .B(net210670), .C(net210650), .D(net213687),
        .Y(n39840) );
  AOI21X1 U26445 ( .A0(n39709), .A1(n39710), .B0(n39711), .Y(n39708) );
  NOR2X1 U26446 ( .A(n39843), .B(n39841), .Y(n39842) );
  NAND2X1 U26447 ( .A(n10126), .B(n10128), .Y(n39841) );
  NAND2X1 U26448 ( .A(net209565), .B(net210460), .Y(n39843) );
  NOR2BX1 U26449 ( .AN(n10393), .B(n39844), .Y(n39845) );
  NAND2X1 U26450 ( .A(n10395), .B(n10394), .Y(n39844) );
  NAND2X1 U26451 ( .A(net209291), .B(n39948), .Y(n39947) );
  CLKINVX1 U26452 ( .A(net210539), .Y(n39948) );
  AOI21X1 U26453 ( .A0(n39499), .A1(n39500), .B0(n37514), .Y(n39498) );
  NOR2X1 U26454 ( .A(net210548), .B(n39945), .Y(n39500) );
  OAI21XL U26455 ( .A0(n39497), .A1(net210552), .B0(n37468), .Y(n39499) );
  NAND2BX1 U26456 ( .AN(net210416), .B(n40031), .Y(n39374) );
  OAI21XL U26457 ( .A0(n39643), .A1(net210520), .B0(n40008), .Y(n40030) );
  CLKINVX1 U26458 ( .A(net210516), .Y(n40008) );
  NAND2X1 U26459 ( .A(n39881), .B(net210848), .Y(n39375) );
  NOR2X1 U26460 ( .A(n39882), .B(n39883), .Y(n39881) );
  CLKINVX1 U26461 ( .A(n10045), .Y(n39882) );
  CLKINVX1 U26462 ( .A(n10044), .Y(n39883) );
  CLKINVX1 U26463 ( .A(n13017), .Y(n50102) );
  NOR2X1 U26464 ( .A(n39314), .B(n39315), .Y(n39313) );
  AOI21X1 U26465 ( .A0(n39572), .A1(net210435), .B0(n39573), .Y(n39314) );
  OR2X1 U26466 ( .A(n10182), .B(n39793), .Y(n39573) );
  NOR2X1 U26467 ( .A(n10572), .B(n10570), .Y(n39796) );
  NAND3X1 U26468 ( .A(n12749), .B(n12085), .C(n39795), .Y(n39794) );
  CLKINVX1 U26469 ( .A(n10577), .Y(n39795) );
  NAND2X1 U26470 ( .A(n10573), .B(n12793), .Y(n39797) );
  AOI21X1 U26471 ( .A0(n39717), .A1(n39718), .B0(n39719), .Y(n39716) );
  NAND2X1 U26472 ( .A(n39845), .B(n11770), .Y(n39719) );
  CLKINVX1 U26473 ( .A(n10419), .Y(n39718) );
  NAND4X1 U26474 ( .A(n10384), .B(n10383), .C(n10385), .D(n10387), .Y(n39721)
         );
  NOR3BXL U26475 ( .AN(n10381), .B(net209543), .C(n40393), .Y(n39846) );
  NOR2X1 U26476 ( .A(net210528), .B(n39421), .Y(n39501) );
  AOI21X1 U26477 ( .A0(n37513), .A1(n39422), .B0(n39423), .Y(n39421) );
  OR2X1 U26478 ( .A(net210561), .B(net210537), .Y(n39423) );
  NOR2X1 U26479 ( .A(net209302), .B(n39947), .Y(n39422) );
  NAND2X1 U26480 ( .A(n11149), .B(n10257), .Y(n39503) );
  OAI21XL U26481 ( .A0(n10729), .A1(n39373), .B0(n39888), .Y(n39645) );
  NOR2X1 U26482 ( .A(n39889), .B(net210140), .Y(n39888) );
  AOI21X1 U26483 ( .A0(n37018), .A1(n39374), .B0(n39375), .Y(n39373) );
  NAND3X1 U26484 ( .A(n10732), .B(n10734), .C(n10730), .Y(n39889) );
  NOR2X1 U26485 ( .A(n39893), .B(n39891), .Y(n39892) );
  CLKINVX1 U26486 ( .A(n10724), .Y(n39893) );
  NAND2X1 U26487 ( .A(n10726), .B(n10725), .Y(n39891) );
  AO21X1 U26488 ( .A0(n48260), .A1(n11984), .B0(net209760), .Y(n41770) );
  OAI21XL U26489 ( .A0(n39335), .A1(n48259), .B0(n12800), .Y(n48260) );
  AOI21X1 U26490 ( .A0(n48258), .A1(n11988), .B0(net209763), .Y(n48259) );
  AO21X1 U26491 ( .A0(n48103), .A1(n11334), .B0(net151444), .Y(n41691) );
  OAI2BB1X1 U26492 ( .A0N(n10754), .A1N(n41690), .B0(n10757), .Y(n48103) );
  AO21X1 U26493 ( .A0(n48102), .A1(n10755), .B0(net151481), .Y(n41690) );
  OAI21XL U26494 ( .A0(net210067), .A1(n48101), .B0(n12901), .Y(n48102) );
  NAND2X1 U26495 ( .A(n40005), .B(n39798), .Y(n39320) );
  NOR2X1 U26496 ( .A(n39799), .B(n39797), .Y(n39798) );
  OAI21XL U26497 ( .A0(n39794), .A1(n39313), .B0(n39796), .Y(n40005) );
  NAND2X1 U26498 ( .A(n10566), .B(n10567), .Y(n39799) );
  NAND2X1 U26499 ( .A(n10378), .B(n12535), .Y(n39848) );
  OAI21XL U26500 ( .A0(n39847), .A1(n39720), .B0(n40037), .Y(n39724) );
  CLKINVX1 U26501 ( .A(n10420), .Y(n40037) );
  CLKINVX1 U26502 ( .A(n39846), .Y(n39847) );
  NOR2X1 U26503 ( .A(n39721), .B(n39716), .Y(n39720) );
  NOR3BXL U26504 ( .AN(n10863), .B(n39957), .C(net171435), .Y(n39956) );
  NAND2X1 U26505 ( .A(n11131), .B(n11132), .Y(n39957) );
  NAND3X1 U26506 ( .A(n10872), .B(net209253), .C(n39952), .Y(n39954) );
  NOR2X1 U26507 ( .A(n39953), .B(net209255), .Y(n39952) );
  NOR3X1 U26508 ( .A(n39506), .B(n10877), .C(net209259), .Y(n39507) );
  NOR2X1 U26509 ( .A(n39505), .B(n39502), .Y(n39506) );
  NOR4X1 U26510 ( .A(n39501), .B(n39503), .C(n39504), .D(net210531), .Y(n39502) );
  CLKINVX1 U26511 ( .A(n11147), .Y(n39504) );
  NAND2X1 U26512 ( .A(n39958), .B(net151599), .Y(n39429) );
  NOR2X1 U26513 ( .A(net171486), .B(net171489), .Y(n39958) );
  CLKINVX1 U26514 ( .A(n9915), .Y(n40012) );
  NOR2X1 U26515 ( .A(n39895), .B(n39648), .Y(n39894) );
  AOI21X1 U26516 ( .A0(n37345), .A1(n39645), .B0(n39646), .Y(n39644) );
  NAND2X1 U26517 ( .A(n13015), .B(n12960), .Y(n39895) );
  NOR2X1 U26518 ( .A(net210238), .B(n39897), .Y(n39896) );
  CLKINVX1 U26519 ( .A(n10709), .Y(n39897) );
  AOI21X1 U26520 ( .A0(n48263), .A1(n10506), .B0(net209753), .Y(n48264) );
  OAI2BB1X2 U26521 ( .A0N(n11978), .A1N(n41770), .B0(n11979), .Y(n48261) );
  OAI2BB1X1 U26522 ( .A0N(n12896), .A1N(n41691), .B0(n12892), .Y(n48104) );
  NOR2X1 U26523 ( .A(n10177), .B(n39319), .Y(n39574) );
  AOI21X1 U26524 ( .A0(n39320), .A1(n39321), .B0(n39322), .Y(n39319) );
  NAND3BX1 U26525 ( .AN(n39801), .B(n12794), .C(n10559), .Y(n39322) );
  CLKINVX1 U26526 ( .A(n10564), .Y(n39321) );
  NAND2X1 U26527 ( .A(n10556), .B(n10553), .Y(n39805) );
  CLKINVX1 U26528 ( .A(n10606), .Y(n39807) );
  OAI21XL U26529 ( .A0(n39723), .A1(n10113), .B0(n40036), .Y(n39727) );
  CLKINVX1 U26530 ( .A(n10421), .Y(n40036) );
  AOI21X1 U26531 ( .A0(n39724), .A1(n39725), .B0(n10112), .Y(n39723) );
  NOR3X1 U26532 ( .A(n39848), .B(net171185), .C(net151308), .Y(n39725) );
  NOR2X1 U26533 ( .A(n10254), .B(n39426), .Y(n39508) );
  AOI21X1 U26534 ( .A0(n39427), .A1(n39428), .B0(n39429), .Y(n39426) );
  CLKINVX1 U26535 ( .A(n10865), .Y(n39428) );
  OAI21XL U26536 ( .A0(n39954), .A1(n39507), .B0(n39956), .Y(n39427) );
  NAND2X1 U26537 ( .A(n10855), .B(n10852), .Y(n39965) );
  AOI21X1 U26538 ( .A0(n39650), .A1(n39651), .B0(n39652), .Y(n39649) );
  CLKINVX1 U26539 ( .A(n10705), .Y(n39651) );
  NAND3X1 U26540 ( .A(n10708), .B(n39896), .C(n10706), .Y(n39652) );
  OAI21XL U26541 ( .A0(n9913), .A1(n37475), .B0(n40012), .Y(n39650) );
  NOR2X1 U26542 ( .A(n10702), .B(net171551), .Y(n39898) );
  NAND2X1 U26543 ( .A(n10751), .B(net211667), .Y(n39901) );
  CLKINVX1 U26544 ( .A(n40390), .Y(net171469) );
  OAI211X1 U26545 ( .A0(n11332), .A1(n11333), .B0(n11334), .C0(n11335), .Y(
        n11329) );
  CLKINVX1 U26546 ( .A(n13019), .Y(net151445) );
  NAND2X1 U26547 ( .A(n11968), .B(n11967), .Y(n40883) );
  AO21X1 U26548 ( .A0(n48108), .A1(n12887), .B0(n36943), .Y(n41692) );
  OAI21XL U26549 ( .A0(n39628), .A1(n48107), .B0(n11515), .Y(n48108) );
  CLKINVX1 U26550 ( .A(n11325), .Y(net210057) );
  AOI21X1 U26551 ( .A0(n39577), .A1(n39578), .B0(n39579), .Y(n39576) );
  NAND4BX1 U26552 ( .AN(n39807), .B(n10608), .C(n10607), .D(n12150), .Y(n39579) );
  NOR3X1 U26553 ( .A(n39805), .B(n39806), .C(net171257), .Y(n39578) );
  OAI21XL U26554 ( .A0(n39574), .A1(n40401), .B0(n37349), .Y(n39577) );
  CLKINVX1 U26555 ( .A(n10609), .Y(n40023) );
  NAND2X1 U26556 ( .A(n10544), .B(n10543), .Y(n39809) );
  OAI21XL U26557 ( .A0(n39726), .A1(n39730), .B0(n10355), .Y(n39736) );
  AOI21X1 U26558 ( .A0(n39727), .A1(n39728), .B0(n39729), .Y(n39726) );
  NAND4BX1 U26559 ( .AN(net209516), .B(n11733), .C(n10422), .D(n10423), .Y(
        n39729) );
  NOR3X1 U26560 ( .A(n39849), .B(net171249), .C(net209529), .Y(n39728) );
  OAI21XL U26561 ( .A0(n39509), .A1(n39510), .B0(n39964), .Y(n40017) );
  NOR2X1 U26562 ( .A(n39965), .B(n39963), .Y(n39964) );
  NOR2X1 U26563 ( .A(n39508), .B(n10253), .Y(n39509) );
  NAND2X1 U26564 ( .A(n10854), .B(n10853), .Y(n39963) );
  CLKINVX1 U26565 ( .A(n10842), .Y(n40016) );
  NAND2X1 U26566 ( .A(n10845), .B(n10843), .Y(n39970) );
  AOI21X1 U26567 ( .A0(n39655), .A1(n39656), .B0(n10699), .Y(n39654) );
  NOR2BX1 U26568 ( .AN(n39899), .B(n39901), .Y(n39655) );
  OAI21XL U26569 ( .A0(n39649), .A1(n39653), .B0(n39898), .Y(n39656) );
  NOR2X1 U26570 ( .A(n39900), .B(net151737), .Y(n39899) );
  OR2X1 U26571 ( .A(n37516), .B(net171111), .Y(n40945) );
  NAND2X1 U26572 ( .A(n11967), .B(n11968), .Y(n40970) );
  CLKINVX1 U26573 ( .A(n40388), .Y(net171103) );
  NAND4BBXL U26574 ( .AN(n40882), .BN(n40971), .C(n10503), .D(n40975), .Y(
        n40974) );
  NOR2X1 U26575 ( .A(net260277), .B(n40883), .Y(n40882) );
  NAND3BX1 U26576 ( .AN(n11969), .B(n11968), .C(n11967), .Y(n40975) );
  NAND3X1 U26577 ( .A(n11961), .B(net261020), .C(n11960), .Y(n40971) );
  CLKINVX1 U26578 ( .A(n40945), .Y(n40973) );
  CLKINVX1 U26579 ( .A(n11961), .Y(n_cell_301249_net269482) );
  NAND2X1 U26580 ( .A(net209746), .B(n11961), .Y(n40916) );
  CLKINVX1 U26581 ( .A(n11960), .Y(n_cell_301249_net269481) );
  NOR2X1 U26582 ( .A(n39555), .B(n39556), .Y(n40977) );
  OAI2BB1X1 U26583 ( .A0N(n11960), .A1N(n41771), .B0(n11961), .Y(n48268) );
  AO21X1 U26584 ( .A0(n48267), .A1(n10501), .B0(net209746), .Y(n41771) );
  NAND2X1 U26585 ( .A(n41258), .B(n10503), .Y(n48267) );
  OR2X1 U26586 ( .A(net171327), .B(n48266), .Y(n41258) );
  CLKINVX1 U26587 ( .A(net259649), .Y(n_cell_303546_net277470) );
  CLKINVX1 U26588 ( .A(net260527), .Y(n_cell_303546_net277469) );
  NOR2X1 U26589 ( .A(n10170), .B(n39581), .Y(n39584) );
  AOI21X1 U26590 ( .A0(n39582), .A1(n39583), .B0(n10169), .Y(n39581) );
  NOR2X1 U26591 ( .A(n10542), .B(n39809), .Y(n39583) );
  OAI21XL U26592 ( .A0(n39576), .A1(n39580), .B0(n40023), .Y(n39582) );
  NOR2X1 U26593 ( .A(net171210), .B(net171214), .Y(n39814) );
  CLKINVX1 U26594 ( .A(n10166), .Y(n39811) );
  CLKINVX1 U26595 ( .A(n10098), .Y(n39850) );
  OAI21XL U26596 ( .A0(n39734), .A1(n40403), .B0(n40035), .Y(n39739) );
  CLKINVX1 U26597 ( .A(n10102), .Y(n40035) );
  AOI21X1 U26598 ( .A0(n39735), .A1(n39736), .B0(n10105), .Y(n39734) );
  NOR2X1 U26599 ( .A(net171300), .B(n10357), .Y(n39735) );
  AOI21X1 U26600 ( .A0(n39512), .A1(n39513), .B0(n39511), .Y(n39431) );
  NOR2X1 U26601 ( .A(n39971), .B(n39970), .Y(n39513) );
  NAND2X1 U26602 ( .A(n40017), .B(n40016), .Y(n39512) );
  NAND2X1 U26603 ( .A(n10846), .B(n10847), .Y(n39971) );
  NAND2X1 U26604 ( .A(n39972), .B(n40398), .Y(n39432) );
  CLKINVX1 U26605 ( .A(n10839), .Y(n39972) );
  AOI21X1 U26606 ( .A0(n39660), .A1(n39661), .B0(n10026), .Y(n39659) );
  CLKINVX1 U26607 ( .A(n10028), .Y(n39661) );
  OAI21XL U26608 ( .A0(n39654), .A1(n39657), .B0(n40029), .Y(n39660) );
  CLKINVX1 U26609 ( .A(n10032), .Y(n40029) );
  OR2X1 U26610 ( .A(n10025), .B(net171548), .Y(n39904) );
  OR2X1 U26611 ( .A(net171535), .B(net238947), .Y(n40829) );
  NOR2X1 U26612 ( .A(net151426), .B(n37510), .Y(n41075) );
  NAND2X1 U26613 ( .A(n39345), .B(n11299), .Y(n40921) );
  NOR2X1 U26614 ( .A(n39676), .B(n39677), .Y(n41079) );
  NAND2X1 U26615 ( .A(n39345), .B(n11299), .Y(n40923) );
  NAND2X1 U26616 ( .A(n_cell_303546_net275956), .B(n11291), .Y(n41083) );
  AOI21X1 U26617 ( .A0(n40973), .A1(n37515), .B0(n40974), .Y(n40972) );
  NOR3X1 U26618 ( .A(n40978), .B(n40915), .C(n40914), .Y(n40979) );
  NAND3X1 U26619 ( .A(net260251), .B(n40977), .C(net260247), .Y(n40978) );
  NOR2X1 U26620 ( .A(n_cell_301249_net269481), .B(n40916), .Y(n40915) );
  NOR3X1 U26621 ( .A(n_cell_301249_net269481), .B(n_cell_301249_net269482),
        .C(n10501), .Y(n40914) );
  NOR2X1 U26622 ( .A(n_cell_301249_net269564), .B(net209736), .Y(n40985) );
  CLKINVX1 U26623 ( .A(n10485), .Y(n_cell_301249_net269564) );
  NAND2X1 U26624 ( .A(n40983), .B(n40981), .Y(n40982) );
  NOR2X1 U26625 ( .A(net171156), .B(net171160), .Y(n40981) );
  NAND3BX1 U26626 ( .AN(net260427), .B(net260251), .C(net260247), .Y(n40983)
         );
  CLKINVX1 U26627 ( .A(net260431), .Y(net171160) );
  NOR2X1 U26628 ( .A(net259747), .B(net151504), .Y(n40980) );
  CLKINVX1 U26629 ( .A(net260251), .Y(net151504) );
  NAND2X1 U26630 ( .A(n41634), .B(net259747), .Y(n48270) );
  OR2X1 U26631 ( .A(net171148), .B(n48269), .Y(n41634) );
  CLKINVX1 U26632 ( .A(net260427), .Y(net171148) );
  AOI21X1 U26633 ( .A0(n48268), .A1(n11958), .B0(n39555), .Y(n48269) );
  CLKINVX1 U26634 ( .A(n40389), .Y(net171156) );
  NOR2X1 U26635 ( .A(n40603), .B(n40601), .Y(n40602) );
  NAND2X1 U26636 ( .A(n_cell_303546_net275934), .B(n11613), .Y(n40601) );
  OAI21XL U26637 ( .A0(net260367), .A1(n_cell_303546_net277667), .B0(n40604),
        .Y(n40603) );
  AND2X2 U26638 ( .A(net259649), .B(net260527), .Y(n40604) );
  NAND2X1 U26639 ( .A(n39444), .B(net259641), .Y(n40600) );
  NOR4X1 U26640 ( .A(net151283), .B(n_cell_303546_net277470), .C(n11614), .D(
        n_cell_303546_net277469), .Y(n40570) );
  NOR3X1 U26641 ( .A(n_cell_303546_net277469), .B(n39470), .C(
        n_cell_303546_net277470), .Y(n40492) );
  NAND2X1 U26642 ( .A(net260900), .B(n40606), .Y(n40605) );
  NAND2BX1 U26643 ( .AN(net259653), .B(net260527), .Y(n40606) );
  NOR2X1 U26644 ( .A(n_cell_303546_net277632), .B(n_cell_303546_net277671),
        .Y(n40607) );
  CLKINVX1 U26645 ( .A(n11606), .Y(n_cell_303546_net277671) );
  CLKINVX1 U26646 ( .A(n40411), .Y(n40764) );
  CLKINVX1 U26647 ( .A(n11600), .Y(n_cell_303546_net277632) );
  OAI2BB1X1 U26648 ( .A0N(n12876), .A1N(n41693), .B0(n12872), .Y(n48113) );
  AO21X1 U26649 ( .A0(n48112), .A1(net210043), .B0(net238868), .Y(n41693) );
  NAND2X1 U26650 ( .A(n41204), .B(n12878), .Y(n48112) );
  OR2X1 U26651 ( .A(n36945), .B(n48111), .Y(n41204) );
  NAND2X1 U26652 ( .A(n10801), .B(n39532), .Y(n40542) );
  OAI21XL U26653 ( .A0(n39585), .A1(n39810), .B0(n39813), .Y(n39587) );
  NAND2X1 U26654 ( .A(n39811), .B(n40386), .Y(n39810) );
  NOR3BXL U26655 ( .AN(n39814), .B(n39815), .C(net171205), .Y(n39813) );
  NOR2X1 U26656 ( .A(n39584), .B(n40402), .Y(n39585) );
  CLKINVX1 U26657 ( .A(n10532), .Y(n39588) );
  OAI21XL U26658 ( .A0(n39737), .A1(n10097), .B0(n10091), .Y(n39744) );
  AOI21X1 U26659 ( .A0(n39738), .A1(n39739), .B0(n39740), .Y(n39737) );
  NOR2X1 U26660 ( .A(n10101), .B(net171198), .Y(n39738) );
  NAND2X1 U26661 ( .A(n39850), .B(n11688), .Y(n39740) );
  NOR2X1 U26662 ( .A(n10093), .B(n10094), .Y(n39743) );
  NOR2X1 U26663 ( .A(net151662), .B(net171456), .Y(n39973) );
  AOI21X1 U26664 ( .A0(n39515), .A1(n39516), .B0(n10240), .Y(n39514) );
  CLKINVX1 U26665 ( .A(n10242), .Y(n39516) );
  OAI21XL U26666 ( .A0(n10246), .A1(n39430), .B0(net168852), .Y(n39515) );
  NOR2X1 U26667 ( .A(n39431), .B(n39432), .Y(n39430) );
  AOI21X1 U26668 ( .A0(n39663), .A1(n39664), .B0(n10020), .Y(n39662) );
  CLKINVX1 U26669 ( .A(n10018), .Y(n39664) );
  OAI21XL U26670 ( .A0(n39659), .A1(n39904), .B0(n40028), .Y(n39663) );
  CLKINVX1 U26671 ( .A(n10024), .Y(n40028) );
  NOR2X1 U26672 ( .A(net151462), .B(n10686), .Y(n39905) );
  CLKINVX1 U26673 ( .A(n10754), .Y(n39907) );
  CLKINVX1 U26674 ( .A(n10757), .Y(n39906) );
  NAND2X1 U26675 ( .A(n41229), .B(n41230), .Y(n44148) );
  NAND2X1 U26676 ( .A(n41260), .B(n41261), .Y(n44048) );
  CLKINVX1 U26677 ( .A(net219450), .Y(net258961) );
  XOR2X1 U26678 ( .A(n41829), .B(n42605), .Y(n44643) );
  NAND2X1 U26679 ( .A(n10904), .B(n10992), .Y(n41142) );
  NAND2X1 U26680 ( .A(n10904), .B(n_cell_301249_net269794), .Y(n40925) );
  CLKINVX1 U26681 ( .A(n10990), .Y(n_cell_301249_net269794) );
  OAI21XL U26682 ( .A0(n11308), .A1(n41074), .B0(n41075), .Y(n40831) );
  OR2X1 U26683 ( .A(net171535), .B(net238947), .Y(n41074) );
  OAI21XL U26684 ( .A0(n10010), .A1(net259841), .B0(n41077), .Y(n40833) );
  NOR2X1 U26685 ( .A(n_cell_301249_net269688), .B(n41076), .Y(n41077) );
  CLKINVX1 U26686 ( .A(n12873), .Y(n_cell_301249_net269688) );
  NAND3X1 U26687 ( .A(n39345), .B(net260488), .C(n11299), .Y(n41076) );
  NOR3X1 U26688 ( .A(n41078), .B(n40922), .C(n40920), .Y(n41080) );
  NOR2X1 U26689 ( .A(n11300), .B(n40923), .Y(n40922) );
  NAND2X1 U26690 ( .A(n11519), .B(n41079), .Y(n41078) );
  NOR2X1 U26691 ( .A(n11301), .B(n40921), .Y(n40920) );
  NOR2X1 U26692 ( .A(n41084), .B(n41086), .Y(n41085) );
  OAI22XL U26693 ( .A0(n13022), .A1(n41082), .B0(n12867), .B1(n41083), .Y(
        n41086) );
  NAND2X1 U26694 ( .A(n_cell_303546_net276009), .B(net260492), .Y(n41084) );
  NAND2X1 U26695 ( .A(n_cell_303546_net275956), .B(n11291), .Y(n41082) );
  NOR2X1 U26696 ( .A(n39623), .B(n_cell_303546_net277530), .Y(n41091) );
  NAND2X1 U26697 ( .A(n39919), .B(net260492), .Y(n41090) );
  NAND2X1 U26698 ( .A(n11625), .B(n11626), .Y(n40859) );
  NAND2X1 U26699 ( .A(n11626), .B(n11625), .Y(n41019) );
  NOR3BXL U26700 ( .AN(net259645), .B(n_cell_301249_net269613), .C(n41020),
        .Y(n41021) );
  CLKINVX1 U26701 ( .A(n11621), .Y(n_cell_301249_net269613) );
  NAND2X1 U26702 ( .A(net259641), .B(n11622), .Y(n41020) );
  NAND4X1 U26703 ( .A(n39444), .B(n_cell_303546_net275934), .C(n39470), .D(
        net260367), .Y(n41023) );
  CLKINVX1 U26704 ( .A(n10425), .Y(n_cell_301249_net269950) );
  NOR2X1 U26705 ( .A(n_cell_301249_net269488), .B(net171169), .Y(n41025) );
  NAND3BX1 U26706 ( .AN(n11614), .B(n39470), .C(n_cell_303546_net275934), .Y(
        n41028) );
  NAND2X1 U26707 ( .A(n40411), .B(n40415), .Y(n40929) );
  AOI21X1 U26708 ( .A0(n40980), .A1(net260247), .B0(n40982), .Y(n40886) );
  NAND2X1 U26709 ( .A(n10481), .B(n40985), .Y(n40887) );
  NAND2X1 U26710 ( .A(n40979), .B(n41194), .Y(n40885) );
  OAI21XL U26711 ( .A0(n37347), .A1(n_cell_301249_net269449), .B0(n40987), .Y(
        n40889) );
  NOR3BXL U26712 ( .AN(n12640), .B(n_cell_301249_net269568), .C(n40986), .Y(
        n40987) );
  NAND2X1 U26713 ( .A(n_cell_303546_net275967), .B(n_cell_303546_net275987),
        .Y(n40986) );
  NOR2X1 U26714 ( .A(n40936), .B(n40934), .Y(n40996) );
  NOR2X1 U26715 ( .A(net260412), .B(n40935), .Y(n40934) );
  NOR3BXL U26716 ( .AN(n11934), .B(n12804), .C(n39554), .Y(n40936) );
  NAND2X1 U26717 ( .A(n11934), .B(n11935), .Y(n40935) );
  NAND2X1 U26718 ( .A(n_cell_303546_net276178), .B(n40995), .Y(n40994) );
  NOR2X1 U26719 ( .A(n_cell_301249_net269578), .B(n39552), .Y(n40995) );
  NOR2X1 U26720 ( .A(n39554), .B(n_cell_301249_net269571), .Y(n40989) );
  NAND3X1 U26721 ( .A(n39605), .B(n_cell_303546_net275967), .C(
        n_cell_303546_net275987), .Y(n40993) );
  NAND3X1 U26722 ( .A(n_cell_303546_net275987), .B(n_cell_303546_net275967),
        .C(n_cell_301249_net269969), .Y(n40992) );
  CLKINVX1 U26723 ( .A(n11943), .Y(n_cell_301249_net269969) );
  NAND2X1 U26724 ( .A(n10480), .B(n12165), .Y(n40990) );
  NAND2X1 U26725 ( .A(n_cell_303546_net276178), .B(n_cell_303546_net277942),
        .Y(n40942) );
  NAND2X1 U26726 ( .A(n_cell_303546_net276178), .B(n_cell_301249_net269583),
        .Y(n40944) );
  CLKINVX1 U26727 ( .A(net271999), .Y(net171175) );
  NAND2BX1 U26728 ( .AN(net209733), .B(n12803), .Y(n40468) );
  NOR2X1 U26729 ( .A(n40465), .B(n40723), .Y(n40724) );
  NAND2X1 U26730 ( .A(n11943), .B(n_cell_303546_net275967), .Y(n40723) );
  NOR2X1 U26731 ( .A(net209733), .B(n40466), .Y(n40465) );
  NAND2BX1 U26732 ( .AN(n12643), .B(n12803), .Y(n40466) );
  NAND2X1 U26733 ( .A(n40726), .B(n12804), .Y(n40727) );
  NOR2X1 U26734 ( .A(n_cell_303546_net277834), .B(n_cell_303546_net277630),
        .Y(n40726) );
  AOI21X1 U26735 ( .A0(n40494), .A1(n40495), .B0(n40496), .Y(n40493) );
  OAI21XL U26736 ( .A0(net171169), .A1(n11607), .B0(n40607), .Y(n40496) );
  NOR4X1 U26737 ( .A(n40570), .B(n40605), .C(net171169), .D(n40492), .Y(n40495) );
  OAI21XL U26738 ( .A0(net209446), .A1(n40600), .B0(n40602), .Y(n40494) );
  AND3X2 U26739 ( .A(n40611), .B(n40612), .C(n40609), .Y(n40610) );
  NAND2BX1 U26740 ( .AN(n12433), .B(net260376), .Y(n40612) );
  NOR2BX1 U26741 ( .AN(n40418), .B(n_cell_301249_net269943), .Y(n40609) );
  NAND3X1 U26742 ( .A(net260376), .B(n40415), .C(n40764), .Y(n40611) );
  NAND4BX1 U26743 ( .AN(n40576), .B(n40415), .C(net260376), .D(n11601), .Y(
        n40608) );
  NOR2X1 U26744 ( .A(n_cell_303546_net277632), .B(n11605), .Y(n40576) );
  NAND2BX1 U26745 ( .AN(n40613), .B(n40615), .Y(n40614) );
  NAND2X1 U26746 ( .A(n10302), .B(n40422), .Y(n40613) );
  NAND2X1 U26747 ( .A(n_cell_301249_net269941), .B(n40418), .Y(n40615) );
  NOR2X1 U26748 ( .A(net171315), .B(n40618), .Y(n40617) );
  CLKINVX1 U26749 ( .A(n12427), .Y(n40618) );
  NAND2X1 U26750 ( .A(n40616), .B(net261422), .Y(n40619) );
  NOR2BX1 U26751 ( .AN(n10302), .B(n11869), .Y(n40616) );
  NAND2X1 U26752 ( .A(net261422), .B(n_cell_303546_net277892), .Y(n40620) );
  CLKINVX1 U26753 ( .A(net259626), .Y(n_cell_303546_net277892) );
  OAI21XL U26754 ( .A0(n13022), .A1(n39677), .B0(n40688), .Y(n40689) );
  NOR2X1 U26755 ( .A(n_cell_303546_net277772), .B(n39676), .Y(n40688) );
  NOR2X1 U26756 ( .A(n10662), .B(n40518), .Y(n40517) );
  NAND2X1 U26757 ( .A(n_cell_303546_net275956), .B(n12867), .Y(n40518) );
  OR3X2 U26758 ( .A(net171480), .B(net151532), .C(net171398), .Y(n40641) );
  NOR3X1 U26759 ( .A(n40541), .B(n40642), .C(n40543), .Y(n40643) );
  NAND2X1 U26760 ( .A(n10983), .B(n_cell_303546_net275923), .Y(n40642) );
  NOR2X1 U26761 ( .A(n10905), .B(net171398), .Y(n40543) );
  NOR2X1 U26762 ( .A(net171398), .B(n40542), .Y(n40541) );
  OAI21XL U26763 ( .A0(n_cell_301249_net269797), .A1(n_cell_303546_net275959),
        .B0(net260332), .Y(n40646) );
  CLKINVX1 U26764 ( .A(n10965), .Y(n40574) );
  NAND2BX1 U26765 ( .AN(net259873), .B(n_cell_303546_net275998), .Y(n40648) );
  NAND2X1 U26766 ( .A(n10519), .B(n10520), .Y(n39819) );
  OAI21XL U26767 ( .A0(n39591), .A1(n39592), .B0(n39816), .Y(n39332) );
  NOR2X1 U26768 ( .A(net171139), .B(n10152), .Y(n39816) );
  NOR2X1 U26769 ( .A(n39586), .B(n39589), .Y(n39591) );
  AOI21X1 U26770 ( .A0(n39587), .A1(n39588), .B0(n10155), .Y(n39586) );
  NAND2X1 U26771 ( .A(n39820), .B(net151456), .Y(n39334) );
  NOR2X1 U26772 ( .A(net171117), .B(net209768), .Y(n39820) );
  NAND2X1 U26773 ( .A(n10339), .B(n10336), .Y(n39853) );
  NAND2X1 U26774 ( .A(n10340), .B(n10341), .Y(n39854) );
  OAI21XL U26775 ( .A0(n39742), .A1(n39852), .B0(n37470), .Y(n39748) );
  OR2X1 U26776 ( .A(n10086), .B(n39851), .Y(n39852) );
  AOI21X1 U26777 ( .A0(n39743), .A1(n39744), .B0(n10085), .Y(n39742) );
  NAND2X1 U26778 ( .A(n10089), .B(n10090), .Y(n39851) );
  AOI21X1 U26779 ( .A0(n39519), .A1(net151652), .B0(n39517), .Y(n39518) );
  OAI21XL U26780 ( .A0(n39514), .A1(n39974), .B0(n40015), .Y(n39519) );
  NAND3X1 U26781 ( .A(n10243), .B(n10827), .C(n39973), .Y(n39974) );
  CLKINVX1 U26782 ( .A(n10829), .Y(n40015) );
  NOR2X1 U26783 ( .A(n10231), .B(n39978), .Y(n39977) );
  NAND2X1 U26784 ( .A(n10233), .B(n10232), .Y(n39978) );
  NOR2X1 U26785 ( .A(n39667), .B(n39670), .Y(n39671) );
  AOI21X1 U26786 ( .A0(n39668), .A1(n39669), .B0(n39666), .Y(n39667) );
  NOR4X1 U26787 ( .A(net151481), .B(n39906), .C(n39907), .D(n39908), .Y(n39668) );
  OAI21XL U26788 ( .A0(n39662), .A1(n39665), .B0(n39905), .Y(n39669) );
  XOR2X1 U26789 ( .A(n41812), .B(n42515), .Y(n44940) );
  NAND2X1 U26790 ( .A(n41350), .B(n41351), .Y(n44941) );
  XOR2X1 U26791 ( .A(n42070), .B(n41323), .Y(n44945) );
  XOR2X1 U26792 ( .A(n42090), .B(n41321), .Y(n44756) );
  NAND2X1 U26793 ( .A(n41231), .B(net219468), .Y(n41233) );
  XOR2X1 U26794 ( .A(n41842), .B(n42609), .Y(n27722) );
  OR2X1 U26795 ( .A(n41773), .B(n26750), .Y(n44287) );
  OR2X1 U26796 ( .A(n26757), .B(n26765), .Y(n41773) );
  CLKINVX1 U26797 ( .A(n26755), .Y(n44296) );
  NAND4BBXL U26798 ( .AN(n26745), .BN(n26756), .C(n37210), .D(n44294), .Y(
        n44299) );
  NOR3X1 U26799 ( .A(n26749), .B(n26766), .C(n44293), .Y(n44294) );
  NOR2X1 U26800 ( .A(n26767), .B(n44289), .Y(n44291) );
  CLKINVX1 U26801 ( .A(n26759), .Y(n44290) );
  XOR2X1 U26802 ( .A(n41799), .B(n36867), .Y(n43890) );
  NOR4X1 U26803 ( .A(n43897), .B(n43896), .C(n43895), .D(n43894), .Y(n43903)
         );
  OR4X1 U26804 ( .A(n44013), .B(n44012), .C(n44011), .D(n44010), .Y(n41684) );
  XNOR2X1 U26805 ( .A(n50377), .B(n42711), .Y(n28031) );
  XOR2X1 U26806 ( .A(n42698), .B(n41799), .Y(n43867) );
  XOR2X1 U26807 ( .A(n42709), .B(n42063), .Y(n43869) );
  NOR2X1 U26808 ( .A(n44939), .B(n44938), .Y(n46505) );
  NAND4X1 U26809 ( .A(n44933), .B(n44932), .C(n44931), .D(n44930), .Y(n44939)
         );
  NAND4X1 U26810 ( .A(n44937), .B(n44936), .C(n44935), .D(n44934), .Y(n44938)
         );
  CLKINVX1 U26811 ( .A(n47727), .Y(n48306) );
  NOR2X1 U26812 ( .A(n46489), .B(n48151), .Y(n46499) );
  NOR2X1 U26813 ( .A(n46511), .B(n48156), .Y(n46521) );
  XOR2X1 U26814 ( .A(n41821), .B(n42597), .Y(n45348) );
  NOR4X1 U26815 ( .A(n45354), .B(n45353), .C(n45352), .D(n45351), .Y(n45365)
         );
  XOR2X1 U26816 ( .A(n41821), .B(n36894), .Y(n45298) );
  NOR4X1 U26817 ( .A(n45296), .B(n45295), .C(n45294), .D(n45293), .Y(n45307)
         );
  NOR4X1 U26818 ( .A(n45385), .B(n45384), .C(n45383), .D(n45382), .Y(n45396)
         );
  NAND4X1 U26819 ( .A(n44752), .B(n44751), .C(n44750), .D(n44749), .Y(n48326)
         );
  NOR4X1 U26820 ( .A(n44748), .B(n44747), .C(n44746), .D(n44745), .Y(n44749)
         );
  NAND4X1 U26821 ( .A(n44721), .B(n44720), .C(n44719), .D(n44718), .Y(n48320)
         );
  NOR4BBX1 U26822 ( .AN(n41720), .BN(n41721), .C(n44717), .D(n44716), .Y(
        n44718) );
  NOR4X1 U26823 ( .A(n44707), .B(n44706), .C(n44705), .D(n44704), .Y(n44721)
         );
  OAI21XL U26824 ( .A0(n10993), .A1(n37179), .B0(n41143), .Y(n40807) );
  NOR3BXL U26825 ( .AN(n10991), .B(net171480), .C(n41142), .Y(n41143) );
  NOR4X1 U26826 ( .A(net151532), .B(n_cell_301249_net269797), .C(
        n_cell_301249_net269798), .D(n39991), .Y(n41146) );
  CLKINVX1 U26827 ( .A(n_cell_303546_net275959), .Y(n_cell_301249_net269798)
         );
  NOR2X1 U26828 ( .A(n40926), .B(n40924), .Y(n41147) );
  NOR2X1 U26829 ( .A(n10903), .B(n40927), .Y(n40926) );
  NOR2X1 U26830 ( .A(net171480), .B(n40925), .Y(n40924) );
  NAND2X1 U26831 ( .A(n10904), .B(n10906), .Y(n40927) );
  OAI21X1 U26832 ( .A0(n10983), .A1(n41150), .B0(n41154), .Y(n41153) );
  NAND2X1 U26833 ( .A(n_cell_303546_net275959), .B(n_cell_303546_net275923),
        .Y(n41150) );
  NAND3X1 U26834 ( .A(n_cell_303546_net275959), .B(n_cell_303546_net275923),
        .C(net171398), .Y(n41154) );
  NAND2X1 U26835 ( .A(n_cell_303546_net275998), .B(n10976), .Y(n41152) );
  CLKINVX1 U26836 ( .A(net271956), .Y(net171396) );
  NOR2X1 U26837 ( .A(n39483), .B(n_cell_301249_net269811), .Y(n41156) );
  CLKINVX1 U26838 ( .A(n10973), .Y(n_cell_301249_net269811) );
  NAND3BX1 U26839 ( .AN(net259873), .B(n10976), .C(n_cell_303546_net275998),
        .Y(n41158) );
  NOR2X1 U26840 ( .A(n41092), .B(n40932), .Y(n40836) );
  NOR2X1 U26841 ( .A(n11520), .B(n40933), .Y(n40932) );
  OAI21XL U26842 ( .A0(n_cell_301249_net269711), .A1(n41090), .B0(n41091), .Y(
        n41092) );
  NAND2X1 U26843 ( .A(n_cell_303546_net276009), .B(net260492), .Y(n40933) );
  NAND3X1 U26844 ( .A(n11280), .B(net260494), .C(n41093), .Y(n40837) );
  NOR2X1 U26845 ( .A(net171525), .B(n_cell_301249_net269714), .Y(n41093) );
  NAND3X1 U26846 ( .A(n41095), .B(net260470), .C(n11273), .Y(n41096) );
  NOR2X1 U26847 ( .A(net151554), .B(n39621), .Y(n41095) );
  NOR2X1 U26848 ( .A(net151539), .B(n_cell_301249_net269714), .Y(n41094) );
  NOR2X1 U26849 ( .A(net151555), .B(n40940), .Y(n40939) );
  NAND2X1 U26850 ( .A(n39923), .B(net260474), .Y(n40940) );
  OAI21XL U26851 ( .A0(net151555), .A1(n41098), .B0(n41099), .Y(n41101) );
  NAND2X1 U26852 ( .A(net151550), .B(net260474), .Y(n41098) );
  NOR2X1 U26853 ( .A(net151558), .B(n_cell_303546_net277536), .Y(n41099) );
  CLKINVX1 U26854 ( .A(n13025), .Y(net151558) );
  NOR3X1 U26855 ( .A(n41023), .B(n37528), .C(n37181), .Y(n41024) );
  OAI21XL U26856 ( .A0(n_cell_301249_net269615), .A1(n41019), .B0(n41021), .Y(
        n41022) );
  NOR2X1 U26857 ( .A(n41026), .B(n41027), .Y(n41030) );
  NAND2X1 U26858 ( .A(n41028), .B(n41029), .Y(n41027) );
  NAND3X1 U26859 ( .A(net259653), .B(net259649), .C(n41025), .Y(n41026) );
  NAND3X1 U26860 ( .A(n_cell_303546_net275934), .B(n39470), .C(net171158), .Y(
        n41029) );
  NOR2X1 U26861 ( .A(n40930), .B(n40928), .Y(n41033) );
  NOR2X1 U26862 ( .A(n11601), .B(n40931), .Y(n40930) );
  NOR2X1 U26863 ( .A(n11600), .B(n40929), .Y(n40928) );
  NAND2X1 U26864 ( .A(n40411), .B(n40415), .Y(n40931) );
  AND2X2 U26865 ( .A(net260376), .B(n12433), .Y(n41032) );
  NOR3X1 U26866 ( .A(net260527), .B(n_cell_301249_net269488), .C(net171169),
        .Y(n40919) );
  NAND4X1 U26867 ( .A(n11605), .B(n11606), .C(n40411), .D(n40415), .Y(n41031)
         );
  NOR2X1 U26868 ( .A(net260900), .B(n40918), .Y(n40917) );
  NAND2X1 U26869 ( .A(n10319), .B(n11607), .Y(n40918) );
  NAND4BX1 U26870 ( .AN(n40990), .B(n40989), .C(n40992), .D(n40993), .Y(n40991) );
  NOR3BXL U26871 ( .AN(n40996), .B(n40994), .C(net171175), .Y(n40997) );
  NOR3X1 U26872 ( .A(n40943), .B(n40941), .C(n40998), .Y(n40892) );
  NAND2X1 U26873 ( .A(n11924), .B(n11925), .Y(n40998) );
  NOR2X1 U26874 ( .A(net171175), .B(n40944), .Y(n40943) );
  NOR2X1 U26875 ( .A(net171175), .B(n40942), .Y(n40941) );
  NAND2X1 U26876 ( .A(n10469), .B(n10471), .Y(n40893) );
  CLKINVX1 U26877 ( .A(n12806), .Y(n_cell_301249_net269590) );
  NOR3X1 U26878 ( .A(n40575), .B(n40469), .C(n40729), .Y(n40730) );
  NAND2X1 U26879 ( .A(n11935), .B(n11932), .Y(n40729) );
  NOR2X1 U26880 ( .A(net260412), .B(n39553), .Y(n40469) );
  NOR3BXL U26881 ( .AN(net151542), .B(n39553), .C(n_cell_303546_net277630),
        .Y(n40575) );
  NAND2X1 U26882 ( .A(n_cell_303546_net277942), .B(n12166), .Y(n40732) );
  CLKINVX1 U26883 ( .A(n11924), .Y(n_cell_303546_net277843) );
  NAND2X1 U26884 ( .A(n_cell_301249_net269571), .B(n11932), .Y(n40731) );
  AOI21X1 U26885 ( .A0(n40498), .A1(n40499), .B0(n40500), .Y(n40497) );
  NAND3X1 U26886 ( .A(n40619), .B(n40620), .C(n40617), .Y(n40500) );
  NOR2X1 U26887 ( .A(n40614), .B(net171318), .Y(n40498) );
  OAI21XL U26888 ( .A0(net171315), .A1(n12424), .B0(n40621), .Y(n40622) );
  NOR2BX1 U26889 ( .AN(n10433), .B(n_cell_301249_net269635), .Y(n40621) );
  AOI21X1 U26890 ( .A0(net151304), .A1(n10433), .B0(n40623), .Y(n40624) );
  NAND2X1 U26891 ( .A(n_cell_303546_net276365), .B(net259661), .Y(n40623) );
  NAND2X1 U26892 ( .A(n11578), .B(n11576), .Y(n40625) );
  NOR3BXL U26893 ( .AN(net260352), .B(n11575), .C(n39701), .Y(n40581) );
  NOR3BXL U26894 ( .AN(n40691), .B(n39919), .C(n_cell_301249_net269711), .Y(
        n40521) );
  AOI21X1 U26895 ( .A0(n_cell_301249_net269701), .A1(n10659), .B0(
        n_cell_303546_net277530), .Y(n40691) );
  OAI21XL U26896 ( .A0(n11520), .A1(n40692), .B0(n40693), .Y(n40523) );
  NOR3BXL U26897 ( .AN(n11283), .B(n40519), .C(net171524), .Y(n40693) );
  NAND2X1 U26898 ( .A(n_cell_303546_net276009), .B(n11282), .Y(n40692) );
  NOR2X1 U26899 ( .A(net260492), .B(n_cell_303546_net277530), .Y(n40519) );
  OAI21XL U26900 ( .A0(n_cell_301249_net269714), .A1(n12855), .B0(n11274), .Y(
        n40696) );
  CLKINVX1 U26901 ( .A(net260494), .Y(net151539) );
  CLKINVX1 U26902 ( .A(n12848), .Y(n_cell_303546_net277536) );
  NOR2X1 U26903 ( .A(n40574), .B(n10969), .Y(n40573) );
  CLKINVX1 U26904 ( .A(n10966), .Y(n40652) );
  NAND2X1 U26905 ( .A(n40770), .B(n40645), .Y(n40545) );
  NOR2X1 U26906 ( .A(n40646), .B(n40644), .Y(n40645) );
  OAI21XL U26907 ( .A0(n40641), .A1(net209142), .B0(n40643), .Y(n40770) );
  NAND2X1 U26908 ( .A(n_cell_303546_net275998), .B(net271956), .Y(n40644) );
  OAI2BB1X1 U26909 ( .A0N(n39483), .A1N(n10973), .B0(n40649), .Y(n40547) );
  NOR2X1 U26910 ( .A(n40574), .B(n40650), .Y(n40649) );
  CLKINVX1 U26911 ( .A(n10968), .Y(n40650) );
  NOR2X1 U26912 ( .A(n40647), .B(n40571), .Y(n40546) );
  NOR2X1 U26913 ( .A(net209136), .B(n40572), .Y(n40571) );
  NAND3X1 U26914 ( .A(n10976), .B(n10973), .C(n40648), .Y(n40647) );
  NAND2X1 U26915 ( .A(net260332), .B(n_cell_303546_net275998), .Y(n40572) );
  NAND2X1 U26916 ( .A(n10503), .B(n10502), .Y(n39824) );
  OAI21XL U26917 ( .A0(n39331), .A1(n10512), .B0(n40025), .Y(n39594) );
  CLKINVX1 U26918 ( .A(n10509), .Y(n40025) );
  AOI21X1 U26919 ( .A0(n39332), .A1(n39333), .B0(n39334), .Y(n39331) );
  NOR2X1 U26920 ( .A(n10522), .B(n39819), .Y(n39333) );
  NAND3X1 U26921 ( .A(n10506), .B(n40388), .C(n39822), .Y(n39595) );
  NOR2BX1 U26922 ( .AN(n10504), .B(net171105), .Y(n39822) );
  OAI21XL U26923 ( .A0(n39747), .A1(n10334), .B0(n40007), .Y(n39754) );
  CLKINVX1 U26924 ( .A(n10082), .Y(n40007) );
  AOI21X1 U26925 ( .A0(n39748), .A1(n39749), .B0(n10338), .Y(n39747) );
  NOR2X1 U26926 ( .A(n39854), .B(n39853), .Y(n39749) );
  NAND2X1 U26927 ( .A(n39979), .B(n40006), .Y(n39523) );
  NOR2X1 U26928 ( .A(n10821), .B(n39980), .Y(n39979) );
  OAI21XL U26929 ( .A0(n10230), .A1(n39518), .B0(n39977), .Y(n40006) );
  CLKINVX1 U26930 ( .A(n10820), .Y(n39980) );
  NOR2X1 U26931 ( .A(n10819), .B(n39981), .Y(n39524) );
  NAND2X1 U26932 ( .A(n40390), .B(n11034), .Y(n39981) );
  CLKINVX1 U26933 ( .A(n10657), .Y(n39919) );
  CLKINVX1 U26934 ( .A(n39345), .Y(n39917) );
  CLKINVX1 U26935 ( .A(n11299), .Y(net151514) );
  OAI21XL U26936 ( .A0(n10671), .A1(n39672), .B0(n39910), .Y(n39674) );
  NOR3BXL U26937 ( .AN(n10672), .B(n39911), .C(net171533), .Y(n39910) );
  NOR2X1 U26938 ( .A(n39671), .B(n10679), .Y(n39672) );
  NAND2X1 U26939 ( .A(n40405), .B(n11315), .Y(n39911) );
  OR2X1 U26940 ( .A(n_cell_301249_net269861), .B(net259841), .Y(n39675) );
  NOR2X1 U26941 ( .A(n12326), .B(n47218), .Y(n47222) );
  NOR2X1 U26942 ( .A(n10869), .B(n47887), .Y(n47891) );
  OR2X1 U26943 ( .A(n29147), .B(n29139), .Y(n41754) );
  NOR4X1 U26944 ( .A(n45499), .B(n45498), .C(n45497), .D(n45496), .Y(n45510)
         );
  XOR2X1 U26945 ( .A(n42078), .B(n42665), .Y(n45497) );
  XOR2X1 U26946 ( .A(n41821), .B(n42523), .Y(n45398) );
  XOR2X1 U26947 ( .A(n42081), .B(n41322), .Y(n45370) );
  NOR2X1 U26948 ( .A(n12270), .B(n47917), .Y(n47921) );
  CLKINVX1 U26949 ( .A(net210695), .Y(net209899) );
  NAND4X1 U26950 ( .A(n45288), .B(n45287), .C(n45286), .D(n45285), .Y(n46573)
         );
  NOR2X1 U26951 ( .A(n45278), .B(n45277), .Y(n45288) );
  NOR2X1 U26952 ( .A(n45284), .B(n45283), .Y(n45285) );
  XOR2X1 U26953 ( .A(n42073), .B(n41321), .Y(n45129) );
  XOR2X1 U26954 ( .A(n41807), .B(n42529), .Y(n44995) );
  CLKINVX1 U26955 ( .A(net213679), .Y(net209624) );
  NOR2BX1 U26956 ( .AN(n41765), .B(n41710), .Y(n45052) );
  NOR2X1 U26957 ( .A(n45046), .B(n45045), .Y(n45054) );
  NAND2X1 U26958 ( .A(n41223), .B(n41224), .Y(n44821) );
  NOR4X1 U26959 ( .A(n44848), .B(n44847), .C(n44846), .D(n44845), .Y(n44849)
         );
  NAND4X2 U26960 ( .A(n44672), .B(n44671), .C(n44670), .D(n44669), .Y(n48175)
         );
  NOR4X1 U26961 ( .A(n44668), .B(n44667), .C(n44666), .D(n44665), .Y(n44669)
         );
  NOR2X1 U26962 ( .A(n44662), .B(n48325), .Y(n44672) );
  NOR2X1 U26963 ( .A(n44122), .B(net209595), .Y(n44132) );
  NOR2X1 U26964 ( .A(n44091), .B(net210643), .Y(n44101) );
  NOR2X1 U26965 ( .A(n43937), .B(net209572), .Y(n43947) );
  NOR4X1 U26966 ( .A(n28012), .B(n28011), .C(n28010), .D(n28009), .Y(n43821)
         );
  NOR4X1 U26967 ( .A(n26673), .B(n26674), .C(n26675), .D(n26676), .Y(n44304)
         );
  NOR2X1 U26968 ( .A(n44238), .B(n48370), .Y(n44242) );
  NOR2X1 U26969 ( .A(n11718), .B(n44521), .Y(n44525) );
  XOR2X1 U26970 ( .A(n42070), .B(n36888), .Y(n45150) );
  NAND2X1 U26971 ( .A(n41271), .B(n41272), .Y(n45149) );
  NAND2X1 U26972 ( .A(n41270), .B(n41385), .Y(n41272) );
  XOR2X1 U26973 ( .A(n41813), .B(n42611), .Y(n45138) );
  NAND2X1 U26974 ( .A(n41639), .B(n41640), .Y(n45109) );
  NAND2BX1 U26975 ( .AN(n41348), .B(n36919), .Y(n41639) );
  XOR2X1 U26976 ( .A(n42072), .B(n42660), .Y(n45113) );
  NAND2X1 U26977 ( .A(n41377), .B(n41378), .Y(n45202) );
  NAND2X1 U26978 ( .A(n42073), .B(n41376), .Y(n41377) );
  NOR4X1 U26979 ( .A(n45212), .B(n45211), .C(n45210), .D(n45209), .Y(n45213)
         );
  NAND4X1 U26980 ( .A(n43967), .B(n43966), .C(n43965), .D(n43964), .Y(n48334)
         );
  XOR2X1 U26981 ( .A(n41847), .B(n36900), .Y(n27399) );
  OR4X1 U26982 ( .A(n27448), .B(n27449), .C(n27450), .D(n27451), .Y(n41670) );
  NOR2X1 U26983 ( .A(n44909), .B(n44908), .Y(n46473) );
  NAND4X1 U26984 ( .A(n44903), .B(n44902), .C(n44901), .D(n44900), .Y(n44909)
         );
  NAND4X1 U26985 ( .A(n44907), .B(n44906), .C(n44905), .D(n44904), .Y(n44908)
         );
  NOR2X1 U26986 ( .A(n36996), .B(n37317), .Y(n39949) );
  NOR2X1 U26987 ( .A(n12799), .B(n45895), .Y(n45899) );
  NAND4X2 U26988 ( .A(n45366), .B(n45365), .C(n45364), .D(n45363), .Y(
        net209602) );
  NOR4X1 U26989 ( .A(n45362), .B(n45361), .C(n45360), .D(n45359), .Y(n45363)
         );
  NOR4X1 U26990 ( .A(n45358), .B(n45357), .C(n45356), .D(n45355), .Y(n45364)
         );
  NOR4X1 U26991 ( .A(n45350), .B(n45349), .C(n45348), .D(n45347), .Y(n45366)
         );
  NOR4X1 U26992 ( .A(n45292), .B(n45291), .C(n45290), .D(n45289), .Y(n45308)
         );
  NOR4X1 U26993 ( .A(n45300), .B(n45299), .C(n45298), .D(n45297), .Y(n45306)
         );
  NOR4X1 U26994 ( .A(n45304), .B(n45303), .C(n45302), .D(n45301), .Y(n45305)
         );
  NAND4X1 U26995 ( .A(n45397), .B(n45396), .C(n45395), .D(n45394), .Y(
        net210669) );
  NOR4X1 U26996 ( .A(n45389), .B(n45388), .C(n45387), .D(n45386), .Y(n45395)
         );
  NOR4X1 U26997 ( .A(n45381), .B(n45380), .C(n45379), .D(n45378), .Y(n45397)
         );
  NOR4X1 U26998 ( .A(n45393), .B(n45392), .C(n45391), .D(n45390), .Y(n45394)
         );
  NAND4X1 U26999 ( .A(n44783), .B(n44782), .C(n44781), .D(n44780), .Y(
        net213687) );
  NOR4X1 U27000 ( .A(n44779), .B(n44778), .C(n44777), .D(n44776), .Y(n44780)
         );
  NOR4X1 U27001 ( .A(n44775), .B(n44774), .C(n44773), .D(n44772), .Y(n44781)
         );
  NAND3X1 U27002 ( .A(net214433), .B(net214435), .C(n37196), .Y(net209583) );
  NOR4X1 U27003 ( .A(n44833), .B(n44832), .C(n44831), .D(n44830), .Y(net214433) );
  NOR4BBX1 U27004 ( .AN(n41728), .BN(n41729), .C(n44839), .D(n44838), .Y(
        net214435) );
  NAND2X1 U27005 ( .A(n41644), .B(n41645), .Y(n45038) );
  NOR4X1 U27006 ( .A(n45036), .B(n45035), .C(n45034), .D(n45033), .Y(n45042)
         );
  XOR2X1 U27007 ( .A(n9667), .B(n41283), .Y(n45270) );
  NOR4X1 U27008 ( .A(n45268), .B(n45267), .C(n45266), .D(n45265), .Y(n45274)
         );
  XOR2X1 U27009 ( .A(n41807), .B(n42607), .Y(n45064) );
  XOR2X1 U27010 ( .A(n41803), .B(n40039), .Y(n45073) );
  NAND2X1 U27011 ( .A(n41712), .B(n41713), .Y(n41711) );
  XNOR2X1 U27012 ( .A(n42062), .B(n42706), .Y(n41712) );
  NOR2X1 U27013 ( .A(n45068), .B(n41734), .Y(n45079) );
  NAND2X1 U27014 ( .A(n41346), .B(n41347), .Y(n45008) );
  NOR4X1 U27015 ( .A(n45014), .B(n45013), .C(n45012), .D(n45011), .Y(n45020)
         );
  XOR2X1 U27016 ( .A(n42064), .B(n42659), .Y(n45013) );
  NOR4X1 U27017 ( .A(n44883), .B(n44882), .C(n44881), .D(n44880), .Y(n44899)
         );
  NOR2X1 U27018 ( .A(n41157), .B(n40937), .Y(n40810) );
  NOR2X1 U27019 ( .A(net260332), .B(n40938), .Y(n40937) );
  NAND2X1 U27020 ( .A(n41158), .B(n41156), .Y(n41157) );
  NAND2X1 U27021 ( .A(n_cell_303546_net275998), .B(n10976), .Y(n40938) );
  NAND2X1 U27022 ( .A(n10969), .B(n10968), .Y(n40811) );
  NOR2X1 U27023 ( .A(n41101), .B(n40939), .Y(n41100) );
  AOI21X2 U27024 ( .A0(n40835), .A1(n40836), .B0(n40837), .Y(n40834) );
  NAND2X1 U27025 ( .A(n11263), .B(n11262), .Y(n40841) );
  NOR2X1 U27026 ( .A(n39343), .B(n_cell_301249_net269731), .Y(n40839) );
  CLKINVX1 U27027 ( .A(n11264), .Y(n_cell_301249_net269731) );
  CLKINVX1 U27028 ( .A(net271515), .Y(net151562) );
  NAND3BX1 U27029 ( .AN(n41034), .B(n41035), .C(n41036), .Y(n40865) );
  NAND2X1 U27030 ( .A(n10302), .B(n11869), .Y(n41034) );
  NAND3X1 U27031 ( .A(n40418), .B(n40422), .C(n_cell_301249_net269943), .Y(
        n41036) );
  NAND3X1 U27032 ( .A(n40418), .B(n40422), .C(n_cell_301249_net269941), .Y(
        n41035) );
  NOR2X1 U27033 ( .A(net171315), .B(n_cell_301249_net269635), .Y(n41038) );
  NAND3X1 U27034 ( .A(n_cell_303546_net276365), .B(n11578), .C(n11870), .Y(
        n41039) );
  CLKINVX1 U27035 ( .A(n10433), .Y(n_cell_301249_net269638) );
  CLKINVX1 U27036 ( .A(net259665), .Y(net171183) );
  NAND3X1 U27037 ( .A(n_cell_303546_net276365), .B(n11578), .C(net171182), .Y(
        n41043) );
  CLKINVX1 U27038 ( .A(net259661), .Y(net171182) );
  NOR2X1 U27039 ( .A(net171180), .B(n_cell_301249_net269590), .Y(n41003) );
  NAND2X1 U27040 ( .A(n10470), .B(n12168), .Y(n41001) );
  NOR2X1 U27041 ( .A(n_cell_303546_net277852), .B(n_cell_301249_net269593),
        .Y(n41004) );
  CLKINVX1 U27042 ( .A(n11916), .Y(n_cell_301249_net269593) );
  NAND4X1 U27043 ( .A(n47335), .B(n47334), .C(n47333), .D(n47332), .Y(n47995)
         );
  NOR4X1 U27044 ( .A(n47331), .B(n47330), .C(n47329), .D(n47328), .Y(n47332)
         );
  NAND4X1 U27045 ( .A(n47324), .B(n47323), .C(n47322), .D(n47321), .Y(n47989)
         );
  NOR2X1 U27046 ( .A(n47316), .B(n47315), .Y(n47322) );
  NAND3X1 U27047 ( .A(n47313), .B(n47312), .C(net210583), .Y(n47979) );
  NAND4X1 U27048 ( .A(n47303), .B(n47302), .C(n47301), .D(n47300), .Y(n47990)
         );
  NAND4X1 U27049 ( .A(n47357), .B(n47356), .C(n47355), .D(n47354), .Y(n48000)
         );
  NOR4X1 U27050 ( .A(n47353), .B(n47352), .C(n47351), .D(n47350), .Y(n47354)
         );
  NAND4X1 U27051 ( .A(n47346), .B(n47345), .C(n47344), .D(n47343), .Y(n47996)
         );
  NAND4X1 U27052 ( .A(n47379), .B(n47378), .C(n47377), .D(n47376), .Y(n47997)
         );
  NAND4X1 U27053 ( .A(n47368), .B(n47367), .C(n47366), .D(n47365), .Y(n47974)
         );
  NOR4X1 U27054 ( .A(n47364), .B(n47363), .C(n47362), .D(n47361), .Y(n47365)
         );
  NAND4X1 U27055 ( .A(n47412), .B(n47411), .C(n47410), .D(n47409), .Y(n48011)
         );
  NAND4X1 U27056 ( .A(n47423), .B(n47422), .C(n47421), .D(n47420), .Y(n48019)
         );
  NOR4X1 U27057 ( .A(n47419), .B(n47418), .C(n47417), .D(n47416), .Y(n47420)
         );
  NAND4X1 U27058 ( .A(n47390), .B(n47389), .C(n47388), .D(n47387), .Y(n48007)
         );
  NAND4X1 U27059 ( .A(n47401), .B(n47400), .C(n47399), .D(n47398), .Y(n48005)
         );
  NAND4X1 U27060 ( .A(n47445), .B(n47444), .C(n47443), .D(n47442), .Y(n47975)
         );
  NAND4X1 U27061 ( .A(n47434), .B(n47433), .C(n47432), .D(n47431), .Y(n47998)
         );
  NAND4X1 U27062 ( .A(n47467), .B(n47466), .C(n47465), .D(n47464), .Y(n48009)
         );
  NOR4X1 U27063 ( .A(n47463), .B(n47462), .C(n47461), .D(n47460), .Y(n47464)
         );
  NAND4X1 U27064 ( .A(n47456), .B(n47455), .C(n47454), .D(n47453), .Y(n48006)
         );
  AOI21X1 U27065 ( .A0(n40471), .A1(n40472), .B0(n40473), .Y(n40470) );
  NOR3BXL U27066 ( .AN(n40731), .B(n_cell_301249_net269583), .C(
        n_cell_301249_net269578), .Y(n40471) );
  NAND3BX1 U27067 ( .AN(n_cell_303546_net277843), .B(n40732), .C(net271999),
        .Y(n40473) );
  NAND2X1 U27068 ( .A(n40761), .B(n40730), .Y(n40472) );
  NAND3X1 U27069 ( .A(n11925), .B(n10471), .C(n40733), .Y(n40475) );
  NAND2X1 U27070 ( .A(n39551), .B(n11924), .Y(n40733) );
  NAND2X1 U27071 ( .A(n_cell_303546_net277936), .B(n10471), .Y(n40735) );
  NAND2X1 U27072 ( .A(n12806), .B(n11917), .Y(n40736) );
  CLKINVX1 U27073 ( .A(net271996), .Y(net171180) );
  CLKINVX1 U27074 ( .A(n12614), .Y(n_cell_303546_net277412) );
  CLKINVX1 U27075 ( .A(n10436), .Y(n_cell_303546_net277698) );
  NOR2BX1 U27076 ( .AN(n40628), .B(n40627), .Y(n40504) );
  NAND2X1 U27077 ( .A(n11568), .B(net214783), .Y(n40627) );
  NOR2X1 U27078 ( .A(n40501), .B(n40581), .Y(n40628) );
  NOR2BX1 U27079 ( .AN(net260352), .B(net260355), .Y(n40501) );
  OAI211X1 U27080 ( .A0(net171280), .A1(net214782), .B0(n11567), .C0(n11566),
        .Y(n40505) );
  CLKINVX1 U27081 ( .A(n11566), .Y(n_cell_303546_net277696) );
  AOI21X1 U27082 ( .A0(n39622), .A1(n11274), .B0(n40699), .Y(n40698) );
  NAND3X1 U27083 ( .A(n10646), .B(n12848), .C(net260474), .Y(n40699) );
  NAND2X1 U27084 ( .A(n11265), .B(n13025), .Y(n40701) );
  AOI21X1 U27085 ( .A0(n40700), .A1(net260474), .B0(n40524), .Y(n40702) );
  NOR2X1 U27086 ( .A(net260470), .B(n_cell_303546_net277536), .Y(n40524) );
  NOR2X1 U27087 ( .A(n_cell_303546_net277536), .B(n11272), .Y(n40700) );
  NOR2X1 U27088 ( .A(n_cell_303546_net277795), .B(net171530), .Y(n40703) );
  CLKINVX1 U27089 ( .A(n11524), .Y(n_cell_303546_net277795) );
  NOR2X1 U27090 ( .A(n37096), .B(n37448), .Y(n40596) );
  NOR2X1 U27091 ( .A(n40544), .B(n40549), .Y(n40548) );
  NAND2X1 U27092 ( .A(net209124), .B(n40651), .Y(n40549) );
  AOI21X1 U27093 ( .A0(n40545), .A1(n40546), .B0(n40547), .Y(n40544) );
  NOR2X1 U27094 ( .A(n40573), .B(n40652), .Y(n40651) );
  OAI21XL U27095 ( .A0(net171408), .A1(net212037), .B0(n40653), .Y(n40654) );
  NOR2X1 U27096 ( .A(net171416), .B(net151571), .Y(n40653) );
  AOI21X1 U27097 ( .A0(net151566), .A1(n10959), .B0(n40656), .Y(n40657) );
  NAND2X1 U27098 ( .A(n10960), .B(n10957), .Y(n40656) );
  NAND2X1 U27099 ( .A(net212088), .B(n10206), .Y(n40658) );
  CLKINVX1 U27100 ( .A(n10958), .Y(n_cell_303546_net277735) );
  NOR2X1 U27101 ( .A(n_cell_303546_net277738), .B(net151586), .Y(n40659) );
  NAND2X1 U27102 ( .A(n10485), .B(n40389), .Y(n39827) );
  OAI21XL U27103 ( .A0(n39593), .A1(n39597), .B0(n39825), .Y(n39600) );
  AND2X2 U27104 ( .A(net261020), .B(n39826), .Y(n39825) );
  AOI21X1 U27105 ( .A0(n39594), .A1(net151430), .B0(n39595), .Y(n39593) );
  NOR2X1 U27106 ( .A(n39824), .B(net171108), .Y(n39826) );
  NAND4BX1 U27107 ( .AN(net209739), .B(net260251), .C(net259747), .D(net260427), .Y(n39602) );
  CLKINVX1 U27108 ( .A(n10492), .Y(n39601) );
  NOR2X1 U27109 ( .A(n39753), .B(n39757), .Y(n39756) );
  NAND2BX1 U27110 ( .AN(n40404), .B(n_cell_301249_net269615), .Y(n39757) );
  AOI21X1 U27111 ( .A0(n39754), .A1(n39755), .B0(n39750), .Y(n39753) );
  CLKINVX1 U27112 ( .A(n10083), .Y(n39755) );
  NAND2X1 U27113 ( .A(n11613), .B(n11614), .Y(n39857) );
  AND2X2 U27114 ( .A(net259645), .B(net259641), .Y(n39856) );
  NOR2X1 U27115 ( .A(net171474), .B(n39987), .Y(n39986) );
  OAI21XL U27116 ( .A0(n39526), .A1(n10227), .B0(n40014), .Y(n40018) );
  CLKINVX1 U27117 ( .A(n10228), .Y(n40014) );
  NOR2X1 U27118 ( .A(n39522), .B(n39525), .Y(n39526) );
  AOI21X1 U27119 ( .A0(n39523), .A1(n39524), .B0(n10814), .Y(n39522) );
  CLKINVX1 U27120 ( .A(n10223), .Y(n40013) );
  NOR2X1 U27121 ( .A(n37042), .B(n37444), .Y(n40588) );
  NOR2X1 U27122 ( .A(n39919), .B(n_cell_301249_net269701), .Y(n39918) );
  OAI21XL U27123 ( .A0(n10661), .A1(n39673), .B0(n39914), .Y(n40032) );
  NOR3BXL U27124 ( .AN(n39915), .B(n39916), .C(net210034), .Y(n39914) );
  AOI21X1 U27125 ( .A0(n36926), .A1(n39674), .B0(n39675), .Y(n39673) );
  NOR2X1 U27126 ( .A(net151514), .B(n39917), .Y(n39915) );
  CLKINVX1 U27127 ( .A(n10758), .Y(n40033) );
  NOR2X1 U27128 ( .A(n11742), .B(n46172), .Y(n46176) );
  NOR2X1 U27129 ( .A(n12153), .B(n45818), .Y(n45822) );
  NOR2X1 U27130 ( .A(n45803), .B(n40386), .Y(n45807) );
  NAND4X1 U27131 ( .A(n44246), .B(n44245), .C(n44244), .D(n44243), .Y(n11732)
         );
  NAND2X1 U27132 ( .A(n41247), .B(n41218), .Y(n41249) );
  NAND4X1 U27133 ( .A(n44602), .B(n44601), .C(n44600), .D(n44599), .Y(n11743)
         );
  NOR4X1 U27134 ( .A(n26725), .B(n26726), .C(n26727), .D(n26728), .Y(n44606)
         );
  OR2X1 U27135 ( .A(n47948), .B(n47947), .Y(net207653) );
  NAND4X1 U27136 ( .A(n47531), .B(n47530), .C(n47529), .D(n47528), .Y(n48029)
         );
  NAND4X1 U27137 ( .A(n47520), .B(n47519), .C(n47518), .D(n47517), .Y(n48034)
         );
  NAND4X1 U27138 ( .A(n47542), .B(n47541), .C(n47540), .D(n47539), .Y(n48032)
         );
  NAND4X1 U27139 ( .A(n47551), .B(n47550), .C(n47549), .D(n47548), .Y(n48027)
         );
  NAND4X1 U27140 ( .A(n47290), .B(n47289), .C(n47288), .D(n47287), .Y(
        net210234) );
  NAND4X1 U27141 ( .A(n47285), .B(n47284), .C(n47283), .D(n47282), .Y(
        net210148) );
  NAND4X1 U27142 ( .A(n47577), .B(n47576), .C(n47575), .D(n47574), .Y(n48036)
         );
  NAND4X1 U27143 ( .A(n47566), .B(n47565), .C(n47564), .D(n47563), .Y(n48038)
         );
  NAND4X1 U27144 ( .A(n47556), .B(n47555), .C(n47554), .D(n47553), .Y(n48040)
         );
  NAND4X1 U27145 ( .A(n47500), .B(n47499), .C(n47498), .D(n47497), .Y(n48028)
         );
  NAND3BX1 U27146 ( .AN(n41719), .B(n47509), .C(net209288), .Y(n48030) );
  OR4X1 U27147 ( .A(n47504), .B(n47503), .C(n47502), .D(n47501), .Y(n41719) );
  NAND4X1 U27148 ( .A(n47489), .B(n47488), .C(n47487), .D(n47486), .Y(n48018)
         );
  NAND4X1 U27149 ( .A(n47478), .B(n47477), .C(n47476), .D(n47475), .Y(n48020)
         );
  NAND4X1 U27150 ( .A(n47035), .B(n47034), .C(n47033), .D(n47032), .Y(
        net210132) );
  NAND4X1 U27151 ( .A(n47896), .B(n47895), .C(n47894), .D(n47893), .Y(n12970)
         );
  XOR2X1 U27152 ( .A(n36757), .B(n41806), .Y(n47664) );
  NAND2X1 U27153 ( .A(n47688), .B(n47687), .Y(n47693) );
  NAND4X1 U27154 ( .A(n47622), .B(n47621), .C(n47620), .D(n47619), .Y(
        net210615) );
  NOR4X1 U27155 ( .A(n47618), .B(n47617), .C(n47616), .D(n47615), .Y(n47619)
         );
  NAND4X1 U27156 ( .A(n47611), .B(n47610), .C(n47609), .D(n47608), .Y(
        net210213) );
  NOR4X1 U27157 ( .A(n47585), .B(n47584), .C(n47583), .D(n47582), .Y(n47586)
         );
  NAND4X1 U27158 ( .A(n47600), .B(n47599), .C(n47598), .D(n47597), .Y(
        net210207) );
  NOR4X1 U27159 ( .A(n47596), .B(n47595), .C(n47594), .D(n47593), .Y(n47597)
         );
  NOR2X1 U27160 ( .A(n12297), .B(n47853), .Y(n47857) );
  NOR4X1 U27161 ( .A(n29320), .B(n29321), .C(n29322), .D(n29323), .Y(n43636)
         );
  NOR4X1 U27162 ( .A(n45495), .B(n45494), .C(n45493), .D(n45492), .Y(n45511)
         );
  NOR4X1 U27163 ( .A(n45503), .B(n45502), .C(n45501), .D(n45500), .Y(n45509)
         );
  NOR4X1 U27164 ( .A(n45507), .B(n45506), .C(n45505), .D(n45504), .Y(n45508)
         );
  NOR4X1 U27165 ( .A(n45477), .B(n45476), .C(n45475), .D(n45474), .Y(n45483)
         );
  AND2X2 U27166 ( .A(net213733), .B(net213732), .Y(n39777) );
  NOR2X1 U27167 ( .A(n11688), .B(n43755), .Y(n43759) );
  NAND4X1 U27168 ( .A(n45842), .B(n45841), .C(n45840), .D(n45839), .Y(n48522)
         );
  NOR2X1 U27169 ( .A(n23178), .B(n23177), .Y(n45840) );
  NAND4X1 U27170 ( .A(n47926), .B(n47925), .C(n47924), .D(n47923), .Y(n12909)
         );
  NOR2X1 U27171 ( .A(n12264), .B(n46680), .Y(n46684) );
  NOR2X1 U27172 ( .A(n12316), .B(n47204), .Y(n47208) );
  NAND4X1 U27173 ( .A(n47163), .B(n47162), .C(n47161), .D(n47160), .Y(
        net210109) );
  NAND4X1 U27174 ( .A(n47881), .B(n47880), .C(n47879), .D(n47878), .Y(n12942)
         );
  NOR2X1 U27175 ( .A(n19791), .B(n19790), .Y(n47879) );
  NAND4X1 U27176 ( .A(n47886), .B(n47885), .C(n47884), .D(n47883), .Y(n12940)
         );
  NAND4X1 U27177 ( .A(n47062), .B(n47061), .C(n47060), .D(n47059), .Y(n12918)
         );
  NOR2X1 U27178 ( .A(n19982), .B(n19981), .Y(n47060) );
  NOR2X1 U27179 ( .A(n37383), .B(n37116), .Y(n39909) );
  NAND3X1 U27180 ( .A(net212171), .B(net212170), .C(net212172), .Y(
        n_cell_301249_net267269) );
  NAND3X1 U27181 ( .A(net212176), .B(net212175), .C(net212177), .Y(
        n_cell_301249_net267275) );
  NOR2BX1 U27182 ( .AN(net209622), .B(n46573), .Y(net256309) );
  XOR2X1 U27183 ( .A(n41815), .B(n42519), .Y(n45217) );
  XOR2X1 U27184 ( .A(n41816), .B(n42518), .Y(n45186) );
  NAND2X1 U27185 ( .A(net212262), .B(n36934), .Y(n48143) );
  NOR2X2 U27186 ( .A(n45107), .B(n45106), .Y(n46482) );
  NAND4X1 U27187 ( .A(n45101), .B(n45100), .C(n45099), .D(n45098), .Y(n45107)
         );
  NAND4X1 U27188 ( .A(n45105), .B(n45104), .C(n45103), .D(n45102), .Y(n45106)
         );
  NOR4X1 U27189 ( .A(n44860), .B(n44859), .C(n44858), .D(n44857), .Y(n44871)
         );
  NAND2X1 U27190 ( .A(n48175), .B(n48172), .Y(net210682) );
  NOR2X1 U27191 ( .A(n10394), .B(n44164), .Y(n44168) );
  NOR2X1 U27192 ( .A(n12582), .B(n44173), .Y(n44177) );
  OR4X1 U27193 ( .A(n27478), .B(n27479), .C(n27480), .D(n27481), .Y(n41672) );
  NAND4X1 U27194 ( .A(n43854), .B(n43853), .C(n43852), .D(n43851), .Y(n48132)
         );
  NOR2X1 U27195 ( .A(n43850), .B(n45530), .Y(n43854) );
  NAND4X1 U27196 ( .A(n43916), .B(n43915), .C(n43914), .D(n43913), .Y(n48130)
         );
  NOR4X1 U27197 ( .A(n43912), .B(n43911), .C(n43910), .D(n43909), .Y(n43913)
         );
  NOR4X1 U27198 ( .A(n43881), .B(n43880), .C(n43879), .D(n43878), .Y(n43882)
         );
  NOR2X1 U27199 ( .A(n43875), .B(n48335), .Y(n43885) );
  NOR4X1 U27200 ( .A(n26669), .B(n26670), .C(n26671), .D(n26672), .Y(n44305)
         );
  NOR4X1 U27201 ( .A(n26677), .B(n26678), .C(n26679), .D(n26680), .Y(n44303)
         );
  NOR4X1 U27202 ( .A(n26665), .B(n26666), .C(n26667), .D(n26668), .Y(n44306)
         );
  NAND4X1 U27203 ( .A(n44507), .B(n44506), .C(n44505), .D(n44504), .Y(n12702)
         );
  NOR2X1 U27204 ( .A(n24947), .B(n24946), .Y(n44505) );
  NOR4X1 U27205 ( .A(n24945), .B(n24944), .C(n24943), .D(n24942), .Y(n44504)
         );
  NAND4X1 U27206 ( .A(n44516), .B(n44515), .C(n44514), .D(n44513), .Y(n12706)
         );
  NAND2X1 U27207 ( .A(n37299), .B(net171305), .Y(n10544) );
  NAND4X1 U27208 ( .A(n44484), .B(n44483), .C(n44482), .D(n44481), .Y(n12049)
         );
  CLKBUFX3 U27209 ( .A(n12048), .Y(n40392) );
  NAND2BX1 U27210 ( .AN(n44570), .B(n44466), .Y(n12151) );
  NOR2X1 U27211 ( .A(n25094), .B(n25097), .Y(n44464) );
  NAND4BBX1 U27212 ( .AN(n47948), .BN(n47947), .C(n44451), .D(n44450), .Y(
        n12152) );
  NAND4X1 U27213 ( .A(n44431), .B(n44430), .C(n44429), .D(n44428), .Y(n12711)
         );
  NOR2X1 U27214 ( .A(n37053), .B(n37465), .Y(n40962) );
  NOR4X1 U27215 ( .A(n44925), .B(n44924), .C(n44923), .D(n44922), .Y(n44926)
         );
  NOR4X1 U27216 ( .A(n44976), .B(n44975), .C(n44974), .D(n44973), .Y(n44982)
         );
  OR4X1 U27217 ( .A(n44968), .B(n44967), .C(n44966), .D(n44965), .Y(n41697) );
  NOR4X1 U27218 ( .A(n45148), .B(n45147), .C(n45146), .D(n45145), .Y(n45154)
         );
  NOR4X1 U27219 ( .A(n45140), .B(n45139), .C(n45138), .D(n45137), .Y(n45156)
         );
  NOR4X1 U27220 ( .A(n45152), .B(n45151), .C(n45150), .D(n45149), .Y(n45153)
         );
  NAND2X1 U27221 ( .A(n41657), .B(n41658), .Y(n44948) );
  OR4X1 U27222 ( .A(n44961), .B(n44960), .C(n44959), .D(n44958), .Y(n41705) );
  NOR4BBX1 U27223 ( .AN(n41730), .BN(n41731), .C(n45121), .D(n45120), .Y(
        n45122) );
  NOR4X1 U27224 ( .A(n45119), .B(n45118), .C(n45117), .D(n45116), .Y(n45123)
         );
  NOR4X1 U27225 ( .A(n45208), .B(n45207), .C(n45206), .D(n45205), .Y(n45214)
         );
  NOR4X1 U27226 ( .A(n45200), .B(n45199), .C(n45198), .D(n45197), .Y(n45216)
         );
  XOR2X1 U27227 ( .A(n41816), .B(n42595), .Y(n45418) );
  NOR4X1 U27228 ( .A(n45175), .B(n45174), .C(n45173), .D(n45172), .Y(n45184)
         );
  NAND2X1 U27229 ( .A(n48336), .B(n48288), .Y(net210635) );
  NOR4X1 U27230 ( .A(n31543), .B(n31544), .C(n31545), .D(n31546), .Y(n43221)
         );
  NOR4X1 U27231 ( .A(n31303), .B(n31304), .C(n31305), .D(n31306), .Y(n43292)
         );
  NOR2X1 U27232 ( .A(n37001), .B(n37226), .Y(n39419) );
  NOR2X1 U27233 ( .A(n37211), .B(n39779), .Y(n39418) );
  NOR2X1 U27234 ( .A(n46376), .B(n48138), .Y(net212474) );
  NAND2X1 U27235 ( .A(net212476), .B(net212475), .Y(n39779) );
  NOR2X1 U27236 ( .A(n46332), .B(net209898), .Y(n46342) );
  NAND4X2 U27237 ( .A(n46353), .B(n46352), .C(n46351), .D(n46350), .Y(
        net209316) );
  NOR4X1 U27238 ( .A(n46327), .B(n46326), .C(n46325), .D(n46324), .Y(n46328)
         );
  NAND3X1 U27239 ( .A(net212387), .B(net212386), .C(net212388), .Y(n39416) );
  NAND2BX1 U27240 ( .AN(n39417), .B(net212374), .Y(net209313) );
  NAND2X1 U27241 ( .A(n39778), .B(net212377), .Y(n39417) );
  NOR2X1 U27242 ( .A(n46463), .B(net209930), .Y(net212374) );
  NOR2X1 U27243 ( .A(n37000), .B(n37229), .Y(n39778) );
  NAND4X1 U27244 ( .A(n46400), .B(n46399), .C(n46398), .D(n46397), .Y(
        net209298) );
  NAND4X2 U27245 ( .A(n46422), .B(n46421), .C(n46420), .D(n46419), .Y(
        net209296) );
  AND2X2 U27246 ( .A(n48449), .B(n48446), .Y(net234488) );
  NAND4X2 U27247 ( .A(n46554), .B(n46553), .C(n46552), .D(n46551), .Y(
        net209320) );
  NAND4X1 U27248 ( .A(n46543), .B(n46542), .C(n46541), .D(n46540), .Y(
        net209323) );
  NOR4X1 U27249 ( .A(n46539), .B(n46538), .C(n46537), .D(n46536), .Y(n46540)
         );
  NAND2X1 U27250 ( .A(n47705), .B(n48436), .Y(net210581) );
  NAND3BX2 U27251 ( .AN(n41724), .B(n46596), .C(n48142), .Y(net210580) );
  OR4X1 U27252 ( .A(n46590), .B(n46589), .C(n46588), .D(n46587), .Y(n41724) );
  NAND4X1 U27253 ( .A(n47011), .B(n47010), .C(n47009), .D(n47008), .Y(n12342)
         );
  NAND4X1 U27254 ( .A(n44070), .B(n44069), .C(n44068), .D(n44067), .Y(n48166)
         );
  NOR4X1 U27255 ( .A(n44066), .B(n44065), .C(n44064), .D(n44063), .Y(n44067)
         );
  NAND2BX1 U27256 ( .AN(n39414), .B(net212642), .Y(net209291) );
  NAND2X1 U27257 ( .A(n39780), .B(net212643), .Y(n39414) );
  NOR2X1 U27258 ( .A(n46232), .B(n48171), .Y(net212642) );
  NAND4X1 U27259 ( .A(n46259), .B(n46258), .C(n46257), .D(n46256), .Y(
        net210919) );
  NOR4X1 U27260 ( .A(n46255), .B(n46254), .C(n46253), .D(n46252), .Y(n46256)
         );
  NAND4X1 U27261 ( .A(n46270), .B(n46269), .C(n46268), .D(n46267), .Y(
        net209303) );
  NAND4X1 U27262 ( .A(n46292), .B(n46291), .C(n46290), .D(n46289), .Y(n48464)
         );
  NAND4X1 U27263 ( .A(n46281), .B(n46280), .C(n46279), .D(n46278), .Y(n48461)
         );
  NOR2X1 U27264 ( .A(n46273), .B(n46272), .Y(n46279) );
  NOR4X1 U27265 ( .A(n46277), .B(n46276), .C(n46275), .D(n46274), .Y(n46278)
         );
  NOR2X1 U27266 ( .A(n46179), .B(n48187), .Y(n46183) );
  NAND2X1 U27267 ( .A(n48465), .B(n48427), .Y(net210584) );
  NAND2X1 U27268 ( .A(n48467), .B(n48426), .Y(net210559) );
  NOR2X1 U27269 ( .A(n43736), .B(n48383), .Y(n43740) );
  NOR2X1 U27270 ( .A(n12007), .B(n45930), .Y(n45934) );
  NOR2X1 U27271 ( .A(n37022), .B(n37451), .Y(n_cell_301249_net267308) );
  NAND3X4 U27272 ( .A(net213901), .B(net213902), .C(n39461), .Y(net209603) );
  NOR4X1 U27273 ( .A(n45331), .B(n45330), .C(n45329), .D(n45328), .Y(net213901) );
  NOR4X1 U27274 ( .A(n45335), .B(n45334), .C(n45333), .D(n45332), .Y(net213902) );
  NOR2X2 U27275 ( .A(n36940), .B(n37198), .Y(n39461) );
  CLKINVX1 U27276 ( .A(net213687), .Y(net209582) );
  CLKINVX1 U27277 ( .A(net209583), .Y(net209592) );
  NAND4X2 U27278 ( .A(n44692), .B(n44691), .C(n44690), .D(n44689), .Y(
        net210670) );
  NOR4X1 U27279 ( .A(n44676), .B(n44675), .C(n44674), .D(n44673), .Y(n44692)
         );
  NOR4X1 U27280 ( .A(n44810), .B(n44809), .C(n44808), .D(n44807), .Y(n44811)
         );
  NOR4X1 U27281 ( .A(n44798), .B(n44797), .C(n44796), .D(n44795), .Y(n44814)
         );
  CLKINVX1 U27282 ( .A(n39712), .Y(net235251) );
  NAND2BX1 U27283 ( .AN(net210641), .B(n39713), .Y(n39712) );
  CLKINVX1 U27284 ( .A(net210646), .Y(n39713) );
  NOR4X1 U27285 ( .A(n45040), .B(n45039), .C(n45038), .D(n45037), .Y(n45041)
         );
  NOR4X1 U27286 ( .A(n45028), .B(n45027), .C(n45026), .D(n45025), .Y(n45044)
         );
  NAND4X1 U27287 ( .A(n45276), .B(n45275), .C(n45274), .D(n45273), .Y(
        net213680) );
  NOR4X1 U27288 ( .A(n45264), .B(n45263), .C(n45262), .D(n45261), .Y(n45275)
         );
  NOR4X1 U27289 ( .A(n45260), .B(n45259), .C(n45258), .D(n45257), .Y(n45276)
         );
  NOR4X1 U27290 ( .A(n45272), .B(n45271), .C(n45270), .D(n45269), .Y(n45273)
         );
  NAND4X2 U27291 ( .A(n45022), .B(n45021), .C(n45020), .D(n45019), .Y(
        net213679) );
  NOR4X1 U27292 ( .A(n45010), .B(n45009), .C(n45008), .D(n45007), .Y(n45021)
         );
  NOR4X1 U27293 ( .A(n45006), .B(n45005), .C(n45004), .D(n45003), .Y(n45022)
         );
  NOR4X1 U27294 ( .A(n44891), .B(n44890), .C(n44889), .D(n44888), .Y(n44897)
         );
  NOR4X1 U27295 ( .A(n44895), .B(n44894), .C(n44893), .D(n44892), .Y(n44896)
         );
  NOR4X1 U27296 ( .A(n44887), .B(n44886), .C(n44885), .D(n44884), .Y(n44898)
         );
  NAND4X1 U27297 ( .A(n45254), .B(n45253), .C(n45252), .D(n45251), .Y(
        net210665) );
  NOR4X1 U27298 ( .A(n45243), .B(n45242), .C(n45241), .D(n45240), .Y(n45253)
         );
  NOR4BX1 U27299 ( .AN(n41725), .B(n45250), .C(n45249), .D(n45248), .Y(n45251)
         );
  NAND2X1 U27300 ( .A(n41389), .B(n41390), .Y(n45086) );
  XOR2X1 U27301 ( .A(n42066), .B(n42659), .Y(n45087) );
  NOR4X1 U27302 ( .A(n45093), .B(n45092), .C(n45091), .D(n45090), .Y(net214154) );
  NAND2X1 U27303 ( .A(n41235), .B(n41236), .Y(n45090) );
  NAND2X1 U27304 ( .A(n41369), .B(n41370), .Y(n45084) );
  NAND2X1 U27305 ( .A(n41637), .B(n41638), .Y(n45083) );
  NAND2X1 U27306 ( .A(n41808), .B(n41636), .Y(n41637) );
  NAND2X1 U27307 ( .A(n37200), .B(n42609), .Y(n41638) );
  CLKINVX1 U27308 ( .A(n42597), .Y(n41636) );
  NOR2X1 U27309 ( .A(net151571), .B(net151566), .Y(n40813) );
  NAND2X1 U27310 ( .A(n10959), .B(n10960), .Y(n40815) );
  CLKINVX1 U27311 ( .A(n12213), .Y(net171403) );
  CLKINVX1 U27312 ( .A(n10635), .Y(n_cell_301249_net269740) );
  AOI31X1 U27313 ( .A0(n39342), .A1(n10761), .A2(n10641), .B0(n41105), .Y(
        n40844) );
  NAND2X1 U27314 ( .A(n10760), .B(n10759), .Y(n41105) );
  NAND2X1 U27315 ( .A(n10638), .B(n_cell_301249_net269738), .Y(n40845) );
  NOR2X1 U27316 ( .A(n41042), .B(n41041), .Y(n40868) );
  NAND2X1 U27317 ( .A(n41043), .B(n41044), .Y(n41042) );
  NAND2X1 U27318 ( .A(n11575), .B(n11576), .Y(n41041) );
  NAND3X1 U27319 ( .A(n_cell_303546_net276365), .B(n11578), .C(net171183), .Y(
        n41044) );
  NAND2X1 U27320 ( .A(net260352), .B(net260355), .Y(n40869) );
  CLKINVX1 U27321 ( .A(n11567), .Y(n_cell_301249_net269646) );
  NAND2X1 U27322 ( .A(n12807), .B(net260403), .Y(n40899) );
  NAND2X1 U27323 ( .A(net272583), .B(net260925), .Y(n41008) );
  NAND2X1 U27324 ( .A(n48011), .B(n48019), .Y(net210598) );
  NAND2X1 U27325 ( .A(n48007), .B(n48005), .Y(net210596) );
  NAND2X1 U27326 ( .A(n47998), .B(n47975), .Y(net210618) );
  NAND2X1 U27327 ( .A(n48006), .B(n48009), .Y(net210601) );
  NAND3X1 U27328 ( .A(n40739), .B(n40740), .C(n40741), .Y(n40479) );
  NAND3X1 U27329 ( .A(net260403), .B(net260299), .C(n39835), .Y(n40741) );
  NAND2BX1 U27330 ( .AN(net260295), .B(net260403), .Y(n40740) );
  NOR2X1 U27331 ( .A(n_cell_303546_net277854), .B(n39550), .Y(n40739) );
  NOR3BXL U27332 ( .AN(n10464), .B(n40738), .C(n_cell_303546_net277405), .Y(
        n40478) );
  CLKINVX1 U27333 ( .A(net260299), .Y(n_cell_303546_net277405) );
  OAI21XL U27334 ( .A0(n_cell_303546_net277852), .A1(n11916), .B0(net260403),
        .Y(n40738) );
  AOI21X1 U27335 ( .A0(n_cell_303546_net277859), .A1(n11906), .B0(
        n_cell_303546_net277412), .Y(n40742) );
  CLKINVX1 U27336 ( .A(n11907), .Y(n_cell_303546_net277859) );
  NOR2X1 U27337 ( .A(net260925), .B(n_cell_303546_net277412), .Y(n40480) );
  NAND2X1 U27338 ( .A(n12611), .B(net209697), .Y(n40744) );
  NOR2BX1 U27339 ( .AN(net272625), .B(net151380), .Y(n40630) );
  CLKINVX1 U27340 ( .A(net259677), .Y(n_cell_303546_net277490) );
  NOR2X1 U27341 ( .A(n40507), .B(n40502), .Y(n40506) );
  OAI21XL U27342 ( .A0(n_cell_303546_net277696), .A1(n11565), .B0(n40629), .Y(
        n40507) );
  AOI21X1 U27343 ( .A0(n40503), .A1(n40504), .B0(n40505), .Y(n40502) );
  NOR2X1 U27344 ( .A(n_cell_303546_net277490), .B(n_cell_303546_net277698),
        .Y(n40629) );
  NAND3X1 U27345 ( .A(n11525), .B(net271515), .C(n40704), .Y(n40530) );
  NAND2X1 U27346 ( .A(n_cell_303546_net277994), .B(n11524), .Y(n40704) );
  CLKINVX1 U27347 ( .A(n11263), .Y(n_cell_303546_net277994) );
  NAND2X1 U27348 ( .A(n10761), .B(n10760), .Y(n40707) );
  NOR2X1 U27349 ( .A(n_cell_303546_net277636), .B(n12838), .Y(n40578) );
  NAND2X1 U27350 ( .A(net171528), .B(net271515), .Y(n40706) );
  NOR2X1 U27351 ( .A(n37491), .B(n37119), .Y(n40948) );
  NOR2X1 U27352 ( .A(n37137), .B(n37442), .Y(n40684) );
  NOR2X1 U27353 ( .A(n37138), .B(n37406), .Y(n40682) );
  AOI21X1 U27354 ( .A0(n40666), .A1(net211640), .B0(n40664), .Y(n40665) );
  CLKINVX1 U27355 ( .A(n12207), .Y(n40666) );
  NAND2X1 U27356 ( .A(n10947), .B(net209111), .Y(n40664) );
  NAND2X1 U27357 ( .A(net211640), .B(n40660), .Y(n40662) );
  AOI21X1 U27358 ( .A0(net171403), .A1(n12392), .B0(n40661), .Y(n40660) );
  CLKINVX1 U27359 ( .A(n12210), .Y(n40661) );
  CLKINVX1 U27360 ( .A(n12196), .Y(n40671) );
  NOR2X1 U27361 ( .A(n39599), .B(n39604), .Y(n39603) );
  NAND2X1 U27362 ( .A(net260431), .B(n39828), .Y(n39604) );
  AOI21X1 U27363 ( .A0(n39600), .A1(n39601), .B0(n39602), .Y(n39599) );
  NOR2BX1 U27364 ( .AN(n10487), .B(n39827), .Y(n39828) );
  OR2X1 U27365 ( .A(n_cell_301249_net269449), .B(n39831), .Y(n39830) );
  NAND2X1 U27366 ( .A(n10483), .B(n10484), .Y(n39831) );
  CLKINVX1 U27367 ( .A(n10610), .Y(n40026) );
  CLKINVX1 U27368 ( .A(n10480), .Y(n_cell_303546_net277630) );
  NAND2X1 U27369 ( .A(n39470), .B(n39859), .Y(n39860) );
  AND2X2 U27370 ( .A(net259649), .B(net259653), .Y(n39859) );
  NOR2BX1 U27371 ( .AN(n11607), .B(n39862), .Y(n39861) );
  NAND2X1 U27372 ( .A(net260527), .B(n10319), .Y(n39862) );
  OAI21XL U27373 ( .A0(n39855), .A1(n39758), .B0(n39858), .Y(n39472) );
  NAND3X1 U27374 ( .A(n10425), .B(n11620), .C(n39856), .Y(n39855) );
  NOR3BXL U27375 ( .AN(net260367), .B(n39857), .C(n_cell_303546_net277667),
        .Y(n39858) );
  NOR2X1 U27376 ( .A(n39756), .B(n10331), .Y(n39758) );
  AOI21X1 U27377 ( .A0(n39528), .A1(n39529), .B0(n10902), .Y(n39527) );
  NOR2X1 U27378 ( .A(net209155), .B(n39985), .Y(n39529) );
  NAND2X1 U27379 ( .A(n40018), .B(n40013), .Y(n39528) );
  NAND2X1 U27380 ( .A(n39986), .B(n10810), .Y(n39985) );
  NAND4X1 U27381 ( .A(n10806), .B(n40391), .C(n10808), .D(n10807), .Y(n39531)
         );
  CLKINVX1 U27382 ( .A(n10798), .Y(n39989) );
  NOR2X1 U27383 ( .A(n11521), .B(net171525), .Y(n39921) );
  AOI21X1 U27384 ( .A0(n39679), .A1(n39680), .B0(n10651), .Y(n39678) );
  NOR2X1 U27385 ( .A(n39920), .B(net151530), .Y(n39680) );
  NAND2X1 U27386 ( .A(n40032), .B(n40033), .Y(n39679) );
  NAND2X1 U27387 ( .A(n10659), .B(n39918), .Y(n39920) );
  CLKBUFX3 U27388 ( .A(n42455), .Y(n42475) );
  NAND4X1 U27389 ( .A(n45637), .B(n45636), .C(n45635), .D(n45634), .Y(n12386)
         );
  NOR2X1 U27390 ( .A(n24101), .B(n24100), .Y(n45635) );
  NAND4X1 U27391 ( .A(n45627), .B(n45626), .C(n45625), .D(n45624), .Y(n11204)
         );
  NOR2X1 U27392 ( .A(n24121), .B(n24120), .Y(n45625) );
  CLKBUFX3 U27393 ( .A(n11205), .Y(n40396) );
  NOR2X1 U27394 ( .A(n37082), .B(n37439), .Y(n39960) );
  NOR2X1 U27395 ( .A(n37079), .B(n37440), .Y(n39961) );
  NOR2X1 U27396 ( .A(n37078), .B(n37438), .Y(n39959) );
  NAND4X1 U27397 ( .A(n46117), .B(n46116), .C(n46115), .D(n46114), .Y(n12324)
         );
  NOR2X1 U27398 ( .A(n22421), .B(n22420), .Y(n46115) );
  NAND4X1 U27399 ( .A(n46092), .B(n46091), .C(n46090), .D(n46089), .Y(n11201)
         );
  NAND4X1 U27400 ( .A(n46102), .B(n46101), .C(n46100), .D(n46099), .Y(n12333)
         );
  NOR2X1 U27401 ( .A(n22441), .B(n22440), .Y(n46105) );
  NOR2X1 U27402 ( .A(n12025), .B(n45813), .Y(n45817) );
  NAND4X1 U27403 ( .A(n45863), .B(n45862), .C(n45861), .D(n45860), .Y(
        net209202) );
  NAND4X1 U27404 ( .A(n45852), .B(n45851), .C(n45850), .D(n45849), .Y(n11065)
         );
  NAND3X2 U27405 ( .A(net215209), .B(net215210), .C(n39451), .Y(n10369) );
  NOR4X1 U27406 ( .A(n26819), .B(n26820), .C(n26821), .D(n26822), .Y(net215210) );
  NOR2X1 U27407 ( .A(n36953), .B(n37260), .Y(n39451) );
  NAND3X1 U27408 ( .A(n39467), .B(n11741), .C(n11743), .Y(n10421) );
  NOR2BX1 U27409 ( .AN(n11744), .B(net209528), .Y(n39467) );
  NOR4X1 U27410 ( .A(n24784), .B(n24785), .C(n24786), .D(n24787), .Y(n44552)
         );
  NOR4X1 U27411 ( .A(n24922), .B(n24923), .C(n24924), .D(n24925), .Y(n44511)
         );
  NOR4X1 U27412 ( .A(n24802), .B(n24803), .C(n24804), .D(n24805), .Y(n44546)
         );
  CLKINVX1 U27413 ( .A(n11723), .Y(net171305) );
  NAND4X1 U27414 ( .A(n44426), .B(n44425), .C(n44424), .D(n44423), .Y(n11721)
         );
  NAND4BX1 U27415 ( .AN(n41671), .B(n44528), .C(n44527), .D(n44526), .Y(n12585) );
  OR4X1 U27416 ( .A(n24862), .B(n24863), .C(n24864), .D(n24865), .Y(n41671) );
  NAND4X1 U27417 ( .A(n44488), .B(n44487), .C(n44486), .D(n44485), .Y(n11722)
         );
  NAND4BX1 U27418 ( .AN(n41676), .B(n44434), .C(n44433), .D(n44432), .Y(
        net209503) );
  OR4X1 U27419 ( .A(n25162), .B(n25163), .C(n25164), .D(n25165), .Y(n41676) );
  NAND2X1 U27420 ( .A(n41273), .B(n42714), .Y(n41275) );
  NOR4X1 U27421 ( .A(n29109), .B(n29110), .C(n29111), .D(n29112), .Y(n43646)
         );
  CLKINVX1 U27422 ( .A(n48057), .Y(n12951) );
  NOR2X1 U27423 ( .A(n11116), .B(n47149), .Y(n47153) );
  NAND4X2 U27424 ( .A(n46193), .B(n46192), .C(n46191), .D(n46190), .Y(n11149)
         );
  NOR2X1 U27425 ( .A(n37027), .B(n37325), .Y(n39879) );
  NOR2X1 U27426 ( .A(n37080), .B(n37326), .Y(n39880) );
  NAND2BX1 U27427 ( .AN(n39365), .B(net211483), .Y(n10725) );
  NAND2X1 U27428 ( .A(n39890), .B(net211485), .Y(n39365) );
  NOR2X1 U27429 ( .A(n37065), .B(n37300), .Y(n39890) );
  NAND2BX1 U27430 ( .AN(n39364), .B(net211488), .Y(n10726) );
  NAND3X1 U27431 ( .A(net211490), .B(net211489), .C(net211491), .Y(n39364) );
  CLKINVX1 U27432 ( .A(net210132), .Y(net171547) );
  CLKINVX1 U27433 ( .A(n12970), .Y(net151720) );
  CLKINVX1 U27434 ( .A(net210142), .Y(net171546) );
  NAND4X1 U27435 ( .A(n46996), .B(n46995), .C(n46994), .D(n46993), .Y(n12976)
         );
  NAND4X1 U27436 ( .A(n47021), .B(n47020), .C(n47019), .D(n47018), .Y(n11442)
         );
  NAND4X1 U27437 ( .A(n47006), .B(n47005), .C(n47004), .D(n47003), .Y(n13014)
         );
  NAND3X1 U27438 ( .A(n47684), .B(n47683), .C(n47682), .Y(n47980) );
  NOR4X1 U27439 ( .A(n47681), .B(n47680), .C(n47679), .D(n47678), .Y(n47683)
         );
  CLKINVX1 U27440 ( .A(n48436), .Y(n47682) );
  NOR4X1 U27441 ( .A(n47700), .B(n47699), .C(n47698), .D(n47697), .Y(n47707)
         );
  XNOR2X1 U27442 ( .A(n36753), .B(n41809), .Y(n47696) );
  NOR2X1 U27443 ( .A(n47693), .B(n47692), .Y(n47694) );
  NOR2X1 U27444 ( .A(n47686), .B(n47685), .Y(n47695) );
  NAND4X1 U27445 ( .A(n47656), .B(n47655), .C(n47654), .D(n47653), .Y(n47662)
         );
  NAND4X1 U27446 ( .A(n47660), .B(n47659), .C(n47658), .D(n47657), .Y(n47661)
         );
  NAND4X1 U27447 ( .A(n46954), .B(n46953), .C(n46952), .D(n46951), .Y(n11389)
         );
  NAND4X1 U27448 ( .A(n45772), .B(n45771), .C(n45770), .D(n45769), .Y(n11082)
         );
  NAND4X1 U27449 ( .A(n43289), .B(n43288), .C(n43287), .D(n43286), .Y(n12006)
         );
  OR4X1 U27450 ( .A(n43607), .B(n43606), .C(n41687), .D(n41688), .Y(n12145) );
  OR2X1 U27451 ( .A(n43605), .B(n43604), .Y(n41688) );
  NAND4X1 U27452 ( .A(n43586), .B(n43585), .C(n43584), .D(n43583), .Y(n12078)
         );
  NOR2X1 U27453 ( .A(n43618), .B(n43617), .Y(n43622) );
  NAND4X1 U27454 ( .A(n43614), .B(n43613), .C(n43612), .D(n43611), .Y(n43623)
         );
  NAND2BX2 U27455 ( .AN(n39309), .B(net213731), .Y(net209898) );
  NAND2X1 U27456 ( .A(n39777), .B(net213734), .Y(n39309) );
  NOR4X1 U27457 ( .A(n45491), .B(n45490), .C(n45489), .D(n45488), .Y(net213734) );
  NAND2X1 U27458 ( .A(n39812), .B(net215915), .Y(n39328) );
  NOR2X1 U27459 ( .A(n37101), .B(n37319), .Y(n39812) );
  NAND4X1 U27460 ( .A(n43713), .B(n43712), .C(n43711), .D(n43710), .Y(n12692)
         );
  NAND2X1 U27461 ( .A(n41070), .B(net211790), .Y(n_cell_301249_net267141) );
  NAND2X1 U27462 ( .A(n41069), .B(net211785), .Y(n_cell_301249_net267135) );
  NAND4X1 U27463 ( .A(n43320), .B(n43319), .C(n43318), .D(n43317), .Y(n12479)
         );
  NAND4X1 U27464 ( .A(n43158), .B(n43157), .C(n43156), .D(n43155), .Y(n12476)
         );
  CLKINVX1 U27465 ( .A(n11697), .Y(net171198) );
  NAND4BX1 U27466 ( .AN(n41678), .B(n43266), .C(n43265), .D(n43264), .Y(n12488) );
  OR4X1 U27467 ( .A(n31389), .B(n31390), .C(n31391), .D(n31392), .Y(n41678) );
  NAND4X1 U27468 ( .A(n43284), .B(n43283), .C(n43282), .D(n43281), .Y(n12485)
         );
  CLKINVX1 U27469 ( .A(net214724), .Y(net171098) );
  CLKINVX1 U27470 ( .A(net214669), .Y(net171321) );
  NOR2X1 U27471 ( .A(n36978), .B(n37282), .Y(n40792) );
  NAND3X2 U27472 ( .A(net216515), .B(net216516), .C(n40781), .Y(n11626) );
  NOR2X1 U27473 ( .A(n36973), .B(n37264), .Y(n40781) );
  NAND3X1 U27474 ( .A(net216461), .B(net216462), .C(n40787), .Y(n11621) );
  NOR2X1 U27475 ( .A(n36979), .B(n37283), .Y(n40787) );
  NAND3X2 U27476 ( .A(net216506), .B(net216507), .C(n40775), .Y(n11625) );
  NOR2X1 U27477 ( .A(n36980), .B(n37263), .Y(n40775) );
  NAND4BX1 U27478 ( .AN(n41679), .B(n43342), .C(n43341), .D(n43340), .Y(n11657) );
  NAND4X1 U27479 ( .A(n43368), .B(n43367), .C(n43366), .D(n43365), .Y(n11652)
         );
  NAND4X1 U27480 ( .A(n43351), .B(n43350), .C(n43349), .D(n43348), .Y(n11658)
         );
  NAND4BX1 U27481 ( .AN(n41680), .B(n43359), .C(n43358), .D(n43357), .Y(n11651) );
  OR4X1 U27482 ( .A(n31058), .B(n31059), .C(n31060), .D(n31061), .Y(n41680) );
  NAND4X1 U27483 ( .A(n43395), .B(n43394), .C(n43393), .D(n43392), .Y(n12466)
         );
  NAND4X1 U27484 ( .A(n43086), .B(n43085), .C(n43084), .D(n43083), .Y(n12588)
         );
  NAND4X2 U27485 ( .A(n43377), .B(n43376), .C(n43375), .D(n43374), .Y(n11649)
         );
  NAND4X1 U27486 ( .A(n43386), .B(n43385), .C(n43384), .D(n43383), .Y(n11650)
         );
  CLKBUFX3 U27487 ( .A(n12417), .Y(net260355) );
  CLKINVX1 U27488 ( .A(net213653), .Y(net171290) );
  NAND2BX1 U27489 ( .AN(n40439), .B(net215015), .Y(net209697) );
  NAND2X1 U27490 ( .A(n40591), .B(net215018), .Y(n40439) );
  AND2X2 U27491 ( .A(net215017), .B(net215016), .Y(n40591) );
  NAND3X1 U27492 ( .A(net215062), .B(net215061), .C(net215063), .Y(
        n_cell_301249_net267948) );
  NOR2X1 U27493 ( .A(n37085), .B(n37501), .Y(n41173) );
  NOR2X1 U27494 ( .A(n37097), .B(n37456), .Y(n41127) );
  AND4X1 U27495 ( .A(n46728), .B(n46727), .C(n46726), .D(n46725), .Y(n41735)
         );
  NOR2X1 U27496 ( .A(n37075), .B(n37446), .Y(n40638) );
  NOR2X1 U27497 ( .A(n37164), .B(n37498), .Y(n40663) );
  NOR2X1 U27498 ( .A(n37142), .B(n37443), .Y(n40589) );
  NOR2X1 U27499 ( .A(n37130), .B(n37441), .Y(n40683) );
  NOR4X1 U27500 ( .A(n19698), .B(n19697), .C(n19696), .D(n19695), .Y(net211264) );
  NAND2X1 U27501 ( .A(n39903), .B(net211351), .Y(n39379) );
  NAND4X1 U27502 ( .A(n47092), .B(n47091), .C(n47090), .D(n47089), .Y(n11369)
         );
  CLKBUFX3 U27503 ( .A(n11368), .Y(n40394) );
  NAND4X1 U27504 ( .A(n47112), .B(n47111), .C(n47110), .D(n47109), .Y(n11509)
         );
  NAND4X1 U27505 ( .A(n47122), .B(n47121), .C(n47120), .D(n47119), .Y(n11360)
         );
  NOR2X1 U27506 ( .A(n37063), .B(n37485), .Y(n39913) );
  CLKBUFX3 U27507 ( .A(n13024), .Y(net260494) );
  NAND3X1 U27508 ( .A(net212146), .B(net212145), .C(net212147), .Y(
        n_cell_301249_net267343) );
  NAND3X1 U27509 ( .A(net212161), .B(net212160), .C(net212162), .Y(
        n_cell_301249_net267349) );
  NAND2X1 U27510 ( .A(n40795), .B(net212164), .Y(n11280) );
  NOR2X1 U27511 ( .A(n37379), .B(n41066), .Y(n40795) );
  NAND2X1 U27512 ( .A(net212166), .B(net212165), .Y(n41066) );
  NAND2X1 U27513 ( .A(n40413), .B(net212194), .Y(n12855) );
  NOR2X1 U27514 ( .A(n37365), .B(n40695), .Y(n40413) );
  NAND2X1 U27515 ( .A(n40414), .B(net212189), .Y(n12858) );
  NOR2X1 U27516 ( .A(n37400), .B(n40686), .Y(n40414) );
  CLKBUFX3 U27517 ( .A(n13023), .Y(net260492) );
  NOR2X1 U27518 ( .A(n37170), .B(n37447), .Y(n41162) );
  NAND3X1 U27519 ( .A(net212156), .B(net212155), .C(net212157), .Y(
        n_cell_301249_net267391) );
  NOR2X1 U27520 ( .A(n37049), .B(n37452), .Y(n41005) );
  NOR2X1 U27521 ( .A(n36974), .B(n37324), .Y(n40956) );
  NOR2X1 U27522 ( .A(n37054), .B(n37331), .Y(n41002) );
  NOR2X1 U27523 ( .A(n37050), .B(n37434), .Y(n40957) );
  NAND2X1 U27524 ( .A(net234998), .B(net214265), .Y(net210494) );
  NAND3X2 U27525 ( .A(net209617), .B(n45080), .C(n45081), .Y(net209919) );
  NOR4X1 U27526 ( .A(n45062), .B(n45061), .C(n45060), .D(n45059), .Y(n45080)
         );
  NOR4X1 U27527 ( .A(n45058), .B(n45057), .C(n45056), .D(n45055), .Y(n45081)
         );
  NAND4X1 U27528 ( .A(n44163), .B(n44162), .C(n44161), .D(n44160), .Y(
        net209873) );
  NOR4X1 U27529 ( .A(n44035), .B(n44034), .C(n44033), .D(n44032), .Y(n44036)
         );
  NAND4X1 U27530 ( .A(n44009), .B(n44008), .C(n44007), .D(n44006), .Y(
        net210677) );
  NAND2X1 U27531 ( .A(n48187), .B(n48132), .Y(net210673) );
  NOR4X1 U27532 ( .A(n27170), .B(n27169), .C(n27168), .D(n27167), .Y(n44213)
         );
  NAND4X1 U27533 ( .A(n44221), .B(n44220), .C(n44219), .D(n44218), .Y(n12744)
         );
  NAND2BX1 U27534 ( .AN(n39295), .B(net215204), .Y(n10556) );
  NAND2X1 U27535 ( .A(n39803), .B(net215207), .Y(n39295) );
  NOR2X1 U27536 ( .A(n10369), .B(n44314), .Y(net215204) );
  NOR2X1 U27537 ( .A(n37102), .B(n37310), .Y(n39803) );
  NAND2X2 U27538 ( .A(n39294), .B(net215231), .Y(n10553) );
  NOR2X1 U27539 ( .A(n37256), .B(n39804), .Y(n39294) );
  NAND2X1 U27540 ( .A(net215233), .B(net215232), .Y(n39804) );
  NOR2X1 U27541 ( .A(n37100), .B(n37308), .Y(n39297) );
  NAND2X1 U27542 ( .A(n39802), .B(net215216), .Y(n39296) );
  NOR2X1 U27543 ( .A(n36949), .B(n37333), .Y(n39802) );
  OR2X1 U27544 ( .A(net151758), .B(n39563), .Y(n39575) );
  CLKINVX1 U27545 ( .A(n12062), .Y(n39563) );
  NAND2X1 U27546 ( .A(n12049), .B(n39326), .Y(n10609) );
  NOR2X1 U27547 ( .A(n39783), .B(n39562), .Y(n39326) );
  NAND2X1 U27548 ( .A(n12152), .B(n12151), .Y(n39783) );
  CLKINVX1 U27549 ( .A(n40392), .Y(n39562) );
  NAND2X1 U27550 ( .A(n12711), .B(n12708), .Y(n10542) );
  XOR2X1 U27551 ( .A(n41948), .B(n42520), .Y(n31833) );
  NOR2X1 U27552 ( .A(n37098), .B(n37413), .Y(n40976) );
  NAND3X2 U27553 ( .A(n40777), .B(net216916), .C(net216913), .Y(n11967) );
  AND2X2 U27554 ( .A(net216915), .B(net216914), .Y(n40777) );
  NAND4X2 U27555 ( .A(n45185), .B(n45184), .C(n45183), .D(n45182), .Y(
        net209605) );
  NOR4X1 U27556 ( .A(n45179), .B(n45178), .C(n45177), .D(n45176), .Y(n45183)
         );
  NOR4X1 U27557 ( .A(n45171), .B(n45170), .C(n45169), .D(n45168), .Y(n45185)
         );
  NOR4BBX1 U27558 ( .AN(n41726), .BN(n41727), .C(n45181), .D(n45180), .Y(
        n45182) );
  OR2X1 U27559 ( .A(net210639), .B(net210635), .Y(net210426) );
  NOR2X1 U27560 ( .A(n39479), .B(net209570), .Y(n39460) );
  CLKINVX1 U27561 ( .A(n47750), .Y(n45531) );
  NOR2X1 U27562 ( .A(net171314), .B(net209638), .Y(n39464) );
  NAND4X1 U27563 ( .A(n43231), .B(n43230), .C(n43229), .D(n43228), .Y(n11673)
         );
  AND2X2 U27564 ( .A(net213222), .B(net213221), .Y(n40721) );
  NOR2X1 U27565 ( .A(n36961), .B(n37262), .Y(n40786) );
  NAND4X2 U27566 ( .A(n46364), .B(n46363), .C(n46362), .D(n46361), .Y(
        net209308) );
  AND2X4 U27567 ( .A(net209344), .B(net209313), .Y(n41763) );
  NAND4X2 U27568 ( .A(n46455), .B(n46454), .C(n46453), .D(n46452), .Y(
        net209341) );
  NAND3X1 U27569 ( .A(net209296), .B(net209300), .C(n39415), .Y(net210543) );
  NOR2X1 U27570 ( .A(net210567), .B(n39478), .Y(n39415) );
  CLKINVX1 U27571 ( .A(net209298), .Y(n39478) );
  OR2X1 U27572 ( .A(net210582), .B(net210579), .Y(net210550) );
  NAND3X1 U27573 ( .A(net209323), .B(net209320), .C(net234488), .Y(net210552)
         );
  NAND2BX2 U27574 ( .AN(n39420), .B(net209923), .Y(net210553) );
  NAND2X1 U27575 ( .A(net212213), .B(net212212), .Y(n39420) );
  NAND3BX1 U27576 ( .AN(net210581), .B(net209335), .C(net210580), .Y(net210554) );
  NAND4X1 U27577 ( .A(n44206), .B(n44205), .C(n44204), .D(n44203), .Y(n12746)
         );
  NOR2X1 U27578 ( .A(n10387), .B(n44207), .Y(n44211) );
  NAND2BX1 U27579 ( .AN(n39301), .B(net215370), .Y(n10573) );
  NAND2X1 U27580 ( .A(n39788), .B(net215373), .Y(n39301) );
  NOR2X1 U27581 ( .A(n10385), .B(n44222), .Y(net215370) );
  NOR2X1 U27582 ( .A(n36998), .B(n37223), .Y(n39788) );
  NOR4X1 U27583 ( .A(n23766), .B(n23765), .C(n23764), .D(n23763), .Y(net213360) );
  AND2X2 U27584 ( .A(net209291), .B(net209287), .Y(n41761) );
  NAND4X1 U27585 ( .A(n46231), .B(n46230), .C(n46229), .D(n46228), .Y(
        net209277) );
  OR2X1 U27586 ( .A(net210584), .B(net210559), .Y(net210528) );
  CLKINVX1 U27587 ( .A(n11148), .Y(net210531) );
  NAND2X1 U27588 ( .A(n41132), .B(net213560), .Y(n_cell_301249_net267257) );
  NOR2X1 U27589 ( .A(n37089), .B(n37506), .Y(n41132) );
  NAND2X1 U27590 ( .A(n_cell_301249_net267302), .B(net216346), .Y(n11943) );
  NOR2X1 U27591 ( .A(n37258), .B(n40988), .Y(n_cell_301249_net267302) );
  NAND2X1 U27592 ( .A(net216348), .B(net216347), .Y(n40988) );
  NAND2X1 U27593 ( .A(n37124), .B(net216364), .Y(n12803) );
  NOR2X1 U27594 ( .A(n37052), .B(n37462), .Y(n40960) );
  NOR2X1 U27595 ( .A(n37366), .B(n37143), .Y(n41130) );
  NOR2X1 U27596 ( .A(n37369), .B(n37043), .Y(n41165) );
  NOR2X1 U27597 ( .A(n37064), .B(n37417), .Y(n39829) );
  NOR2X1 U27598 ( .A(n37032), .B(n37431), .Y(n41144) );
  NAND2X1 U27599 ( .A(net213680), .B(net209623), .Y(net210476) );
  CLKINVX1 U27600 ( .A(net210665), .Y(net210475) );
  NAND2X1 U27601 ( .A(n10942), .B(n41169), .Y(n40819) );
  NOR2X1 U27602 ( .A(net171403), .B(n_cell_303546_net277738), .Y(n41169) );
  NOR2X1 U27603 ( .A(net151586), .B(net151584), .Y(n40817) );
  OR2X1 U27604 ( .A(net171390), .B(n_cell_301249_net268916), .Y(
        n_cell_301249_net269022) );
  CLKINVX1 U27605 ( .A(net211640), .Y(net171390) );
  CLKINVX1 U27606 ( .A(net209111), .Y(n_cell_301249_net268916) );
  NOR2X1 U27607 ( .A(n_cell_303546_net278017), .B(n_cell_301249_net269828),
        .Y(n41170) );
  CLKINVX1 U27608 ( .A(n10947), .Y(n_cell_301249_net269828) );
  CLKINVX1 U27609 ( .A(n10941), .Y(n_cell_301249_net269831) );
  OAI21XL U27610 ( .A0(n10632), .A1(n41107), .B0(n41108), .Y(n40849) );
  NOR2X1 U27611 ( .A(net171542), .B(net238789), .Y(n41108) );
  NAND2X1 U27612 ( .A(n10635), .B(n39341), .Y(n41107) );
  CLKINVX1 U27613 ( .A(n10630), .Y(n_cell_301249_net269745) );
  NAND2X1 U27614 ( .A(net214783), .B(net214782), .Y(n41045) );
  NOR2X1 U27615 ( .A(net171280), .B(n_cell_301249_net269646), .Y(n41046) );
  NOR2BX1 U27616 ( .AN(n11566), .B(n_cell_301249_net269647), .Y(n40871) );
  CLKINVX1 U27617 ( .A(n11565), .Y(n_cell_301249_net269647) );
  NAND2X1 U27618 ( .A(n10436), .B(n10434), .Y(n40873) );
  NOR2X1 U27619 ( .A(n41008), .B(n40900), .Y(n41009) );
  NAND2X1 U27620 ( .A(n11906), .B(n11907), .Y(n41007) );
  NOR2X1 U27621 ( .A(n40894), .B(n40899), .Y(n40898) );
  AOI21X1 U27622 ( .A0(n11904), .A1(n11897), .B0(n41010), .Y(n40902) );
  NAND2X1 U27623 ( .A(n11902), .B(n11901), .Y(n41010) );
  NAND2X1 U27624 ( .A(n11895), .B(n11896), .Y(n40904) );
  NAND2X1 U27625 ( .A(net234521), .B(net234523), .Y(n39642) );
  OR2X1 U27626 ( .A(net210598), .B(net210596), .Y(net210516) );
  OR2X1 U27627 ( .A(net210601), .B(net210618), .Y(net210520) );
  AOI21X1 U27628 ( .A0(net171290), .A1(net209697), .B0(n40746), .Y(n40747) );
  NAND2X1 U27629 ( .A(n11901), .B(n11895), .Y(n40746) );
  NAND2X1 U27630 ( .A(n11896), .B(n11894), .Y(n40748) );
  NOR2X1 U27631 ( .A(n40583), .B(n11902), .Y(n40582) );
  CLKINVX1 U27632 ( .A(n11895), .Y(n40583) );
  CLKINVX1 U27633 ( .A(n11893), .Y(n40749) );
  NAND2X1 U27634 ( .A(n40766), .B(net214756), .Y(n40509) );
  OAI21XL U27635 ( .A0(n40506), .A1(n40631), .B0(n40632), .Y(n40766) );
  OAI21XL U27636 ( .A0(n_cell_303546_net277490), .A1(n10434), .B0(n40630), .Y(
        n40631) );
  OA21XL U27637 ( .A0(net151380), .A1(n10292), .B0(net272620), .Y(n40632) );
  NOR4X1 U27638 ( .A(n_cell_303546_net277804), .B(n40579), .C(n40710), .D(
        net151790), .Y(n40709) );
  NOR2X1 U27639 ( .A(n39927), .B(n10759), .Y(n40579) );
  NOR2X1 U27640 ( .A(net171542), .B(net151809), .Y(n40715) );
  CLKINVX1 U27641 ( .A(n39341), .Y(n_cell_303546_net277814) );
  NAND2X1 U27642 ( .A(n40685), .B(net210356), .Y(n40436) );
  NOR2X1 U27643 ( .A(n37028), .B(n37422), .Y(n40685) );
  NAND3X1 U27644 ( .A(n39341), .B(n40713), .C(n40714), .Y(n40712) );
  NAND2BX1 U27645 ( .AN(net260461), .B(net209996), .Y(n40714) );
  NOR2X1 U27646 ( .A(n40710), .B(n_cell_301249_net269738), .Y(n40711) );
  NOR2X1 U27647 ( .A(n37152), .B(n37487), .Y(n40590) );
  NOR2X1 U27648 ( .A(n40669), .B(n40577), .Y(n40556) );
  NAND3X1 U27649 ( .A(n10938), .B(net272417), .C(net260830), .Y(n40669) );
  NOR2X1 U27650 ( .A(n_cell_301249_net269836), .B(n10941), .Y(n40577) );
  NAND3X1 U27651 ( .A(n40670), .B(n40672), .C(n40673), .Y(n40557) );
  NAND2BX1 U27652 ( .AN(net209101), .B(net272417), .Y(n40672) );
  NOR2X1 U27653 ( .A(net171394), .B(n40671), .Y(n40670) );
  NAND3BX1 U27654 ( .AN(net211602), .B(net260830), .C(net272417), .Y(n40673)
         );
  NAND2X1 U27655 ( .A(net171392), .B(n12196), .Y(n40675) );
  NAND2X1 U27656 ( .A(n10776), .B(n10771), .Y(n40676) );
  NOR2X1 U27657 ( .A(n37135), .B(n37494), .Y(n40598) );
  AOI21X1 U27658 ( .A0(n39608), .A1(n39609), .B0(n10143), .Y(n39607) );
  NOR4X1 U27659 ( .A(net151542), .B(n_cell_303546_net277630), .C(n39606), .D(
        n_cell_303546_net277834), .Y(n39609) );
  OAI21XL U27660 ( .A0(n39830), .A1(n39603), .B0(n40026), .Y(n39608) );
  CLKINVX1 U27661 ( .A(n_cell_303546_net275967), .Y(n39606) );
  CLKINVX1 U27662 ( .A(n10611), .Y(n40022) );
  CLKINVX1 U27663 ( .A(n11915), .Y(n39835) );
  AND2X2 U27664 ( .A(net259665), .B(net259661), .Y(n39866) );
  OAI21XL U27665 ( .A0(n10311), .A1(n39471), .B0(net168848), .Y(n39760) );
  AOI21X1 U27666 ( .A0(n39472), .A1(n39473), .B0(n39474), .Y(n39471) );
  NAND2X1 U27667 ( .A(n39861), .B(net260900), .Y(n39474) );
  NOR2X1 U27668 ( .A(n39860), .B(net151283), .Y(n39473) );
  NAND2X1 U27669 ( .A(net261422), .B(n39864), .Y(n39761) );
  NOR2X1 U27670 ( .A(net151299), .B(n39863), .Y(n39864) );
  NAND2X1 U27671 ( .A(net259626), .B(n10302), .Y(n39863) );
  OAI21XL U27672 ( .A0(n39530), .A1(n39988), .B0(n39990), .Y(n39534) );
  NAND2X1 U27673 ( .A(n10903), .B(n39989), .Y(n39988) );
  NOR4BX1 U27674 ( .AN(n10801), .B(n39991), .C(n39532), .D(net171480), .Y(
        n39990) );
  NOR2X1 U27675 ( .A(n39527), .B(n39531), .Y(n39530) );
  NOR2X1 U27676 ( .A(n39992), .B(net171398), .Y(n39535) );
  NAND3X1 U27677 ( .A(n_cell_303546_net275923), .B(n_cell_303546_net275959),
        .C(n10983), .Y(n39992) );
  NAND3X1 U27678 ( .A(net259873), .B(net271956), .C(n39993), .Y(n39536) );
  NOR2X1 U27679 ( .A(net171401), .B(net151536), .Y(n39993) );
  NAND2X1 U27680 ( .A(n40586), .B(net211629), .Y(n40713) );
  NOR2X1 U27681 ( .A(n37376), .B(n40585), .Y(n40586) );
  OAI21XL U27682 ( .A0(n39681), .A1(n39683), .B0(n39922), .Y(n39687) );
  NOR2X1 U27683 ( .A(n39923), .B(n39685), .Y(n39922) );
  NOR2X1 U27684 ( .A(n39678), .B(n39682), .Y(n39681) );
  NAND2X1 U27685 ( .A(n39921), .B(n11280), .Y(n39682) );
  CLKINVX1 U27686 ( .A(n9900), .Y(n39688) );
  CLKINVX1 U27687 ( .A(n39342), .Y(n_cell_303546_net277636) );
  CLKINVX1 U27688 ( .A(n10759), .Y(n39928) );
  CLKINVX1 U27689 ( .A(n10641), .Y(n39925) );
  NOR2X1 U27690 ( .A(n37489), .B(n37180), .Y(n41119) );
  NAND2BX1 U27691 ( .AN(n39401), .B(net212731), .Y(n10845) );
  NAND2X1 U27692 ( .A(n39967), .B(net212734), .Y(n39401) );
  NOR2X1 U27693 ( .A(n37167), .B(n37405), .Y(n39967) );
  NAND2BX2 U27694 ( .AN(n39402), .B(net213422), .Y(n10843) );
  NAND2X1 U27695 ( .A(n39966), .B(net213423), .Y(n39402) );
  NOR2X1 U27696 ( .A(n45638), .B(net209814), .Y(net213422) );
  NAND3X1 U27697 ( .A(n12311), .B(n12386), .C(n39403), .Y(n10842) );
  NOR2X1 U27698 ( .A(n39493), .B(n39494), .Y(n39403) );
  CLKINVX1 U27699 ( .A(n40396), .Y(n39494) );
  CLKINVX1 U27700 ( .A(n11204), .Y(n39493) );
  NAND2BX2 U27701 ( .AN(n39400), .B(net212741), .Y(n10846) );
  NAND2X1 U27702 ( .A(n39968), .B(net212744), .Y(n39400) );
  NOR2X1 U27703 ( .A(n12717), .B(n46168), .Y(net212741) );
  NAND2BX1 U27704 ( .AN(n39399), .B(net212736), .Y(n10847) );
  NAND2X1 U27705 ( .A(n39969), .B(net212739), .Y(n39399) );
  NOR2X1 U27706 ( .A(n37168), .B(n37409), .Y(n39969) );
  NAND4X1 U27707 ( .A(n46142), .B(n46141), .C(n46140), .D(n46139), .Y(n12385)
         );
  NOR2X1 U27708 ( .A(n22391), .B(n22390), .Y(n46140) );
  NAND3X1 U27709 ( .A(n12333), .B(n12384), .C(n39409), .Y(n10865) );
  NOR2X1 U27710 ( .A(net209362), .B(n39495), .Y(n39409) );
  CLKINVX1 U27711 ( .A(n11201), .Y(n39495) );
  NAND2BX1 U27712 ( .AN(n39436), .B(net213115), .Y(n10243) );
  NAND2X1 U27713 ( .A(n39944), .B(net213116), .Y(n39436) );
  NOR2X1 U27714 ( .A(n37059), .B(n37318), .Y(n39944) );
  NOR2X1 U27715 ( .A(n23218), .B(n23217), .Y(n45830) );
  NOR4X1 U27716 ( .A(n23216), .B(n23215), .C(n23214), .D(n23213), .Y(n45829)
         );
  NAND4X1 U27717 ( .A(n45827), .B(n45826), .C(n45825), .D(n45824), .Y(n11211)
         );
  NOR2X1 U27718 ( .A(n23228), .B(n23227), .Y(n45825) );
  NAND4X1 U27719 ( .A(n45837), .B(n45836), .C(n45835), .D(n45834), .Y(n12292)
         );
  NAND4X1 U27720 ( .A(n45812), .B(n45811), .C(n45810), .D(n45809), .Y(n11072)
         );
  CLKINVX1 U27721 ( .A(net209202), .Y(net171456) );
  CLKINVX1 U27722 ( .A(n12287), .Y(net151662) );
  CLKINVX1 U27723 ( .A(n39730), .Y(n10362) );
  NAND4X1 U27724 ( .A(n44537), .B(n44536), .C(n44535), .D(n44534), .Y(n11709)
         );
  NOR4X1 U27725 ( .A(n24814), .B(n24815), .C(n24816), .D(n24817), .Y(n44543)
         );
  NOR4X1 U27726 ( .A(n24806), .B(n24807), .C(n24808), .D(n24809), .Y(n44545)
         );
  NOR4X1 U27727 ( .A(n24810), .B(n24811), .C(n24812), .D(n24813), .Y(n44544)
         );
  NAND4X1 U27728 ( .A(n44564), .B(n44563), .C(n44562), .D(n44561), .Y(n11710)
         );
  CLKINVX1 U27729 ( .A(n39732), .Y(n10355) );
  NAND2BX1 U27730 ( .AN(net171301), .B(n39733), .Y(n39732) );
  NOR3X1 U27731 ( .A(net151394), .B(net171305), .C(net209509), .Y(n39733) );
  NAND3X1 U27732 ( .A(n11722), .B(n12585), .C(n11721), .Y(n10357) );
  CLKINVX1 U27733 ( .A(net209503), .Y(net171300) );
  NOR4X1 U27734 ( .A(n28512), .B(n28513), .C(n28514), .D(n28515), .Y(n43696)
         );
  NAND4X1 U27735 ( .A(n43790), .B(n43789), .C(n43788), .D(n43787), .Y(n11705)
         );
  NOR4X1 U27736 ( .A(n28182), .B(n28183), .C(n28184), .D(n28185), .Y(n43787)
         );
  NAND4X1 U27737 ( .A(n43772), .B(n43771), .C(n43770), .D(n43769), .Y(n11700)
         );
  NAND4X1 U27738 ( .A(n43690), .B(n43689), .C(n43688), .D(n43687), .Y(n12501)
         );
  NOR4X1 U27739 ( .A(n28542), .B(n28543), .C(n28544), .D(n28545), .Y(n43687)
         );
  NAND4X1 U27740 ( .A(n43763), .B(n43762), .C(n43761), .D(n43760), .Y(n12587)
         );
  NAND4X1 U27741 ( .A(n43681), .B(n43680), .C(n43679), .D(n43678), .Y(n11698)
         );
  NAND4X1 U27742 ( .A(n43717), .B(n43716), .C(n43715), .D(n43714), .Y(n11685)
         );
  NAND4X1 U27743 ( .A(n43726), .B(n43725), .C(n43724), .D(n43723), .Y(n11686)
         );
  NAND4X1 U27744 ( .A(n43749), .B(n43748), .C(n43747), .D(n43746), .Y(n11694)
         );
  NAND4X1 U27745 ( .A(n43708), .B(n43707), .C(n43706), .D(n43705), .Y(n11687)
         );
  NOR2X1 U27746 ( .A(n36954), .B(n37212), .Y(n39455) );
  NAND3X2 U27747 ( .A(net216025), .B(net216026), .C(n39454), .Y(n10378) );
  NOR2X1 U27748 ( .A(n37230), .B(n36995), .Y(n39454) );
  NOR4X1 U27749 ( .A(n29286), .B(n29287), .C(n29288), .D(n29289), .Y(net216026) );
  NAND3X1 U27750 ( .A(n11763), .B(n39466), .C(n12538), .Y(n10420) );
  NOR2X1 U27751 ( .A(n39722), .B(net171189), .Y(n39466) );
  CLKINVX1 U27752 ( .A(n11762), .Y(n39722) );
  NOR4X1 U27753 ( .A(n26789), .B(n26790), .C(n26791), .D(n26792), .Y(n44280)
         );
  NAND4BX1 U27754 ( .AN(n41668), .B(n43663), .C(n43662), .D(n43661), .Y(n11849) );
  OR4X1 U27755 ( .A(n29041), .B(n29042), .C(n29043), .D(n29044), .Y(n41668) );
  NOR4X1 U27756 ( .A(n29474), .B(n29475), .C(n29476), .D(n29477), .Y(n43546)
         );
  NOR4X1 U27757 ( .A(n29444), .B(n29445), .C(n29446), .D(n29447), .Y(n43555)
         );
  NAND4BX1 U27758 ( .AN(n41677), .B(n43655), .C(n43654), .D(n43653), .Y(n11752) );
  OR4X1 U27759 ( .A(n29071), .B(n29072), .C(n29073), .D(n29074), .Y(n41677) );
  NAND4X1 U27760 ( .A(n47232), .B(n47231), .C(n47230), .D(n47229), .Y(n11422)
         );
  NAND4X1 U27761 ( .A(n47237), .B(n47236), .C(n47235), .D(n47234), .Y(n11423)
         );
  NAND4X1 U27762 ( .A(n47143), .B(n47142), .C(n47141), .D(n47140), .Y(n11414)
         );
  NAND4X1 U27763 ( .A(n47148), .B(n47147), .C(n47146), .D(n47145), .Y(n11415)
         );
  NOR2X1 U27764 ( .A(n19831), .B(n19830), .Y(n47146) );
  NAND3X1 U27765 ( .A(net211474), .B(net211476), .C(net211475), .Y(n39363) );
  NOR2X1 U27766 ( .A(n40397), .B(n47044), .Y(net211473) );
  NAND2BX1 U27767 ( .AN(n39362), .B(net211478), .Y(n10724) );
  NAND3X1 U27768 ( .A(net211480), .B(net211479), .C(net211481), .Y(n39362) );
  NAND2X1 U27769 ( .A(n39886), .B(net211516), .Y(n39367) );
  NAND2BX1 U27770 ( .AN(n39369), .B(net211523), .Y(n10730) );
  NAND2X1 U27771 ( .A(n39884), .B(net211526), .Y(n39369) );
  NAND2BX1 U27772 ( .AN(n39366), .B(net211518), .Y(n10734) );
  NAND2X1 U27773 ( .A(n39887), .B(net211521), .Y(n39366) );
  NAND2BX2 U27774 ( .AN(n39368), .B(net211508), .Y(n10732) );
  NAND2X1 U27775 ( .A(n39885), .B(net211511), .Y(n39368) );
  NAND4X1 U27776 ( .A(n12976), .B(n13014), .C(n11441), .D(n11442), .Y(n10729)
         );
  NAND4X1 U27777 ( .A(n46924), .B(n46923), .C(n46922), .D(n46921), .Y(n11379)
         );
  NAND4X1 U27778 ( .A(n46919), .B(n46918), .C(n46917), .D(n46916), .Y(n11378)
         );
  NOR2X1 U27779 ( .A(n21112), .B(n21111), .Y(n46912) );
  NOR4X1 U27780 ( .A(n21110), .B(n21109), .C(n21108), .D(n21107), .Y(n46911)
         );
  NAND3X1 U27781 ( .A(net211642), .B(net211644), .C(net211643), .Y(n39376) );
  NAND3X1 U27782 ( .A(net211652), .B(net211654), .C(net211653), .Y(n39377) );
  NAND2BX1 U27783 ( .AN(n39378), .B(net211657), .Y(n10751) );
  NAND3X1 U27784 ( .A(net211658), .B(net211660), .C(net211659), .Y(n39378) );
  CLKINVX1 U27785 ( .A(net211667), .Y(net171540) );
  NAND3X1 U27786 ( .A(n39355), .B(n11389), .C(n11386), .Y(n10699) );
  NOR2X1 U27787 ( .A(n39637), .B(n39636), .Y(n39355) );
  CLKINVX1 U27788 ( .A(n11387), .Y(n39637) );
  NAND4X1 U27789 ( .A(n45732), .B(n45731), .C(n45730), .D(n45729), .Y(n11208)
         );
  NAND3X1 U27790 ( .A(n12006), .B(n12007), .C(n39590), .Y(n39589) );
  NOR2X1 U27791 ( .A(n39557), .B(net171127), .Y(n39590) );
  OR4X1 U27792 ( .A(net171125), .B(net171126), .C(net171122), .D(net171124),
        .Y(n39592) );
  NAND4X1 U27793 ( .A(n43209), .B(n43208), .C(n43207), .D(n43206), .Y(n12156)
         );
  NAND4X1 U27794 ( .A(n43200), .B(n43199), .C(n43198), .D(n43197), .Y(n12157)
         );
  NAND4X1 U27795 ( .A(n43227), .B(n43226), .C(n43225), .D(n43224), .Y(n12015)
         );
  NAND4X1 U27796 ( .A(n43218), .B(n43217), .C(n43216), .D(n43215), .Y(n12014)
         );
  NAND2X1 U27797 ( .A(n39787), .B(net216050), .Y(n39299) );
  NOR2X1 U27798 ( .A(n37107), .B(n37313), .Y(n39787) );
  NOR2X1 U27799 ( .A(net209956), .B(n39565), .Y(n39300) );
  CLKINVX1 U27800 ( .A(n12078), .Y(n39565) );
  NAND2X1 U27801 ( .A(n37255), .B(n43677), .Y(n12065) );
  NOR2X1 U27802 ( .A(n12530), .B(n43673), .Y(n43677) );
  NAND4X1 U27803 ( .A(n43652), .B(n43651), .C(n43650), .D(n43649), .Y(n12795)
         );
  OR3X2 U27804 ( .A(n41685), .B(n41686), .C(net209635), .Y(net209902) );
  OR4X1 U27805 ( .A(n45416), .B(n45415), .C(n45414), .D(n45413), .Y(n41686) );
  OR4X1 U27806 ( .A(n45412), .B(n45411), .C(n45410), .D(n45409), .Y(n41685) );
  NAND4X2 U27807 ( .A(n45465), .B(n45464), .C(n45463), .D(n45462), .Y(
        net209903) );
  NOR2X1 U27808 ( .A(n45455), .B(net209606), .Y(n45465) );
  NOR4X1 U27809 ( .A(n45461), .B(n45460), .C(n45459), .D(n45458), .Y(n45462)
         );
  NAND2X1 U27810 ( .A(net234529), .B(net213824), .Y(net210490) );
  NAND2X1 U27811 ( .A(n12639), .B(n12643), .Y(n_cell_301249_net269449) );
  NAND4X1 U27812 ( .A(n43786), .B(n43785), .C(n43784), .D(n43783), .Y(n12154)
         );
  NOR2X1 U27813 ( .A(n28195), .B(n28194), .Y(n43784) );
  NOR4X1 U27814 ( .A(n28193), .B(n28192), .C(n28191), .D(n28190), .Y(n43783)
         );
  NOR2X1 U27815 ( .A(n39560), .B(net209791), .Y(n39291) );
  NAND4X1 U27816 ( .A(n46763), .B(n46762), .C(n46761), .D(n46760), .Y(n11348)
         );
  NAND4X1 U27817 ( .A(n46773), .B(n46772), .C(n46771), .D(n46770), .Y(n11349)
         );
  NAND4X1 U27818 ( .A(n46758), .B(n46757), .C(n46756), .D(n46755), .Y(n11511)
         );
  NAND4X1 U27819 ( .A(n46748), .B(n46747), .C(n46746), .D(n46745), .Y(n11512)
         );
  NAND4X1 U27820 ( .A(n46718), .B(n46717), .C(n46716), .D(n46715), .Y(n11350)
         );
  NAND4X1 U27821 ( .A(n46723), .B(n46722), .C(n46721), .D(n46720), .Y(n11351)
         );
  OR3X2 U27822 ( .A(net151465), .B(net151467), .C(n37344), .Y(n39665) );
  NOR2X1 U27823 ( .A(n37129), .B(n37404), .Y(n39878) );
  NOR2X1 U27824 ( .A(n37133), .B(n37445), .Y(n39876) );
  NOR2X1 U27825 ( .A(n37159), .B(n37401), .Y(n39877) );
  NOR2X1 U27826 ( .A(n37371), .B(n37145), .Y(n41089) );
  NOR2X1 U27827 ( .A(n37368), .B(n37148), .Y(n41067) );
  CLKINVX1 U27828 ( .A(n11291), .Y(n39676) );
  NAND2BX1 U27829 ( .AN(n_cell_301249_net267219), .B(net210621), .Y(n11520) );
  NAND2X1 U27830 ( .A(n41088), .B(net210623), .Y(n_cell_301249_net267219) );
  NOR2X1 U27831 ( .A(n37153), .B(n37484), .Y(n41058) );
  CLKBUFX3 U27832 ( .A(n12590), .Y(net260376) );
  NOR2X1 U27833 ( .A(n36993), .B(n37297), .Y(n_cell_301249_net267447) );
  NOR2X1 U27834 ( .A(n37070), .B(n37298), .Y(n_cell_301249_net267441) );
  NAND4X1 U27835 ( .A(n43121), .B(n43120), .C(n43119), .D(n43118), .Y(n11637)
         );
  NAND4X1 U27836 ( .A(n43149), .B(n43148), .C(n43147), .D(n43146), .Y(n11638)
         );
  NAND4BX1 U27837 ( .AN(n41681), .B(n43094), .C(n43093), .D(n43092), .Y(n11645) );
  OR4X1 U27838 ( .A(n32141), .B(n32142), .C(n32143), .D(n32144), .Y(n41681) );
  NAND4X1 U27839 ( .A(n43103), .B(n43102), .C(n43101), .D(n43100), .Y(n11646)
         );
  NAND4X1 U27840 ( .A(n43135), .B(n43134), .C(n43133), .D(n43132), .Y(n11640)
         );
  NAND4X1 U27841 ( .A(n43112), .B(n43111), .C(n43110), .D(n43109), .Y(n11639)
         );
  CLKINVX1 U27842 ( .A(n11688), .Y(net171207) );
  NAND2X1 U27843 ( .A(n12488), .B(n12485), .Y(n10094) );
  NAND2X1 U27844 ( .A(net216264), .B(net216263), .Y(n40421) );
  NOR2X1 U27845 ( .A(n37069), .B(n37295), .Y(n_cell_301249_net267510) );
  NAND2X1 U27846 ( .A(net216273), .B(net216272), .Y(n40419) );
  NOR2X1 U27847 ( .A(n36991), .B(n37294), .Y(n_cell_301249_net267516) );
  NOR2X1 U27848 ( .A(n36964), .B(n37265), .Y(n_cell_301249_net267589) );
  NAND2X1 U27849 ( .A(n39751), .B(n39752), .Y(n39750) );
  NOR2X1 U27850 ( .A(net171098), .B(net151246), .Y(n39751) );
  NOR2X1 U27851 ( .A(net171321), .B(net151243), .Y(n39752) );
  CLKBUFX3 U27852 ( .A(n10427), .Y(net259645) );
  NAND3X1 U27853 ( .A(n11626), .B(n11621), .C(n39445), .Y(n10331) );
  NOR2X1 U27854 ( .A(n39702), .B(n39703), .Y(n39445) );
  CLKINVX1 U27855 ( .A(n11625), .Y(n39703) );
  NAND2BX2 U27856 ( .AN(n39469), .B(n_cell_301249_net267095), .Y(n10425) );
  NOR2X1 U27857 ( .A(n36960), .B(n37279), .Y(n_cell_301249_net267095) );
  NAND2X1 U27858 ( .A(net216471), .B(net216470), .Y(n39469) );
  NAND4X1 U27859 ( .A(n11657), .B(n11658), .C(n11651), .D(n11652), .Y(n10338)
         );
  NAND4X1 U27860 ( .A(n11649), .B(n11650), .C(n12466), .D(n12588), .Y(n10334)
         );
  CLKINVX1 U27861 ( .A(net260355), .Y(net151373) );
  NOR2BX1 U27862 ( .AN(net215116), .B(n37361), .Y(n40952) );
  NAND3X1 U27863 ( .A(n10526), .B(n10527), .C(n10525), .Y(n10152) );
  NAND2BX1 U27864 ( .AN(n40433), .B(net215051), .Y(n12611) );
  NAND3X1 U27865 ( .A(net215053), .B(net215052), .C(net215054), .Y(n40433) );
  NAND2BX1 U27866 ( .AN(n40435), .B(net215042), .Y(n12614) );
  NAND2X1 U27867 ( .A(n40722), .B(net215045), .Y(n40435) );
  AND2X2 U27868 ( .A(net215044), .B(net215043), .Y(n40722) );
  CLKBUFX3 U27869 ( .A(n12618), .Y(net260403) );
  NAND2BX1 U27870 ( .AN(net171290), .B(net209697), .Y(n40900) );
  NAND2BX1 U27871 ( .AN(n_cell_301249_net267319), .B(net213517), .Y(n10969) );
  NAND2X1 U27872 ( .A(n41159), .B(net213520), .Y(n_cell_301249_net267319) );
  NAND2BX1 U27873 ( .AN(n_cell_301249_net267337), .B(net213512), .Y(n10965) );
  NAND2X1 U27874 ( .A(n41161), .B(net213515), .Y(n_cell_301249_net267337) );
  AND2X2 U27875 ( .A(net212080), .B(net212079), .Y(n40639) );
  NAND2X1 U27876 ( .A(n41128), .B(net213621), .Y(n_cell_301249_net267706) );
  CLKINVX1 U27877 ( .A(n_cell_301249_net269022), .Y(n10942) );
  NAND2BX1 U27878 ( .AN(n40432), .B(net212104), .Y(n12838) );
  NAND3X1 U27879 ( .A(net212106), .B(net212105), .C(net212107), .Y(n40432) );
  NAND2BX1 U27880 ( .AN(n40430), .B(net212114), .Y(n12840) );
  NAND3X1 U27881 ( .A(net212116), .B(net212115), .C(net212117), .Y(n40430) );
  NOR2X1 U27882 ( .A(n37131), .B(n37410), .Y(n41060) );
  NAND2BX1 U27883 ( .AN(n40947), .B(net211635), .Y(n_cell_301249_net269738) );
  NAND2X1 U27884 ( .A(n40946), .B(net211637), .Y(n40947) );
  CLKBUFX3 U27885 ( .A(n12831), .Y(net260461) );
  CLKINVX1 U27886 ( .A(n12834), .Y(net151790) );
  NAND3X1 U27887 ( .A(net211258), .B(net211257), .C(net211259), .Y(n39356) );
  NAND2BX1 U27888 ( .AN(n39357), .B(net211251), .Y(n10709) );
  NAND3X1 U27889 ( .A(net211253), .B(net211252), .C(net211254), .Y(n39357) );
  NOR2X1 U27890 ( .A(n10854), .B(n47216), .Y(net211251) );
  NAND2BX1 U27891 ( .AN(n39359), .B(net211261), .Y(n10706) );
  NAND3X1 U27892 ( .A(net211263), .B(net211262), .C(net211264), .Y(n39359) );
  NAND2BX1 U27893 ( .AN(n39358), .B(net211246), .Y(n10708) );
  NAND3X1 U27894 ( .A(net211248), .B(net211247), .C(net211249), .Y(n39358) );
  NAND3X1 U27895 ( .A(n11410), .B(n11411), .C(n39360), .Y(n10705) );
  NOR2X1 U27896 ( .A(n39638), .B(n36944), .Y(n39360) );
  CLKINVX1 U27897 ( .A(n13016), .Y(n39638) );
  CLKINVX1 U27898 ( .A(n39647), .Y(n10719) );
  CLKBUFX3 U27899 ( .A(n13021), .Y(net260488) );
  NAND2BX1 U27900 ( .AN(n40784), .B(net211967), .Y(n11301) );
  NAND3X1 U27901 ( .A(net211969), .B(net211968), .C(net211970), .Y(n40784) );
  NAND2BX1 U27902 ( .AN(n40785), .B(net211972), .Y(n11300) );
  NAND3X1 U27903 ( .A(net211974), .B(net211973), .C(net211975), .Y(n40785) );
  CLKBUFX3 U27904 ( .A(n10013), .Y(n40405) );
  CLKINVX1 U27905 ( .A(n11315), .Y(net171534) );
  CLKINVX1 U27906 ( .A(n11314), .Y(net171533) );
  NAND3X1 U27907 ( .A(n11316), .B(n11317), .C(n39349), .Y(n10671) );
  NOR2X1 U27908 ( .A(n36943), .B(n39626), .Y(n39349) );
  NAND2X1 U27909 ( .A(net210043), .B(n41191), .Y(n_cell_301249_net269861) );
  CLKINVX1 U27910 ( .A(net238868), .Y(n41191) );
  NAND3X1 U27911 ( .A(n12856), .B(net260494), .C(n39684), .Y(n39683) );
  NOR2X1 U27912 ( .A(n39621), .B(n39622), .Y(n39684) );
  OR2X1 U27913 ( .A(net151554), .B(n37352), .Y(n39685) );
  CLKINVX1 U27914 ( .A(n11280), .Y(net171524) );
  NAND3X1 U27915 ( .A(n_cell_303546_net276009), .B(n39344), .C(net260492), .Y(
        n10651) );
  NOR2X1 U27916 ( .A(n39623), .B(n_cell_303546_net277530), .Y(n39344) );
  NAND2X1 U27917 ( .A(n41063), .B(net212020), .Y(n_cell_301249_net267574) );
  NOR2X1 U27918 ( .A(n37139), .B(n37402), .Y(n41063) );
  NOR2X1 U27919 ( .A(n37482), .B(n37172), .Y(n41064) );
  NAND2BX2 U27920 ( .AN(n40443), .B(net213592), .Y(n12196) );
  NAND2X1 U27921 ( .A(n40637), .B(net213595), .Y(n40443) );
  NOR2X1 U27922 ( .A(n37163), .B(n37497), .Y(n40637) );
  NOR2X1 U27923 ( .A(n37477), .B(n37177), .Y(n41059) );
  NAND2X1 U27924 ( .A(n39338), .B(n12640), .Y(n10610) );
  NOR2X1 U27925 ( .A(n39605), .B(n39782), .Y(n39338) );
  NAND2X1 U27926 ( .A(n12803), .B(n11943), .Y(n39782) );
  NAND2X1 U27927 ( .A(n40965), .B(net216338), .Y(n_cell_301249_net267385) );
  NAND2X1 U27928 ( .A(n40963), .B(net216320), .Y(n_cell_301249_net267397) );
  NAND2X1 U27929 ( .A(n40964), .B(net216329), .Y(n_cell_301249_net267379) );
  CLKINVX1 U27930 ( .A(n12804), .Y(n39553) );
  CLKINVX1 U27931 ( .A(n11935), .Y(n39554) );
  NAND2X1 U27932 ( .A(n37121), .B(net216310), .Y(n11934) );
  NAND2BX1 U27933 ( .AN(n_cell_301249_net267550), .B(net216247), .Y(n12166) );
  NAND3X1 U27934 ( .A(net216249), .B(net216248), .C(net216250), .Y(
        n_cell_301249_net267550) );
  CLKINVX1 U27935 ( .A(n11933), .Y(n_cell_301249_net269578) );
  CLKBUFX3 U27936 ( .A(n12624), .Y(net271996) );
  NAND3X1 U27937 ( .A(net209900), .B(net210695), .C(net214016), .Y(n39568) );
  OR2X1 U27938 ( .A(net210699), .B(n39310), .Y(net210441) );
  NAND2X1 U27939 ( .A(net209919), .B(net258199), .Y(n39310) );
  CLKINVX1 U27940 ( .A(n39571), .Y(net234760) );
  NAND2BX2 U27941 ( .AN(n39303), .B(net215831), .Y(n10184) );
  NAND2X1 U27942 ( .A(n39789), .B(net215834), .Y(n39303) );
  NOR2X1 U27943 ( .A(n36999), .B(n37227), .Y(n39789) );
  NAND2X1 U27944 ( .A(n39312), .B(net209873), .Y(net210445) );
  NOR2X1 U27945 ( .A(net210680), .B(net209885), .Y(n39312) );
  OR2X1 U27946 ( .A(net210675), .B(n39306), .Y(net210444) );
  CLKINVX1 U27947 ( .A(n10182), .Y(net171222) );
  NOR2X1 U27948 ( .A(n10128), .B(n43819), .Y(net215822) );
  NAND2X1 U27949 ( .A(n39790), .B(net215825), .Y(n39305) );
  CLKINVX1 U27950 ( .A(n10573), .Y(net171240) );
  NAND3X1 U27951 ( .A(net215361), .B(net215362), .C(n39316), .Y(n10567) );
  NOR2X1 U27952 ( .A(n36977), .B(n37225), .Y(n39316) );
  NOR2X1 U27953 ( .A(n36976), .B(n37224), .Y(n39317) );
  CLKINVX1 U27954 ( .A(n39580), .Y(n10548) );
  NAND2X1 U27955 ( .A(n12036), .B(n12041), .Y(n10169) );
  NAND3X1 U27956 ( .A(n12034), .B(n12035), .C(n39292), .Y(n10170) );
  NOR2X1 U27957 ( .A(net171313), .B(n39561), .Y(n39292) );
  NAND2X1 U27958 ( .A(n40961), .B(net216239), .Y(n_cell_301249_net267619) );
  NOR2X1 U27959 ( .A(n36989), .B(n37292), .Y(n40798) );
  NAND3X1 U27960 ( .A(n40425), .B(net216210), .C(net216207), .Y(n12424) );
  NOR2X1 U27961 ( .A(n37066), .B(n37382), .Y(n40425) );
  NOR2X1 U27962 ( .A(n37073), .B(n37463), .Y(n40958) );
  NAND3X1 U27963 ( .A(n40424), .B(net214781), .C(net214778), .Y(n12427) );
  NOR2X1 U27964 ( .A(n37067), .B(n37285), .Y(n40424) );
  NOR2X1 U27965 ( .A(n37109), .B(n37312), .Y(n39337) );
  CLKINVX1 U27966 ( .A(n39288), .Y(net151430) );
  NAND4BX1 U27967 ( .AN(n39289), .B(n11976), .C(n11978), .D(n11979), .Y(n39288) );
  NOR2X1 U27968 ( .A(n36962), .B(n37259), .Y(n40427) );
  NAND3X4 U27969 ( .A(net214759), .B(n_cell_301249_net267780), .C(net214758),
        .Y(n11578) );
  NOR2X1 U27970 ( .A(n37047), .B(n37270), .Y(n_cell_301249_net267780) );
  NAND3X2 U27971 ( .A(net214763), .B(n_cell_301249_net267867), .C(net214762),
        .Y(n11575) );
  NOR2X1 U27972 ( .A(n36968), .B(n37269), .Y(n_cell_301249_net267867) );
  NAND3X1 U27973 ( .A(net216217), .B(n_cell_301249_net267601), .C(net216216),
        .Y(n11869) );
  NOR2X1 U27974 ( .A(n37048), .B(n37271), .Y(n_cell_301249_net267601) );
  NAND2X1 U27975 ( .A(n12427), .B(n12424), .Y(n11584) );
  NAND2X1 U27976 ( .A(n39462), .B(net209635), .Y(net210390) );
  NOR2BX1 U27977 ( .AN(net209605), .B(net210660), .Y(n39462) );
  CLKINVX1 U27978 ( .A(n11770), .Y(net151349) );
  CLKINVX1 U27979 ( .A(n40393), .Y(net151347) );
  NAND3X2 U27980 ( .A(net216758), .B(net216759), .C(n39448), .Y(n10339) );
  NOR2X1 U27981 ( .A(n36958), .B(n37216), .Y(n39448) );
  NAND3X1 U27982 ( .A(net216749), .B(net216750), .C(n39449), .Y(n10336) );
  NOR2X1 U27983 ( .A(n36957), .B(n37277), .Y(n39449) );
  NAND3X1 U27984 ( .A(net214662), .B(net214663), .C(n39447), .Y(n10340) );
  NOR2X1 U27985 ( .A(n36959), .B(n37278), .Y(n39447) );
  NOR2X1 U27986 ( .A(net171319), .B(net171113), .Y(n39745) );
  NOR2X1 U27987 ( .A(net171114), .B(net151253), .Y(n39746) );
  AND2X2 U27988 ( .A(net213207), .B(net213206), .Y(n40750) );
  AND2X2 U27989 ( .A(net215125), .B(net215124), .Y(n40953) );
  AND2X2 U27990 ( .A(net215098), .B(net215097), .Y(n40592) );
  NOR2X1 U27991 ( .A(n37136), .B(n37493), .Y(n40679) );
  CLKBUFX3 U27992 ( .A(n12238), .Y(n40391) );
  CLKBUFX3 U27993 ( .A(n11001), .Y(n40400) );
  CLKBUFX3 U27994 ( .A(n11028), .Y(n40399) );
  OR4X1 U27995 ( .A(net151458), .B(net171462), .C(net171461), .D(net151473),
        .Y(n39517) );
  NAND4X1 U27996 ( .A(n45939), .B(n45938), .C(n45937), .D(n45936), .Y(n11050)
         );
  NOR2X1 U27997 ( .A(n22918), .B(n22917), .Y(n45937) );
  NAND3BX1 U27998 ( .AN(n45951), .B(n37355), .C(n45950), .Y(n11046) );
  NOR2X1 U27999 ( .A(n10526), .B(n22887), .Y(n45950) );
  NAND4X1 U28000 ( .A(n45949), .B(n45948), .C(n45947), .D(n45946), .Y(n11041)
         );
  NAND2BX2 U28001 ( .AN(n_cell_301249_net267183), .B(net213562), .Y(n10976) );
  NAND2X1 U28002 ( .A(n41134), .B(net213565), .Y(n_cell_301249_net267183) );
  NOR2X1 U28003 ( .A(n37093), .B(n37508), .Y(n41134) );
  NAND4X1 U28004 ( .A(n46029), .B(n46028), .C(n46027), .D(n46026), .Y(n11016)
         );
  NAND4X1 U28005 ( .A(n46024), .B(n46023), .C(n46022), .D(n46021), .Y(n11217)
         );
  CLKBUFX3 U28006 ( .A(n11218), .Y(n40395) );
  NAND2BX1 U28007 ( .AN(n40774), .B(net212846), .Y(n10991) );
  NAND2X1 U28008 ( .A(n41141), .B(net212849), .Y(n40774) );
  NOR2X1 U28009 ( .A(n37037), .B(n37432), .Y(n41141) );
  CLKINVX1 U28010 ( .A(net210392), .Y(net210473) );
  NOR2X1 U28011 ( .A(n39482), .B(n_cell_301249_net269836), .Y(n40821) );
  NAND2X1 U28012 ( .A(net260830), .B(net211602), .Y(n40823) );
  NAND2X1 U28013 ( .A(n41176), .B(n10927), .Y(n41177) );
  NOR2X1 U28014 ( .A(net171392), .B(n_cell_301249_net269839), .Y(n41176) );
  CLKINVX1 U28015 ( .A(net211590), .Y(net171394) );
  CLKINVX1 U28016 ( .A(n10928), .Y(n_cell_301249_net269839) );
  NOR2X1 U28017 ( .A(n_cell_301249_net269745), .B(n_cell_301249_net269746),
        .Y(n41110) );
  NAND2X1 U28018 ( .A(n12826), .B(n12824), .Y(n41109) );
  NOR2X2 U28019 ( .A(n40846), .B(n40849), .Y(n40848) );
  NOR2X1 U28020 ( .A(n_cell_301249_net269749), .B(n_cell_303546_net277822),
        .Y(n40851) );
  CLKINVX1 U28021 ( .A(n9992), .Y(n_cell_301249_net269749) );
  NAND2X1 U28022 ( .A(n12821), .B(n13026), .Y(n40853) );
  NAND2X1 U28023 ( .A(net259677), .B(net272625), .Y(n41047) );
  NOR2X1 U28024 ( .A(net151380), .B(n_cell_301249_net269650), .Y(n41048) );
  AOI21X1 U28025 ( .A0(n40871), .A1(n40872), .B0(n40873), .Y(n40870) );
  NOR2BX1 U28026 ( .AN(net272620), .B(net171270), .Y(n40875) );
  NAND2X1 U28027 ( .A(n11558), .B(n11874), .Y(n40877) );
  CLKINVX1 U28028 ( .A(n10064), .Y(n_cell_301249_net269653) );
  NOR2X1 U28029 ( .A(net151788), .B(net151786), .Y(n40906) );
  NAND2X1 U28030 ( .A(n11885), .B(n11886), .Y(n40908) );
  CLKINVX1 U28031 ( .A(n39642), .Y(net234762) );
  CLKINVX1 U28032 ( .A(net211102), .Y(net210523) );
  AOI21X1 U28033 ( .A0(n40482), .A1(n40483), .B0(n40484), .Y(n40481) );
  OAI2BB1X1 U28034 ( .A0N(n40749), .A1N(n11894), .B0(net213230), .Y(n40484) );
  NOR2X1 U28035 ( .A(n40748), .B(n40582), .Y(n40482) );
  NAND2X1 U28036 ( .A(n40747), .B(n40762), .Y(n40483) );
  NOR2X1 U28037 ( .A(n37154), .B(n37476), .Y(n40720) );
  CLKINVX1 U28038 ( .A(n11556), .Y(n_cell_303546_net277957) );
  NOR2X1 U28039 ( .A(n37488), .B(n37147), .Y(n41057) );
  NOR2X1 U28040 ( .A(n37479), .B(n37174), .Y(n41113) );
  NAND3X1 U28041 ( .A(n40716), .B(n10630), .C(n12824), .Y(n40536) );
  NAND2BX1 U28042 ( .AN(n_cell_301249_net269874), .B(n12826), .Y(n40716) );
  NAND2X1 U28043 ( .A(n12821), .B(n9992), .Y(n40717) );
  NOR2X1 U28044 ( .A(n37478), .B(n37173), .Y(n41114) );
  NAND2X1 U28045 ( .A(n40590), .B(net211565), .Y(n40460) );
  NAND3X1 U28046 ( .A(n10619), .B(net266151), .C(n10612), .Y(net209395) );
  AOI21X1 U28047 ( .A0(n_cell_303546_net277761), .A1(n10771), .B0(n40678), .Y(
        n40559) );
  NAND2X1 U28048 ( .A(n10772), .B(n12188), .Y(n40678) );
  CLKINVX1 U28049 ( .A(n10923), .Y(n_cell_303546_net277761) );
  NAND2X1 U28050 ( .A(n40680), .B(net261069), .Y(n40561) );
  NOR2X1 U28051 ( .A(net151767), .B(n40584), .Y(n40680) );
  NOR2X1 U28052 ( .A(n_cell_303546_net277645), .B(n12190), .Y(n40584) );
  CLKINVX1 U28053 ( .A(n12188), .Y(n_cell_303546_net277645) );
  AOI21X1 U28054 ( .A0(n39611), .A1(n39612), .B0(n10463), .Y(n39610) );
  NOR3X1 U28055 ( .A(n39832), .B(n_cell_303546_net277936), .C(n39833), .Y(
        n39612) );
  OAI21XL U28056 ( .A0(n39607), .A1(n10142), .B0(n40022), .Y(n39611) );
  NAND2X1 U28057 ( .A(n10471), .B(n12168), .Y(n39832) );
  CLKINVX1 U28058 ( .A(n10456), .Y(n40021) );
  NAND3X1 U28059 ( .A(net260295), .B(net260299), .C(n39834), .Y(n39836) );
  NOR2X1 U28060 ( .A(n39835), .B(n_cell_301249_net269596), .Y(n39834) );
  NAND2X1 U28061 ( .A(n39838), .B(net260925), .Y(n39837) );
  CLKINVX1 U28062 ( .A(n11904), .Y(n39838) );
  OAI21XL U28063 ( .A0(n39759), .A1(n39762), .B0(n39867), .Y(n39769) );
  NOR2BX1 U28064 ( .AN(n10433), .B(n39865), .Y(n39867) );
  AOI21X1 U28065 ( .A0(n39760), .A1(net168846), .B0(n39761), .Y(n39759) );
  NAND2X1 U28066 ( .A(n11870), .B(n39866), .Y(n39865) );
  CLKINVX1 U28067 ( .A(n10301), .Y(n39768) );
  NAND2X1 U28068 ( .A(net259677), .B(net272625), .Y(n39869) );
  NAND2X1 U28069 ( .A(n10436), .B(n10434), .Y(n39868) );
  NOR2X1 U28070 ( .A(net171414), .B(net151584), .Y(n39995) );
  OAI21XL U28071 ( .A0(n37512), .A1(n39537), .B0(n39994), .Y(n39539) );
  NOR2X1 U28072 ( .A(net171416), .B(n10215), .Y(n39994) );
  AOI21X1 U28073 ( .A0(n39534), .A1(n39535), .B0(n39536), .Y(n39533) );
  NAND2X1 U28074 ( .A(n10635), .B(n39341), .Y(n39930) );
  OAI21XL U28075 ( .A0(n39686), .A1(n39924), .B0(n39926), .Y(n39692) );
  NAND3X1 U28076 ( .A(net210007), .B(net271515), .C(n39925), .Y(n39924) );
  NOR4X1 U28077 ( .A(n39927), .B(n39928), .C(n_cell_303546_net277636), .D(
        n39929), .Y(n39926) );
  AOI21X1 U28078 ( .A0(n39687), .A1(n39688), .B0(n37519), .Y(n39686) );
  NAND2X1 U28079 ( .A(n41118), .B(net211170), .Y(n_cell_301249_net268355) );
  CLKINVX1 U28080 ( .A(n39510), .Y(n10848) );
  NAND4BX1 U28081 ( .AN(n39408), .B(n11117), .C(n11114), .D(n11116), .Y(n10253) );
  NOR2X1 U28082 ( .A(n39490), .B(net171448), .Y(n39433) );
  CLKINVX1 U28083 ( .A(n11211), .Y(n39490) );
  NAND3X1 U28084 ( .A(n39434), .B(n11073), .C(n11072), .Y(n10240) );
  NOR2X1 U28085 ( .A(n39491), .B(net209210), .Y(n39434) );
  NAND4X1 U28086 ( .A(n11699), .B(n11705), .C(n11700), .D(n11706), .Y(n10102)
         );
  NAND3X1 U28087 ( .A(n12587), .B(n11698), .C(n12501), .Y(n10101) );
  NAND3X1 U28088 ( .A(n11694), .B(n11693), .C(n11687), .Y(n10098) );
  NAND4BX1 U28089 ( .AN(n39453), .B(n11752), .C(n11848), .D(n11751), .Y(n10112) );
  CLKINVX1 U28090 ( .A(n11756), .Y(n39453) );
  CLKINVX1 U28091 ( .A(net260900), .Y(net171168) );
  NAND3X1 U28092 ( .A(n11423), .B(n11422), .C(n11418), .Y(n9913) );
  NAND3X1 U28093 ( .A(n11415), .B(n39361), .C(n11417), .Y(n9915) );
  NOR2X1 U28094 ( .A(n39480), .B(net210242), .Y(n39361) );
  CLKINVX1 U28095 ( .A(n11414), .Y(n39480) );
  CLKINVX1 U28096 ( .A(net210416), .Y(net210512) );
  NAND3X1 U28097 ( .A(n11378), .B(n11379), .C(n39354), .Y(n10032) );
  NOR2X1 U28098 ( .A(n39634), .B(n39635), .Y(n39354) );
  CLKINVX1 U28099 ( .A(n11377), .Y(n39634) );
  CLKINVX1 U28100 ( .A(n11376), .Y(n39635) );
  OR2X1 U28101 ( .A(net171537), .B(n39902), .Y(n39658) );
  OR2X1 U28102 ( .A(net151860), .B(net171538), .Y(n39902) );
  CLKINVX1 U28103 ( .A(n10247), .Y(net168852) );
  CLKINVX1 U28104 ( .A(n39511), .Y(n10837) );
  NAND3X1 U28105 ( .A(n11209), .B(n39398), .C(n12297), .Y(n10246) );
  NOR2X1 U28106 ( .A(n39492), .B(net171440), .Y(n39398) );
  CLKINVX1 U28107 ( .A(n11208), .Y(n39492) );
  CLKINVX1 U28108 ( .A(n10527), .Y(net171136) );
  CLKINVX1 U28109 ( .A(n10157), .Y(net171139) );
  CLKINVX1 U28110 ( .A(n39589), .Y(n10162) );
  CLKINVX1 U28111 ( .A(n39592), .Y(n10158) );
  NAND3X1 U28112 ( .A(n12157), .B(n12156), .C(n39290), .Y(n10155) );
  NOR2X1 U28113 ( .A(n39558), .B(n39559), .Y(n39290) );
  CLKINVX1 U28114 ( .A(n12014), .Y(n39559) );
  CLKINVX1 U28115 ( .A(n12015), .Y(n39558) );
  CLKBUFX3 U28116 ( .A(n12648), .Y(n40389) );
  CLKINVX1 U28117 ( .A(n_cell_301249_net269449), .Y(n10481) );
  NOR2X1 U28118 ( .A(n37024), .B(n37321), .Y(n_cell_301249_net267165) );
  CLKBUFX3 U28119 ( .A(n12802), .Y(net260431) );
  NAND4BX1 U28120 ( .AN(n39335), .B(n12800), .C(n11984), .D(n11985), .Y(n10509) );
  NAND4X1 U28121 ( .A(n11990), .B(n11991), .C(n11988), .D(n11989), .Y(n10512)
         );
  NAND2X1 U28122 ( .A(n12264), .B(n12260), .Y(n10819) );
  NAND2BX2 U28123 ( .AN(n39438), .B(net212981), .Y(n10820) );
  NAND2X1 U28124 ( .A(n39942), .B(net212984), .Y(n39438) );
  AND2X2 U28125 ( .A(net212983), .B(net212982), .Y(n39942) );
  NAND3X1 U28126 ( .A(n11040), .B(n11039), .C(n11035), .Y(n10821) );
  CLKBUFX3 U28127 ( .A(n12262), .Y(n40390) );
  CLKINVX1 U28128 ( .A(n10015), .Y(net151462) );
  NAND2X1 U28129 ( .A(n12904), .B(n12901), .Y(n10686) );
  NAND3X1 U28130 ( .A(n11348), .B(n11349), .C(n39351), .Y(n10020) );
  NOR2X1 U28131 ( .A(n39629), .B(n39630), .Y(n39351) );
  CLKINVX1 U28132 ( .A(n11512), .Y(n39630) );
  CLKINVX1 U28133 ( .A(n11511), .Y(n39629) );
  NAND3X1 U28134 ( .A(n11350), .B(n11351), .C(n39352), .Y(n10018) );
  NOR2X1 U28135 ( .A(n39631), .B(n36942), .Y(n39352) );
  CLKINVX1 U28136 ( .A(n39665), .Y(n10016) );
  NAND3X1 U28137 ( .A(n13022), .B(n12867), .C(n39384), .Y(n10758) );
  NOR2X1 U28138 ( .A(n39676), .B(n39677), .Y(n39384) );
  NAND2X1 U28139 ( .A(n41068), .B(net211770), .Y(n_cell_301249_net267213) );
  CLKINVX1 U28140 ( .A(n11520), .Y(net151530) );
  NAND3X1 U28141 ( .A(net211440), .B(net211439), .C(net211441), .Y(
        n_cell_301249_net268217) );
  NAND3X1 U28142 ( .A(n11637), .B(n11638), .C(n39446), .Y(n10083) );
  AND2X2 U28143 ( .A(n12461), .B(n12589), .Y(n39446) );
  NAND4X1 U28144 ( .A(n11645), .B(n11646), .C(n11639), .D(n11640), .Y(n10082)
         );
  CLKBUFX3 U28145 ( .A(n10079), .Y(n40404) );
  CLKINVX1 U28146 ( .A(n39750), .Y(n10077) );
  CLKINVX1 U28147 ( .A(net260367), .Y(net151279) );
  NAND3X1 U28148 ( .A(net215182), .B(net215183), .C(n_cell_301249_net268242),
        .Y(n11550) );
  NOR2X1 U28149 ( .A(n36963), .B(n37289), .Y(n_cell_301249_net268242) );
  NAND4BBX1 U28150 ( .AN(n37397), .BN(n37005), .C(net214754), .D(net214752),
        .Y(n11558) );
  NAND4BBX1 U28151 ( .AN(n37396), .BN(n37004), .C(net215104), .D(net215102),
        .Y(n11874) );
  NAND4BBX1 U28152 ( .AN(n37395), .BN(n37112), .C(net214750), .D(net214748),
        .Y(n11555) );
  NAND4BBX1 U28153 ( .AN(n37398), .BN(n37113), .C(net215131), .D(net215129),
        .Y(n11556) );
  CLKINVX1 U28154 ( .A(net261020), .Y(net171327) );
  CLKBUFX3 U28155 ( .A(net209701), .Y(net260925) );
  CLKBUFX3 U28156 ( .A(net213602), .Y(net272583) );
  NAND2X1 U28157 ( .A(n37473), .B(net214988), .Y(n11902) );
  AND2X2 U28158 ( .A(net214990), .B(net214989), .Y(n40955) );
  NAND2BX1 U28159 ( .AN(n_cell_301249_net268002), .B(net214997), .Y(n11901) );
  NAND2X1 U28160 ( .A(n40954), .B(net215000), .Y(n_cell_301249_net268002) );
  AND2X2 U28161 ( .A(net214999), .B(net214998), .Y(n40954) );
  NAND2BX1 U28162 ( .AN(n_cell_301249_net268142), .B(net214979), .Y(n11893) );
  NAND2X1 U28163 ( .A(n41011), .B(net214982), .Y(n_cell_301249_net268142) );
  NOR2BX1 U28164 ( .AN(net214981), .B(n37359), .Y(n41011) );
  CLKINVX1 U28165 ( .A(n10959), .Y(net171416) );
  NAND3X1 U28166 ( .A(n12392), .B(n12213), .C(n37120), .Y(n10779) );
  OR2X1 U28167 ( .A(net171394), .B(n39545), .Y(n39544) );
  OR2X1 U28168 ( .A(net171392), .B(n10926), .Y(n39545) );
  NAND3X1 U28169 ( .A(n10946), .B(n10947), .C(n10942), .Y(n39541) );
  NAND3X1 U28170 ( .A(net212045), .B(net212044), .C(net212046), .Y(
        n_cell_301249_net267646) );
  NAND2BX2 U28171 ( .AN(n_cell_301249_net267658), .B(net212063), .Y(n11524) );
  NAND2X1 U28172 ( .A(n41062), .B(net212065), .Y(n_cell_301249_net267658) );
  NAND2BX1 U28173 ( .AN(n_cell_301249_net267652), .B(net212058), .Y(n11525) );
  NAND3X1 U28174 ( .A(net212060), .B(net212059), .C(net212061), .Y(
        n_cell_301249_net267652) );
  CLKINVX1 U28175 ( .A(net259841), .Y(net151440) );
  NAND2X1 U28176 ( .A(n40587), .B(net212055), .Y(n40429) );
  NAND2X1 U28177 ( .A(n12840), .B(n12838), .Y(n10641) );
  NAND3X1 U28178 ( .A(net212075), .B(net212074), .C(net212076), .Y(
        n_cell_301249_net267846) );
  NAND2X1 U28179 ( .A(n41061), .B(net212101), .Y(n_cell_301249_net267840) );
  NAND2X1 U28180 ( .A(n41104), .B(net212096), .Y(n_cell_301249_net267885) );
  NAND2BX2 U28181 ( .AN(n_cell_301249_net267891), .B(net212089), .Y(n10759) );
  NAND3X1 U28182 ( .A(net212091), .B(net212090), .C(net212092), .Y(
        n_cell_301249_net267891) );
  CLKBUFX3 U28183 ( .A(n10644), .Y(net271515) );
  OR2X1 U28184 ( .A(n37354), .B(net151809), .Y(n39694) );
  CLKINVX1 U28185 ( .A(n12824), .Y(net151806) );
  NOR2X1 U28186 ( .A(n37158), .B(n37483), .Y(n41111) );
  CLKINVX1 U28187 ( .A(n39653), .Y(n10700) );
  CLKINVX1 U28188 ( .A(n10025), .Y(net151653) );
  CLKINVX1 U28189 ( .A(n10026), .Y(net151666) );
  NAND2X1 U28190 ( .A(n41072), .B(net211965), .Y(n_cell_301249_net267075) );
  NAND3X1 U28191 ( .A(n12873), .B(net260488), .C(n39347), .Y(n10661) );
  NOR2X1 U28192 ( .A(n39624), .B(n39625), .Y(n39347) );
  CLKINVX1 U28193 ( .A(n11300), .Y(n39625) );
  CLKINVX1 U28194 ( .A(n11301), .Y(n39624) );
  CLKBUFX3 U28195 ( .A(n10669), .Y(net259841) );
  CLKINVX1 U28196 ( .A(n40405), .Y(net151435) );
  OR2X1 U28197 ( .A(n36945), .B(net238947), .Y(n39912) );
  CLKINVX1 U28198 ( .A(n_cell_301249_net269861), .Y(n10010) );
  NAND3X1 U28199 ( .A(net212121), .B(net212120), .C(net212122), .Y(
        n_cell_301249_net267490) );
  CLKINVX1 U28200 ( .A(n39683), .Y(n10004) );
  CLKINVX1 U28201 ( .A(n39685), .Y(n10005) );
  NAND2X1 U28202 ( .A(n41065), .B(net212041), .Y(n_cell_301249_net267484) );
  NAND2BX1 U28203 ( .AN(n_cell_301249_net267580), .B(net212027), .Y(n11264) );
  NAND2X1 U28204 ( .A(n41064), .B(net212030), .Y(n_cell_301249_net267580) );
  NAND3X1 U28205 ( .A(net211581), .B(net211580), .C(net211582), .Y(
        n_cell_301249_net268044) );
  NAND3X1 U28206 ( .A(n39284), .B(n11934), .C(net260412), .Y(n10143) );
  NOR2X1 U28207 ( .A(n39554), .B(n39553), .Y(n39284) );
  NAND3X1 U28208 ( .A(n12167), .B(n12166), .C(n39283), .Y(n10142) );
  NOR2X1 U28209 ( .A(n_cell_301249_net269578), .B(n39552), .Y(n39283) );
  NAND2X1 U28210 ( .A(n41006), .B(net214691), .Y(n_cell_301249_net267804) );
  NOR2BX1 U28211 ( .AN(net214690), .B(n37357), .Y(n41006) );
  CLKBUFX3 U28212 ( .A(n12169), .Y(net260295) );
  CLKBUFX3 U28213 ( .A(n12170), .Y(net260299) );
  NAND4X1 U28214 ( .A(net271996), .B(n12806), .C(n11916), .D(n11917), .Y(
        n10463) );
  CLKINVX1 U28215 ( .A(n39568), .Y(net234007) );
  CLKINVX1 U28216 ( .A(n12087), .Y(net151705) );
  CLKINVX1 U28217 ( .A(n12089), .Y(net171233) );
  NAND2BX1 U28218 ( .AN(n39330), .B(net214641), .Y(n10519) );
  NAND2X1 U28219 ( .A(n39818), .B(net214644), .Y(n39330) );
  NOR2BX1 U28220 ( .AN(net214643), .B(n37466), .Y(n39818) );
  NAND2BX2 U28221 ( .AN(n39329), .B(net214646), .Y(n10520) );
  NAND2X1 U28222 ( .A(n39817), .B(net214649), .Y(n39329) );
  CLKINVX1 U28223 ( .A(net209767), .Y(net171117) );
  NAND2X1 U28224 ( .A(n12675), .B(n12672), .Y(n10522) );
  CLKINVX1 U28225 ( .A(n39597), .Y(n10498) );
  CLKINVX1 U28226 ( .A(net259747), .Y(net171145) );
  CLKINVX1 U28227 ( .A(n10072), .Y(net168848) );
  CLKINVX1 U28228 ( .A(n10073), .Y(net168846) );
  CLKBUFX3 U28229 ( .A(n10432), .Y(net259665) );
  CLKBUFX3 U28230 ( .A(n10431), .Y(net259661) );
  NAND3X2 U28231 ( .A(n_cell_301249_net267742), .B(net216183), .C(net216180),
        .Y(n10433) );
  NOR2X1 U28232 ( .A(n36967), .B(n37272), .Y(n_cell_301249_net267742) );
  CLKINVX1 U28233 ( .A(n11869), .Y(net151299) );
  CLKINVX1 U28234 ( .A(n10089), .Y(net151264) );
  CLKINVX1 U28235 ( .A(n10090), .Y(net151266) );
  NAND2X1 U28236 ( .A(n40950), .B(net212560), .Y(n_cell_301249_net268342) );
  AND2X2 U28237 ( .A(net212559), .B(net212558), .Y(n40950) );
  NAND2BX1 U28238 ( .AN(n_cell_301249_net268029), .B(net213210), .Y(n10927) );
  NAND3X1 U28239 ( .A(net213212), .B(net213211), .C(net213213), .Y(
        n_cell_301249_net268029) );
  NAND2BX1 U28240 ( .AN(n_cell_301249_net268079), .B(net213215), .Y(n10923) );
  NAND2X1 U28241 ( .A(n41179), .B(net213218), .Y(n_cell_301249_net268079) );
  AND2X2 U28242 ( .A(net213217), .B(net213216), .Y(n41179) );
  NAND2BX2 U28243 ( .AN(n40452), .B(net213231), .Y(n12188) );
  NAND3X1 U28244 ( .A(net213233), .B(net213232), .C(net213234), .Y(n40452) );
  NAND2BX1 U28245 ( .AN(n40455), .B(net213236), .Y(n12190) );
  NAND2X1 U28246 ( .A(n40679), .B(net213239), .Y(n40455) );
  NAND2BX2 U28247 ( .AN(n39386), .B(net212861), .Y(n10808) );
  NAND2X1 U28248 ( .A(n39939), .B(net212864), .Y(n39386) );
  NOR2X1 U28249 ( .A(n37035), .B(n37420), .Y(n39939) );
  NAND2X1 U28250 ( .A(n39940), .B(net212869), .Y(n39387) );
  NOR2X1 U28251 ( .A(n37029), .B(n37419), .Y(n39940) );
  NAND2X1 U28252 ( .A(n39941), .B(net212874), .Y(n39388) );
  NOR2X1 U28253 ( .A(n37171), .B(n37418), .Y(n39941) );
  CLKINVX1 U28254 ( .A(n40391), .Y(net151509) );
  NAND4BX1 U28255 ( .AN(n39440), .B(n11002), .C(n10996), .D(n10997), .Y(n10902) );
  CLKINVX1 U28256 ( .A(n40400), .Y(n39440) );
  CLKINVX1 U28257 ( .A(n11131), .Y(net171430) );
  CLKINVX1 U28258 ( .A(n39505), .Y(n10875) );
  CLKINVX1 U28259 ( .A(n47805), .Y(n46305) );
  NAND2BX2 U28260 ( .AN(n39395), .B(net213016), .Y(n10233) );
  NAND2X1 U28261 ( .A(n39976), .B(net213017), .Y(n39395) );
  NOR2X1 U28262 ( .A(n37056), .B(n37436), .Y(n39976) );
  NOR2X1 U28263 ( .A(n39488), .B(n39489), .Y(n39397) );
  CLKINVX1 U28264 ( .A(n11058), .Y(n39489) );
  CLKINVX1 U28265 ( .A(n39517), .Y(n10237) );
  NAND2BX2 U28266 ( .AN(n39396), .B(net213022), .Y(n10232) );
  NAND2X1 U28267 ( .A(n39975), .B(net213023), .Y(n39396) );
  NOR2X1 U28268 ( .A(n37055), .B(n37407), .Y(n39975) );
  NAND3X1 U28269 ( .A(n11050), .B(n12270), .C(n39437), .Y(n10230) );
  NOR2X1 U28270 ( .A(n39520), .B(n39521), .Y(n39437) );
  CLKINVX1 U28271 ( .A(n12389), .Y(n39521) );
  NAND2X1 U28272 ( .A(n11041), .B(n11046), .Y(n10231) );
  NAND3X1 U28273 ( .A(n10973), .B(n_cell_303546_net275998), .C(n39385), .Y(
        n10219) );
  NOR2X1 U28274 ( .A(n39483), .B(n39484), .Y(n39385) );
  CLKINVX1 U28275 ( .A(n10976), .Y(n39484) );
  CLKINVX1 U28276 ( .A(n10218), .Y(net151557) );
  CLKINVX1 U28277 ( .A(net259873), .Y(net151541) );
  NAND2BX2 U28278 ( .AN(n40796), .B(net213447), .Y(n10959) );
  NAND2X1 U28279 ( .A(n41131), .B(net213450), .Y(n40796) );
  NOR2X1 U28280 ( .A(n37132), .B(n37503), .Y(n41131) );
  NAND3X1 U28281 ( .A(n10958), .B(n10957), .C(n10960), .Y(n10215) );
  NAND2X1 U28282 ( .A(n39983), .B(net212904), .Y(n39390) );
  NOR2X1 U28283 ( .A(n37091), .B(n37416), .Y(n39983) );
  NAND2X1 U28284 ( .A(n39984), .B(net212909), .Y(n39389) );
  NOR2X1 U28285 ( .A(n37030), .B(n37415), .Y(n39984) );
  NOR2X1 U28286 ( .A(n37364), .B(n39982), .Y(n39391) );
  NAND2X1 U28287 ( .A(net212913), .B(net212912), .Y(n39982) );
  NAND3X2 U28288 ( .A(n39392), .B(net212899), .C(net212896), .Y(n10810) );
  NOR2X1 U28289 ( .A(n37034), .B(n37414), .Y(n39392) );
  NAND3X1 U28290 ( .A(n11017), .B(n11018), .C(n39439), .Y(n10227) );
  NOR2X1 U28291 ( .A(n39487), .B(net171472), .Y(n39439) );
  NAND3X1 U28292 ( .A(n11217), .B(n11016), .C(n39393), .Y(n10228) );
  NOR2X1 U28293 ( .A(n39485), .B(n39486), .Y(n39393) );
  CLKINVX1 U28294 ( .A(n40395), .Y(n39486) );
  NAND4X1 U28295 ( .A(n11007), .B(n12246), .C(n12391), .D(n11006), .Y(n10223)
         );
  NAND2X1 U28296 ( .A(n41138), .B(net212834), .Y(n_cell_301249_net266944) );
  NOR2X1 U28297 ( .A(n37038), .B(n37430), .Y(n41138) );
  NAND2X1 U28298 ( .A(n41139), .B(net212829), .Y(n40779) );
  NAND3X1 U28299 ( .A(n10990), .B(n10992), .C(n10991), .Y(n10798) );
  NAND2BX2 U28300 ( .AN(n_cell_301249_net266950), .B(net212836), .Y(n10903) );
  NAND2X1 U28301 ( .A(n41145), .B(net212839), .Y(n_cell_301249_net266950) );
  NOR2X1 U28302 ( .A(n37040), .B(n37428), .Y(n41145) );
  CLKBUFX3 U28303 ( .A(n42457), .Y(n42455) );
  CLKBUFX3 U28304 ( .A(n42481), .Y(n42477) );
  AOI21X1 U28305 ( .A0(n41181), .A1(n10926), .B0(n41182), .Y(n40826) );
  NAND2X1 U28306 ( .A(n10923), .B(n10776), .Y(n41182) );
  NOR2X1 U28307 ( .A(n_cell_301249_net269839), .B(n_cell_303546_net277759),
        .Y(n41181) );
  NAND4X1 U28308 ( .A(n10771), .B(net261069), .C(net209087), .D(n10772), .Y(
        n40827) );
  NAND2X1 U28309 ( .A(n12186), .B(net260302), .Y(n41184) );
  NOR2X1 U28310 ( .A(net171437), .B(net171439), .Y(n41183) );
  NAND2X1 U28311 ( .A(n41123), .B(net213315), .Y(n_cell_301249_net268380) );
  NOR2X1 U28312 ( .A(n37140), .B(n37496), .Y(n41123) );
  NOR2X1 U28313 ( .A(n39934), .B(n_cell_301249_net269758), .Y(n40855) );
  NAND2X1 U28314 ( .A(net209974), .B(net209976), .Y(n40857) );
  CLKINVX1 U28315 ( .A(n10612), .Y(n_cell_301249_net269764) );
  NAND3X1 U28316 ( .A(net211189), .B(net211188), .C(net211190), .Y(
        n_cell_301249_net268398) );
  NOR2X1 U28317 ( .A(n_cell_301249_net269653), .B(n39698), .Y(n41050) );
  NAND2X1 U28318 ( .A(n11556), .B(n11555), .Y(n41049) );
  NOR2BX1 U28319 ( .AN(net260346), .B(n39699), .Y(n40879) );
  NAND2X1 U28320 ( .A(n11549), .B(n11550), .Y(n40881) );
  NAND2X1 U28321 ( .A(net260394), .B(net260449), .Y(n40912) );
  NOR2X1 U28322 ( .A(net151773), .B(net151775), .Y(n40910) );
  CLKINVX1 U28323 ( .A(n_cell_301249_net269477), .Y(n10437) );
  CLKINVX1 U28324 ( .A(n11537), .Y(n39549) );
  CLKBUFX3 U28325 ( .A(net217954), .Y(n40270) );
  CLKBUFX3 U28326 ( .A(net221900), .Y(net266201) );
  CLKBUFX3 U28327 ( .A(net221978), .Y(net221900) );
  CLKBUFX3 U28328 ( .A(net217952), .Y(n40271) );
  CLKBUFX3 U28329 ( .A(n10446), .Y(net271431) );
  CLKINVX1 U28330 ( .A(n11886), .Y(n40488) );
  NOR2X1 U28331 ( .A(n40481), .B(net171274), .Y(n40485) );
  CLKINVX1 U28332 ( .A(n11883), .Y(n40760) );
  NAND2X1 U28333 ( .A(n37474), .B(net215132), .Y(n11884) );
  CLKINVX1 U28334 ( .A(net209395), .Y(n40759) );
  CLKINVX1 U28335 ( .A(n12395), .Y(n40491) );
  NAND3X1 U28336 ( .A(net214739), .B(net214740), .C(n_cell_301249_net268236),
        .Y(n11549) );
  NOR2X1 U28337 ( .A(n37046), .B(n37288), .Y(n_cell_301249_net268236) );
  NAND4BX1 U28338 ( .AN(n37393), .B(net215158), .C(net215155), .D(net215156),
        .Y(n11543) );
  NAND4BBX1 U28339 ( .AN(n37111), .BN(n37399), .C(net214746), .D(net214744),
        .Y(n11544) );
  NAND3X1 U28340 ( .A(net215194), .B(n40799), .C(net215192), .Y(n11541) );
  NOR2X1 U28341 ( .A(n37156), .B(n37380), .Y(n40799) );
  NAND2BX1 U28342 ( .AN(n9747), .B(n40599), .Y(n40567) );
  NOR3BXL U28343 ( .AN(net171380), .B(net260384), .C(net219434), .Y(n40599) );
  NAND3X1 U28344 ( .A(net211445), .B(net211444), .C(net211446), .Y(
        n_cell_301249_net268223) );
  OAI21XL U28345 ( .A0(n40535), .A1(n37518), .B0(n40718), .Y(n40538) );
  AOI21X1 U28346 ( .A0(n_cell_303546_net277822), .A1(n12821), .B0(n39619), .Y(
        n40718) );
  NOR2X1 U28347 ( .A(n40531), .B(n40536), .Y(n40535) );
  NAND2BX1 U28348 ( .AN(n_cell_301249_net268091), .B(net211458), .Y(n11241) );
  NAND2X1 U28349 ( .A(n41114), .B(net211461), .Y(n_cell_301249_net268091) );
  NOR2X1 U28350 ( .A(n12594), .B(n40491), .Y(n40635) );
  NAND2X1 U28351 ( .A(n12395), .B(n12594), .Y(n_cell_301249_net269475) );
  CLKINVX1 U28352 ( .A(net260394), .Y(n39773) );
  OAI21XL U28353 ( .A0(n10136), .A1(n39613), .B0(n40387), .Y(n39617) );
  AOI21X1 U28354 ( .A0(n39614), .A1(n39615), .B0(n10137), .Y(n39613) );
  NOR2BX1 U28355 ( .AN(net272583), .B(n39837), .Y(n39615) );
  OAI21XL U28356 ( .A0(n39836), .A1(n39610), .B0(n40021), .Y(n39614) );
  NAND4X1 U28357 ( .A(net271431), .B(n10447), .C(n10448), .D(n12596), .Y(
        n39618) );
  NAND2BX2 U28358 ( .AN(n9747), .B(n_cell_301249_net269478), .Y(
        n_cell_301249_net269477) );
  CLKINVX1 U28359 ( .A(net264532), .Y(n_cell_301249_net269478) );
  OAI21XL U28360 ( .A0(n39767), .A1(n37529), .B0(n39870), .Y(n39772) );
  NOR2X1 U28361 ( .A(n39869), .B(n39868), .Y(n39870) );
  AOI21X1 U28362 ( .A0(n39768), .A1(n39769), .B0(n39764), .Y(n39767) );
  NOR2BX1 U28363 ( .AN(net272620), .B(n39872), .Y(n39771) );
  NAND2X1 U28364 ( .A(n39871), .B(n12408), .Y(n39872) );
  NOR2BX1 U28365 ( .AN(net214756), .B(n_cell_301249_net269650), .Y(n39871) );
  CLKINVX1 U28366 ( .A(n10062), .Y(net168849) );
  CLKINVX1 U28367 ( .A(net260302), .Y(net151772) );
  CLKINVX1 U28368 ( .A(n10775), .Y(n39997) );
  NAND2X1 U28369 ( .A(n10771), .B(n10772), .Y(n39999) );
  AOI21X1 U28370 ( .A0(n37346), .A1(n39547), .B0(n39544), .Y(n39546) );
  OAI21XL U28371 ( .A0(n39538), .A1(n39541), .B0(n37123), .Y(n39547) );
  AOI21X1 U28372 ( .A0(n39539), .A1(n39540), .B0(n10779), .Y(n39538) );
  NOR3BXL U28373 ( .AN(n39995), .B(net151586), .C(net171412), .Y(n39540) );
  CLKINVX1 U28374 ( .A(n12811), .Y(net151766) );
  CLKINVX1 U28375 ( .A(n12813), .Y(net151769) );
  CLKINVX1 U28376 ( .A(n9988), .Y(n39932) );
  NOR2X1 U28377 ( .A(n39690), .B(n39694), .Y(n39695) );
  AOI21X1 U28378 ( .A0(n39691), .A1(n39692), .B0(n39693), .Y(n39690) );
  OR2X1 U28379 ( .A(n_cell_301249_net269872), .B(n39930), .Y(n39693) );
  NOR2X1 U28380 ( .A(n_cell_303546_net277804), .B(n39689), .Y(n39691) );
  CLKINVX1 U28381 ( .A(n10621), .Y(n40027) );
  NAND2BX1 U28382 ( .AN(n_cell_301249_net268392), .B(net211558), .Y(n10619) );
  NAND3X1 U28383 ( .A(net211560), .B(net211559), .C(net211561), .Y(
        n_cell_301249_net268392) );
  CLKINVX1 U28384 ( .A(n40403), .Y(net151404) );
  CLKINVX1 U28385 ( .A(n40401), .Y(net168842) );
  CLKINVX1 U28386 ( .A(n40402), .Y(net168843) );
  CLKINVX1 U28387 ( .A(n39670), .Y(n10677) );
  CLKINVX1 U28388 ( .A(n39666), .Y(n10683) );
  NAND2X1 U28389 ( .A(n39442), .B(net260346), .Y(n10067) );
  NOR2X1 U28390 ( .A(n39698), .B(n39699), .Y(n39442) );
  CLKINVX1 U28391 ( .A(n39764), .Y(n10293) );
  NAND4X1 U28392 ( .A(n11874), .B(n11558), .C(n11555), .D(n11556), .Y(n10066)
         );
  NAND4X2 U28393 ( .A(net215119), .B(net215121), .C(net215122), .D(net215120),
        .Y(n10064) );
  NAND3X1 U28394 ( .A(n39441), .B(n11542), .C(n11541), .Y(n10063) );
  NOR2X1 U28395 ( .A(n39548), .B(n39549), .Y(n39441) );
  CLKINVX1 U28396 ( .A(net212088), .Y(net171412) );
  NOR2X1 U28397 ( .A(net171386), .B(net171388), .Y(n39543) );
  CLKINVX1 U28398 ( .A(net209101), .Y(net171386) );
  CLKINVX1 U28399 ( .A(net272417), .Y(net171388) );
  CLKINVX1 U28400 ( .A(n39544), .Y(n10199) );
  NOR2X1 U28401 ( .A(n39481), .B(n39482), .Y(n39542) );
  CLKINVX1 U28402 ( .A(n39541), .Y(n10204) );
  NAND3X1 U28403 ( .A(n10630), .B(n10631), .C(n10629), .Y(n9988) );
  NAND3X1 U28404 ( .A(n11524), .B(n11525), .C(n11263), .Y(n9999) );
  CLKINVX1 U28405 ( .A(n39689), .Y(n10639) );
  CLKINVX1 U28406 ( .A(n39694), .Y(n9993) );
  NAND2BX2 U28407 ( .AN(n_cell_301249_net268109), .B(net211574), .Y(n9992) );
  NAND2X1 U28408 ( .A(n41111), .B(net211576), .Y(n_cell_301249_net268109) );
  NAND4BX1 U28409 ( .AN(n39343), .B(n11264), .C(n12848), .D(n13025), .Y(n9900)
         );
  CLKINVX1 U28410 ( .A(net271431), .Y(net171262) );
  CLKINVX1 U28411 ( .A(n12596), .Y(net151775) );
  CLKBUFX3 U28412 ( .A(n12808), .Y(net260449) );
  CLKINVX1 U28413 ( .A(n_cell_301249_net269475), .Y(n10438) );
  CLKBUFX3 U28414 ( .A(n12597), .Y(net260394) );
  CLKBUFX3 U28415 ( .A(n9946), .Y(n40387) );
  CLKINVX1 U28416 ( .A(n10136), .Y(net151819) );
  CLKINVX1 U28417 ( .A(n10137), .Y(net151812) );
  CLKINVX1 U28418 ( .A(n12168), .Y(net171178) );
  CLKINVX1 U28419 ( .A(n10130), .Y(net151779) );
  CLKINVX1 U28420 ( .A(net272620), .Y(net171294) );
  CLKINVX1 U28421 ( .A(n39762), .Y(n10306) );
  NAND3X1 U28422 ( .A(n10923), .B(n10927), .C(n10928), .Y(n10775) );
  NAND2BX2 U28423 ( .AN(n_cell_301249_net268160), .B(net213200), .Y(n10771) );
  NAND3X1 U28424 ( .A(net213202), .B(net213201), .C(net213203), .Y(
        n_cell_301249_net268160) );
  NAND2BX2 U28425 ( .AN(n_cell_301249_net268154), .B(net213195), .Y(n10772) );
  NAND3X1 U28426 ( .A(net213197), .B(net213196), .C(net213198), .Y(
        n_cell_301249_net268154) );
  NAND2BX2 U28427 ( .AN(n_cell_301249_net268085), .B(net213190), .Y(n10776) );
  NAND2X1 U28428 ( .A(n41180), .B(net213193), .Y(n_cell_301249_net268085) );
  AND2X2 U28429 ( .A(net213192), .B(net213191), .Y(n41180) );
  CLKINVX1 U28430 ( .A(n39525), .Y(n10815) );
  NAND2BX2 U28431 ( .AN(n40801), .B(net213661), .Y(n9716) );
  NAND2X1 U28432 ( .A(net213660), .B(net213659), .Y(n40801) );
  CLKBUFX3 U28433 ( .A(net221978), .Y(net221902) );
  CLKBUFX3 U28434 ( .A(net221978), .Y(net221904) );
  CLKINVX1 U28435 ( .A(n42651), .Y(n41285) );
  OAI21X2 U28436 ( .A0(n40824), .A1(n37527), .B0(n41185), .Y(n41192) );
  NOR2X1 U28437 ( .A(n_cell_301249_net269853), .B(n40001), .Y(n41185) );
  NOR2X1 U28438 ( .A(net209402), .B(n41186), .Y(n41187) );
  NAND2X1 U28439 ( .A(n10762), .B(n10763), .Y(n41186) );
  NAND2X1 U28440 ( .A(n12811), .B(n12813), .Y(n41117) );
  NOR2X1 U28441 ( .A(n_cell_301249_net269763), .B(n_cell_301249_net269764),
        .Y(n41120) );
  NOR2X1 U28442 ( .A(net218294), .B(n41121), .Y(n41122) );
  NAND2X1 U28443 ( .A(n10619), .B(n10614), .Y(n41121) );
  NOR2X1 U28444 ( .A(net266549), .B(n41198), .Y(n40913) );
  NAND2X1 U28445 ( .A(n11543), .B(n11544), .Y(n41051) );
  NOR2BX1 U28446 ( .AN(n11541), .B(n_cell_303546_net277506), .Y(n41052) );
  OAI2BB2XL U28447 ( .B0(n40909), .B1(n41018), .A0N(n41056), .A1N(n10437), .Y(
        n41188) );
  NOR2X1 U28448 ( .A(n9716), .B(n36894), .Y(n41056) );
  NAND2X1 U28449 ( .A(n10438), .B(n10437), .Y(n41018) );
  AOI21X1 U28450 ( .A0(n40910), .A1(n40911), .B0(n40912), .Y(n40909) );
  NOR2X1 U28451 ( .A(n41055), .B(n_cell_301249_net269477), .Y(n41054) );
  NAND2X1 U28452 ( .A(n41053), .B(n36928), .Y(n41055) );
  NOR2X1 U28453 ( .A(n39548), .B(n39549), .Y(n41053) );
  CLKBUFX3 U28454 ( .A(net217964), .Y(n40267) );
  CLKINVX1 U28455 ( .A(net266201), .Y(net221822) );
  CLKINVX1 U28456 ( .A(net266201), .Y(net221808) );
  CLKINVX1 U28457 ( .A(net266218), .Y(net221846) );
  CLKINVX1 U28458 ( .A(net266201), .Y(net221824) );
  CLKINVX1 U28459 ( .A(net266201), .Y(net221826) );
  CLKINVX1 U28460 ( .A(net266201), .Y(net221818) );
  CLKINVX1 U28461 ( .A(n40316), .Y(net217010) );
  CLKINVX1 U28462 ( .A(net266201), .Y(net221814) );
  CLKINVX1 U28463 ( .A(net266201), .Y(net221816) );
  CLKINVX1 U28464 ( .A(n40317), .Y(net216980) );
  CLKINVX1 U28465 ( .A(n40317), .Y(net216994) );
  CLKINVX1 U28466 ( .A(n40317), .Y(net216996) );
  CLKBUFX3 U28467 ( .A(net217070), .Y(n40335) );
  CLKINVX1 U28468 ( .A(n40314), .Y(net217070) );
  CLKBUFX3 U28469 ( .A(net217974), .Y(n40264) );
  CLKINVX1 U28470 ( .A(n40183), .Y(net217974) );
  CLKBUFX3 U28471 ( .A(net221754), .Y(net264827) );
  CLKINVX1 U28472 ( .A(net221954), .Y(net221754) );
  CLKINVX1 U28473 ( .A(net218202), .Y(net217934) );
  CLKBUFX3 U28474 ( .A(net217092), .Y(n40325) );
  CLKINVX1 U28475 ( .A(n40313), .Y(net217094) );
  CLKINVX1 U28476 ( .A(net266201), .Y(net221828) );
  CLKINVX1 U28477 ( .A(net218150), .Y(net218050) );
  CLKBUFX3 U28478 ( .A(net217072), .Y(n40334) );
  CLKINVX1 U28479 ( .A(n40314), .Y(net217072) );
  CLKINVX1 U28480 ( .A(net218150), .Y(net218036) );
  CLKINVX1 U28481 ( .A(net266201), .Y(net221820) );
  CLKBUFX3 U28482 ( .A(net217056), .Y(n40342) );
  CLKBUFX3 U28483 ( .A(net217050), .Y(n40345) );
  CLKBUFX3 U28484 ( .A(net217988), .Y(n40257) );
  CLKBUFX3 U28485 ( .A(net217068), .Y(n40336) );
  CLKINVX1 U28486 ( .A(n40314), .Y(net217068) );
  CLKBUFX3 U28487 ( .A(net217978), .Y(n40262) );
  CLKINVX1 U28488 ( .A(n40183), .Y(net217978) );
  CLKBUFX3 U28489 ( .A(net217976), .Y(n40263) );
  CLKINVX1 U28490 ( .A(n40183), .Y(net217976) );
  CLKBUFX3 U28491 ( .A(net217052), .Y(n40344) );
  CLKBUFX3 U28492 ( .A(net221758), .Y(net264865) );
  CLKINVX1 U28493 ( .A(net221954), .Y(net221758) );
  CLKBUFX3 U28494 ( .A(net217060), .Y(n40340) );
  CLKBUFX3 U28495 ( .A(net217980), .Y(n40261) );
  CLKINVX1 U28496 ( .A(net218146), .Y(net217980) );
  CLKBUFX3 U28497 ( .A(net217084), .Y(n40328) );
  CLKINVX1 U28498 ( .A(n40314), .Y(net217084) );
  CLKINVX1 U28499 ( .A(net218150), .Y(net218048) );
  CLKINVX1 U28500 ( .A(n40313), .Y(net217100) );
  CLKINVX1 U28501 ( .A(n40317), .Y(net216992) );
  CLKBUFX3 U28502 ( .A(net217102), .Y(n40320) );
  CLKBUFX3 U28503 ( .A(net217094), .Y(n40324) );
  CLKBUFX3 U28504 ( .A(net218026), .Y(n40238) );
  CLKINVX1 U28505 ( .A(net218148), .Y(net218026) );
  CLKBUFX3 U28506 ( .A(net217064), .Y(n40338) );
  CLKINVX1 U28507 ( .A(n40314), .Y(net217064) );
  CLKBUFX3 U28508 ( .A(net218138), .Y(n40184) );
  CLKINVX1 U28509 ( .A(n40182), .Y(net218138) );
  CLKBUFX3 U28510 ( .A(net217100), .Y(n40321) );
  CLKBUFX3 U28511 ( .A(net218024), .Y(n40239) );
  CLKINVX1 U28512 ( .A(net218148), .Y(net218024) );
  CLKBUFX3 U28513 ( .A(net217984), .Y(n40259) );
  CLKINVX1 U28514 ( .A(net218146), .Y(net217984) );
  CLKINVX1 U28515 ( .A(net266218), .Y(net221832) );
  CLKBUFX3 U28516 ( .A(net217972), .Y(n40265) );
  CLKINVX1 U28517 ( .A(n40183), .Y(net217972) );
  CLKBUFX3 U28518 ( .A(net221752), .Y(net264808) );
  CLKINVX1 U28519 ( .A(net221910), .Y(net221752) );
  CLKBUFX3 U28520 ( .A(net217104), .Y(n40319) );
  CLKINVX1 U28521 ( .A(n40313), .Y(net217104) );
  CLKBUFX3 U28522 ( .A(net218028), .Y(n40237) );
  CLKINVX1 U28523 ( .A(net218148), .Y(net218028) );
  CLKBUFX3 U28524 ( .A(net217970), .Y(n40266) );
  CLKINVX1 U28525 ( .A(n40183), .Y(net217970) );
  CLKINVX1 U28526 ( .A(n40315), .Y(net217050) );
  CLKINVX1 U28527 ( .A(n40315), .Y(net217052) );
  CLKINVX1 U28528 ( .A(net218232), .Y(net217946) );
  CLKBUFX3 U28529 ( .A(net218008), .Y(n40247) );
  CLKINVX1 U28530 ( .A(net218148), .Y(net218008) );
  CLKINVX1 U28531 ( .A(net218148), .Y(net218016) );
  CLKINVX1 U28532 ( .A(net218148), .Y(net218006) );
  CLKINVX1 U28533 ( .A(net218154), .Y(net217938) );
  CLKINVX1 U28534 ( .A(net218148), .Y(net218014) );
  CLKINVX1 U28535 ( .A(net218148), .Y(net218018) );
  CLKINVX1 U28536 ( .A(net218148), .Y(net218010) );
  CLKINVX1 U28537 ( .A(n40183), .Y(net217960) );
  CLKBUFX3 U28538 ( .A(net221724), .Y(net264592) );
  CLKINVX1 U28539 ( .A(net266151), .Y(net221724) );
  CLKBUFX3 U28540 ( .A(net217026), .Y(n40355) );
  CLKBUFX3 U28541 ( .A(net217030), .Y(n40353) );
  CLKBUFX3 U28542 ( .A(net221872), .Y(net265948) );
  CLKINVX1 U28543 ( .A(net266235), .Y(net221872) );
  CLKBUFX3 U28544 ( .A(net221868), .Y(net265910) );
  CLKINVX1 U28545 ( .A(net266235), .Y(net221868) );
  CLKBUFX3 U28546 ( .A(net217180), .Y(n40285) );
  CLKBUFX3 U28547 ( .A(net217028), .Y(n40354) );
  CLKINVX1 U28548 ( .A(net218156), .Y(net218112) );
  CLKBUFX3 U28549 ( .A(net221870), .Y(net265929) );
  CLKINVX1 U28550 ( .A(net266235), .Y(net221870) );
  CLKBUFX3 U28551 ( .A(net217990), .Y(n40256) );
  CLKINVX1 U28552 ( .A(net218146), .Y(net217990) );
  CLKBUFX3 U28553 ( .A(net217024), .Y(n40356) );
  CLKINVX1 U28554 ( .A(n40316), .Y(net217024) );
  CLKINVX1 U28555 ( .A(net218156), .Y(net218108) );
  CLKINVX1 U28556 ( .A(n40315), .Y(net217060) );
  CLKINVX1 U28557 ( .A(n40315), .Y(net217054) );
  CLKINVX1 U28558 ( .A(net218154), .Y(net217932) );
  CLKINVX1 U28559 ( .A(net221986), .Y(net221740) );
  CLKINVX1 U28560 ( .A(net221962), .Y(net221756) );
  CLKBUFX3 U28561 ( .A(net217186), .Y(n40282) );
  CLKINVX1 U28562 ( .A(n40315), .Y(net217046) );
  CLKINVX1 U28563 ( .A(n40317), .Y(net216984) );
  CLKBUFX3 U28564 ( .A(net217002), .Y(n40365) );
  CLKINVX1 U28565 ( .A(n40317), .Y(net217002) );
  CLKBUFX3 U28566 ( .A(net221882), .Y(net266043) );
  CLKINVX1 U28567 ( .A(net266235), .Y(net221882) );
  CLKINVX1 U28568 ( .A(n40317), .Y(net217004) );
  CLKINVX1 U28569 ( .A(net218156), .Y(net218128) );
  CLKBUFX3 U28570 ( .A(net221884), .Y(net266062) );
  CLKINVX1 U28571 ( .A(net266235), .Y(net221884) );
  CLKBUFX3 U28572 ( .A(net221806), .Y(net265321) );
  CLKBUFX3 U28573 ( .A(net218062), .Y(n40221) );
  CLKINVX1 U28574 ( .A(net218152), .Y(net218062) );
  CLKINVX1 U28575 ( .A(net221970), .Y(net221790) );
  CLKINVX1 U28576 ( .A(n40315), .Y(net217048) );
  CLKBUFX3 U28577 ( .A(net218078), .Y(n40213) );
  CLKINVX1 U28578 ( .A(net218152), .Y(net218078) );
  CLKINVX1 U28579 ( .A(net266201), .Y(net221812) );
  CLKINVX1 U28580 ( .A(n40315), .Y(net217034) );
  CLKINVX1 U28581 ( .A(net221908), .Y(net221768) );
  CLKINVX1 U28582 ( .A(n40316), .Y(net217012) );
  CLKINVX1 U28583 ( .A(net221972), .Y(net221798) );
  CLKINVX1 U28584 ( .A(n40315), .Y(net217058) );
  BUFX4 U28585 ( .A(net221796), .Y(net265226) );
  CLKINVX1 U28586 ( .A(net221942), .Y(net221796) );
  BUFX4 U28587 ( .A(net221784), .Y(net265112) );
  CLKINVX1 U28588 ( .A(net221930), .Y(net221784) );
  CLKBUFX3 U28589 ( .A(net218080), .Y(n40212) );
  CLKINVX1 U28590 ( .A(net218152), .Y(net218080) );
  CLKBUFX3 U28591 ( .A(net216962), .Y(n40385) );
  CLKINVX1 U28592 ( .A(n40287), .Y(net216962) );
  CLKBUFX3 U28593 ( .A(net218082), .Y(n40211) );
  CLKINVX1 U28594 ( .A(net218154), .Y(net218082) );
  CLKBUFX3 U28595 ( .A(net216964), .Y(n40384) );
  CLKINVX1 U28596 ( .A(n40314), .Y(net216964) );
  CLKBUFX3 U28597 ( .A(net221846), .Y(net265701) );
  CLKINVX1 U28598 ( .A(net218156), .Y(net218126) );
  CLKBUFX3 U28599 ( .A(net218084), .Y(n40210) );
  CLKINVX1 U28600 ( .A(net218154), .Y(net218084) );
  CLKBUFX3 U28601 ( .A(net221852), .Y(net265758) );
  CLKINVX1 U28602 ( .A(n40317), .Y(net216998) );
  CLKBUFX3 U28603 ( .A(net221878), .Y(net266005) );
  CLKINVX1 U28604 ( .A(net266235), .Y(net221878) );
  CLKBUFX3 U28605 ( .A(net218124), .Y(n40190) );
  CLKBUFX3 U28606 ( .A(net221880), .Y(net266024) );
  CLKBUFX3 U28607 ( .A(net216982), .Y(n40375) );
  CLKINVX1 U28608 ( .A(net218152), .Y(net218060) );
  CLKBUFX3 U28609 ( .A(net218086), .Y(n40209) );
  CLKINVX1 U28610 ( .A(net218154), .Y(net218086) );
  CLKINVX1 U28611 ( .A(net217226), .Y(net216966) );
  CLKBUFX3 U28612 ( .A(net221848), .Y(net265720) );
  CLKINVX1 U28613 ( .A(net218150), .Y(net218044) );
  CLKBUFX3 U28614 ( .A(net217080), .Y(n40330) );
  CLKINVX1 U28615 ( .A(n40314), .Y(net217080) );
  CLKBUFX3 U28616 ( .A(net217032), .Y(n40352) );
  CLKBUFX3 U28617 ( .A(net221874), .Y(net265967) );
  CLKINVX1 U28618 ( .A(net266235), .Y(net221874) );
  CLKBUFX3 U28619 ( .A(net218068), .Y(n40218) );
  CLKINVX1 U28620 ( .A(net218152), .Y(net218068) );
  CLKBUFX3 U28621 ( .A(net216988), .Y(n40372) );
  CLKINVX1 U28622 ( .A(n40317), .Y(net216988) );
  CLKBUFX3 U28623 ( .A(net218070), .Y(n40217) );
  CLKINVX1 U28624 ( .A(net218152), .Y(net218070) );
  CLKBUFX3 U28625 ( .A(net221834), .Y(net265587) );
  CLKBUFX3 U28626 ( .A(net216972), .Y(n40380) );
  CLKINVX1 U28627 ( .A(n40287), .Y(net216972) );
  CLKBUFX3 U28628 ( .A(net218092), .Y(n40206) );
  CLKINVX1 U28629 ( .A(net218154), .Y(net218092) );
  CLKBUFX3 U28630 ( .A(net218094), .Y(n40205) );
  CLKINVX1 U28631 ( .A(net218154), .Y(net218094) );
  CLKBUFX3 U28632 ( .A(net221830), .Y(net265549) );
  CLKBUFX3 U28633 ( .A(net218090), .Y(n40207) );
  CLKINVX1 U28634 ( .A(net218154), .Y(net218090) );
  CLKBUFX3 U28635 ( .A(net216990), .Y(n40371) );
  CLKINVX1 U28636 ( .A(n40317), .Y(net216990) );
  CLKBUFX3 U28637 ( .A(net221800), .Y(net265264) );
  CLKINVX1 U28638 ( .A(net218156), .Y(net218120) );
  CLKBUFX3 U28639 ( .A(net216986), .Y(n40373) );
  CLKINVX1 U28640 ( .A(n40317), .Y(net216986) );
  CLKBUFX3 U28641 ( .A(net218066), .Y(n40219) );
  CLKINVX1 U28642 ( .A(net218152), .Y(net218066) );
  CLKBUFX3 U28643 ( .A(net221832), .Y(net265568) );
  CLKBUFX3 U28644 ( .A(net216974), .Y(n40379) );
  CLKINVX1 U28645 ( .A(n40306), .Y(net216974) );
  CLKBUFX3 U28646 ( .A(net218096), .Y(n40204) );
  CLKINVX1 U28647 ( .A(net218154), .Y(net218096) );
  CLKBUFX3 U28648 ( .A(net218088), .Y(n40208) );
  CLKINVX1 U28649 ( .A(net218154), .Y(net218088) );
  CLKBUFX3 U28650 ( .A(net218072), .Y(n40216) );
  CLKINVX1 U28651 ( .A(net218152), .Y(net218072) );
  CLKBUFX3 U28652 ( .A(net221836), .Y(net265606) );
  CLKINVX1 U28653 ( .A(net266218), .Y(net221836) );
  CLKBUFX3 U28654 ( .A(net216992), .Y(n40370) );
  CLKBUFX3 U28655 ( .A(net218074), .Y(n40215) );
  BUFX4 U28656 ( .A(net221838), .Y(net265625) );
  CLKINVX1 U28657 ( .A(net266218), .Y(net221838) );
  CLKBUFX3 U28658 ( .A(net216994), .Y(n40369) );
  CLKBUFX3 U28659 ( .A(net218076), .Y(n40214) );
  CLKINVX1 U28660 ( .A(net218152), .Y(net218076) );
  BUFX4 U28661 ( .A(net221840), .Y(net265644) );
  CLKINVX1 U28662 ( .A(net266218), .Y(net221840) );
  CLKBUFX3 U28663 ( .A(net216980), .Y(n40376) );
  CLKBUFX3 U28664 ( .A(net218058), .Y(n40223) );
  CLKINVX1 U28665 ( .A(net218152), .Y(net218058) );
  CLKINVX1 U28666 ( .A(net266218), .Y(net221850) );
  CLKBUFX3 U28667 ( .A(net218118), .Y(n40193) );
  CLKBUFX3 U28668 ( .A(net218130), .Y(n40187) );
  CLKBUFX3 U28669 ( .A(net216976), .Y(n40378) );
  CLKINVX1 U28670 ( .A(n40289), .Y(net216976) );
  CLKBUFX3 U28671 ( .A(net218056), .Y(n40224) );
  CLKINVX1 U28672 ( .A(net218152), .Y(net218056) );
  CLKINVX1 U28673 ( .A(net266151), .Y(net221722) );
  BUFX4 U28674 ( .A(net221812), .Y(net265378) );
  CLKINVX1 U28675 ( .A(net221984), .Y(net221744) );
  CLKINVX1 U28676 ( .A(net221962), .Y(net221762) );
  CLKINVX1 U28677 ( .A(net266218), .Y(net221844) );
  CLKBUFX3 U28678 ( .A(net217992), .Y(n40255) );
  CLKINVX1 U28679 ( .A(net218146), .Y(net217992) );
  CLKINVX1 U28680 ( .A(net218156), .Y(net218122) );
  BUFX4 U28681 ( .A(net221770), .Y(net264979) );
  CLKINVX1 U28682 ( .A(net221934), .Y(net221770) );
  CLKBUFX3 U28683 ( .A(net217202), .Y(n40278) );
  CLKBUFX3 U28684 ( .A(net217190), .Y(n40280) );
  BUFX4 U28685 ( .A(net221792), .Y(net265188) );
  CLKINVX1 U28686 ( .A(net221954), .Y(net221792) );
  OAI211X1 U28687 ( .A0(n12813), .A1(net209977), .B0(n40756), .C0(n40757), .Y(
        n40755) );
  NAND2BX1 U28688 ( .AN(net266235), .B(n51445), .Y(n40756) );
  NAND2X1 U28689 ( .A(n_cell_301249_net269763), .B(n40759), .Y(n40757) );
  AND2X2 U28690 ( .A(net172112), .B(n40753), .Y(n40752) );
  NOR3BXL U28691 ( .AN(net171523), .B(n40491), .C(net171264), .Y(n40753) );
  CLKINVX1 U28692 ( .A(net260449), .Y(net171264) );
  NOR2X1 U28693 ( .A(n40514), .B(n_cell_303546_net277506), .Y(n40516) );
  AOI21X1 U28694 ( .A0(n11544), .A1(n40515), .B0(n40513), .Y(n40514) );
  CLKINVX1 U28695 ( .A(n11543), .Y(n40513) );
  NAND2X1 U28696 ( .A(n40767), .B(n11549), .Y(n40515) );
  NAND2X1 U28697 ( .A(n11541), .B(n36929), .Y(n40633) );
  NOR2X1 U28698 ( .A(n40566), .B(n40568), .Y(n40754) );
  NOR2X1 U28699 ( .A(net264532), .B(n40569), .Y(n40568) );
  NOR2X1 U28700 ( .A(n40567), .B(net209402), .Y(n40566) );
  NAND2X1 U28701 ( .A(n10619), .B(n39937), .Y(n40569) );
  AOI21X1 U28702 ( .A0(n40540), .A1(n10626), .B0(n_cell_301249_net269758), .Y(
        n40539) );
  OAI21XL U28703 ( .A0(n39935), .A1(n40537), .B0(n10624), .Y(n40540) );
  AOI21X1 U28704 ( .A0(n40538), .A1(n11241), .B0(n_cell_303546_net277551), .Y(
        n40537) );
  CLKINVX1 U28705 ( .A(n11242), .Y(n_cell_303546_net277551) );
  NOR2X1 U28706 ( .A(net209977), .B(net171545), .Y(n40719) );
  NOR2X1 U28707 ( .A(net209402), .B(n40565), .Y(n40461) );
  NOR2X1 U28708 ( .A(n37471), .B(n40564), .Y(n40565) );
  NOR2X1 U28709 ( .A(n40562), .B(n40003), .Y(n40564) );
  NOR2X1 U28710 ( .A(n10063), .B(net217178), .Y(n39875) );
  NOR3X1 U28711 ( .A(n39616), .B(n39775), .C(n_cell_301249_net269477), .Y(
        n39774) );
  CLKINVX1 U28712 ( .A(n39839), .Y(n39775) );
  AOI21X1 U28713 ( .A0(n39617), .A1(net151779), .B0(n39618), .Y(n39616) );
  NOR3BXL U28714 ( .AN(net260449), .B(n39773), .C(n_cell_301249_net269475),
        .Y(n39839) );
  OAI21XL U28715 ( .A0(n39770), .A1(n39873), .B0(net168849), .Y(n40004) );
  NAND2X1 U28716 ( .A(n39874), .B(n10064), .Y(n39873) );
  AOI21X1 U28717 ( .A0(n39771), .A1(n39772), .B0(n10066), .Y(n39770) );
  CLKINVX1 U28718 ( .A(n10067), .Y(n39874) );
  NAND2X1 U28719 ( .A(n37348), .B(n40019), .Y(n40020) );
  OAI21XL U28720 ( .A0(n39546), .A1(n39996), .B0(n39998), .Y(n40019) );
  NOR2X1 U28721 ( .A(n11228), .B(n39999), .Y(n39998) );
  NAND2X1 U28722 ( .A(n10776), .B(n39997), .Y(n39996) );
  NOR4X1 U28723 ( .A(n40001), .B(n40002), .C(n_cell_301249_net269853), .D(
        n40003), .Y(n40000) );
  OAI2BB1X1 U28724 ( .A0N(n40034), .A1N(n39933), .B0(n37016), .Y(n39696) );
  NOR4X1 U28725 ( .A(n39934), .B(n_cell_301249_net269758), .C(n39935), .D(
        n_cell_301249_net269755), .Y(n39933) );
  OAI21XL U28726 ( .A0(n39695), .A1(n39931), .B0(n40027), .Y(n40034) );
  NAND2X1 U28727 ( .A(n9992), .B(n39932), .Y(n39931) );
  NAND2X1 U28728 ( .A(n37342), .B(n39936), .Y(n39697) );
  NOR2X1 U28729 ( .A(n39937), .B(n39938), .Y(n39936) );
  CLKINVX1 U28730 ( .A(n10619), .Y(n39938) );
  NAND2X1 U28731 ( .A(n40272), .B(net219356), .Y(net208565) );
  CLKBUFX3 U28732 ( .A(net221716), .Y(net264532) );
  CLKINVX1 U28733 ( .A(net266151), .Y(net221716) );
  CLKBUFX3 U28734 ( .A(net218746), .Y(n40096) );
  CLKBUFX3 U28735 ( .A(net218414), .Y(net262988) );
  CLKBUFX3 U28736 ( .A(net218740), .Y(n40099) );
  CLKBUFX3 U28737 ( .A(net218410), .Y(net262950) );
  CLKBUFX3 U28738 ( .A(net218742), .Y(n40098) );
  CLKBUFX3 U28739 ( .A(net218744), .Y(n40097) );
  CLKBUFX3 U28740 ( .A(net218412), .Y(net262969) );
  CLKBUFX3 U28741 ( .A(net218788), .Y(n40076) );
  CLKBUFX3 U28742 ( .A(net218790), .Y(n40075) );
  CLKBUFX3 U28743 ( .A(net218454), .Y(net263368) );
  CLKBUFX3 U28744 ( .A(net218456), .Y(net263387) );
  CLKBUFX3 U28745 ( .A(net218442), .Y(net263254) );
  CLKBUFX3 U28746 ( .A(net218772), .Y(n40083) );
  CLKBUFX3 U28747 ( .A(n42497), .Y(n42496) );
  CLKINVX1 U28748 ( .A(n43015), .Y(n42957) );
  CLKINVX1 U28749 ( .A(n43015), .Y(n42956) );
  CLKBUFX3 U28750 ( .A(net218472), .Y(net263539) );
  CLKBUFX3 U28751 ( .A(n33211), .Y(n42214) );
  CLKINVX1 U28752 ( .A(n43014), .Y(n42951) );
  CLKBUFX3 U28753 ( .A(n33219), .Y(n42213) );
  CLKINVX1 U28754 ( .A(n43014), .Y(n42950) );
  CLKINVX1 U28755 ( .A(n43012), .Y(n42909) );
  CLKBUFX3 U28756 ( .A(n33807), .Y(n41881) );
  CLKBUFX3 U28757 ( .A(n33815), .Y(n41880) );
  CLKBUFX3 U28758 ( .A(n33823), .Y(n41879) );
  CLKBUFX3 U28759 ( .A(net218504), .Y(net263843) );
  CLKBUFX3 U28760 ( .A(net218502), .Y(net263824) );
  CLKBUFX3 U28761 ( .A(net218506), .Y(net263862) );
  CLKBUFX3 U28762 ( .A(net218214), .Y(n40154) );
  CLKBUFX3 U28763 ( .A(net221952), .Y(net266738) );
  CLKBUFX3 U28764 ( .A(net217140), .Y(n40304) );
  CLKBUFX3 U28765 ( .A(net218500), .Y(net263805) );
  CLKBUFX3 U28766 ( .A(net217176), .Y(n40286) );
  CLKBUFX3 U28767 ( .A(net218430), .Y(net263140) );
  CLKBUFX3 U28768 ( .A(net218426), .Y(net263102) );
  CLKBUFX3 U28769 ( .A(net218416), .Y(net263007) );
  CLKBUFX3 U28770 ( .A(net218428), .Y(net263121) );
  CLKBUFX3 U28771 ( .A(net218192), .Y(n40165) );
  CLKBUFX3 U28772 ( .A(net218190), .Y(n40166) );
  BUFX4 U28773 ( .A(net221934), .Y(net266549) );
  CLKBUFX3 U28774 ( .A(net218432), .Y(net263159) );
  CLKBUFX3 U28775 ( .A(net218420), .Y(net263045) );
  CLKBUFX3 U28776 ( .A(net218194), .Y(n40164) );
  CLKBUFX3 U28777 ( .A(net221936), .Y(net266570) );
  CLKBUFX3 U28778 ( .A(net218750), .Y(n40094) );
  CLKBUFX3 U28779 ( .A(net218418), .Y(net263026) );
  CLKBUFX3 U28780 ( .A(net218458), .Y(net263406) );
  CLKBUFX3 U28781 ( .A(net218424), .Y(net263083) );
  CLKBUFX3 U28782 ( .A(net218218), .Y(n40152) );
  CLKBUFX3 U28783 ( .A(net217172), .Y(n40288) );
  CLKBUFX3 U28784 ( .A(net218422), .Y(net263064) );
  CLKBUFX3 U28785 ( .A(net218198), .Y(n40162) );
  CLKBUFX3 U28786 ( .A(net218200), .Y(n40161) );
  CLKBUFX3 U28787 ( .A(net221940), .Y(net266612) );
  CLKBUFX3 U28788 ( .A(net217168), .Y(n40290) );
  CLKBUFX3 U28789 ( .A(net218464), .Y(net263463) );
  CLKBUFX3 U28790 ( .A(n33131), .Y(n42224) );
  CLKBUFX3 U28791 ( .A(net218212), .Y(n40155) );
  CLKBUFX3 U28792 ( .A(net218478), .Y(net263596) );
  CLKBUFX3 U28793 ( .A(n33135), .Y(n41965) );
  CLKBUFX3 U28794 ( .A(n33147), .Y(n42222) );
  CLKBUFX3 U28795 ( .A(n33151), .Y(n41963) );
  CLKBUFX3 U28796 ( .A(net218476), .Y(net263577) );
  CLKBUFX3 U28797 ( .A(n33203), .Y(n42215) );
  CLKBUFX3 U28798 ( .A(n33155), .Y(n42221) );
  CLKBUFX3 U28799 ( .A(n33187), .Y(n42217) );
  CLKBUFX3 U28800 ( .A(n33195), .Y(n42216) );
  CLKBUFX3 U28801 ( .A(n33179), .Y(n42218) );
  CLKBUFX3 U28802 ( .A(n33163), .Y(n42220) );
  CLKBUFX3 U28803 ( .A(n33171), .Y(n42219) );
  CLKBUFX3 U28804 ( .A(net218210), .Y(n40156) );
  CLKBUFX3 U28805 ( .A(net217134), .Y(n40307) );
  CLKBUFX3 U28806 ( .A(n33191), .Y(n41958) );
  CLKBUFX3 U28807 ( .A(n33199), .Y(n41957) );
  CLKBUFX3 U28808 ( .A(n33183), .Y(n41959) );
  CLKBUFX3 U28809 ( .A(net221950), .Y(net266717) );
  CLKBUFX3 U28810 ( .A(n33175), .Y(n41960) );
  CLKBUFX3 U28811 ( .A(net218474), .Y(net263558) );
  CLKBUFX3 U28812 ( .A(n33167), .Y(n41961) );
  CLKBUFX3 U28813 ( .A(n33159), .Y(n41962) );
  CLKBUFX3 U28814 ( .A(n33215), .Y(n41955) );
  CLKBUFX3 U28815 ( .A(n33223), .Y(n41954) );
  CLKBUFX3 U28816 ( .A(n33207), .Y(n41956) );
  CLKBUFX3 U28817 ( .A(n33239), .Y(n41952) );
  CLKBUFX3 U28818 ( .A(n33247), .Y(n41951) );
  CLKBUFX3 U28819 ( .A(n33231), .Y(n41953) );
  CLKBUFX3 U28820 ( .A(net218468), .Y(net263501) );
  CLKBUFX3 U28821 ( .A(n33227), .Y(n42212) );
  CLKBUFX3 U28822 ( .A(n33235), .Y(n42211) );
  CLKBUFX3 U28823 ( .A(n33243), .Y(n42210) );
  CLKBUFX3 U28824 ( .A(net218434), .Y(net263178) );
  CLKBUFX3 U28825 ( .A(net218450), .Y(net263330) );
  CLKBUFX3 U28826 ( .A(net218196), .Y(n40163) );
  CLKBUFX3 U28827 ( .A(net221938), .Y(net266591) );
  CLKBUFX3 U28828 ( .A(net217166), .Y(n40291) );
  CLKBUFX3 U28829 ( .A(net218202), .Y(n40160) );
  CLKBUFX3 U28830 ( .A(net221942), .Y(net266633) );
  CLKBUFX3 U28831 ( .A(net218216), .Y(n40153) );
  CLKBUFX3 U28832 ( .A(net217138), .Y(n40305) );
  CLKBUFX3 U28833 ( .A(net221954), .Y(net266759) );
  CLKBUFX3 U28834 ( .A(net218932), .Y(net218610) );
  CLKBUFX3 U28835 ( .A(n33799), .Y(n41882) );
  CLKBUFX3 U28836 ( .A(n33791), .Y(n41883) );
  INVX4 U28837 ( .A(n49523), .Y(n37597) );
  CLKBUFX3 U28838 ( .A(n34407), .Y(n41807) );
  CLKBUFX3 U28839 ( .A(n33575), .Y(n41910) );
  CLKINVX1 U28840 ( .A(n43023), .Y(n42861) );
  CLKBUFX3 U28841 ( .A(net218614), .Y(n40150) );
  CLKINVX1 U28842 ( .A(n43023), .Y(n42846) );
  CLKBUFX3 U28843 ( .A(net218298), .Y(net261886) );
  CLKBUFX3 U28844 ( .A(n34335), .Y(n41815) );
  CLKBUFX3 U28845 ( .A(n34343), .Y(n41814) );
  CLKBUFX3 U28846 ( .A(n34327), .Y(n41816) );
  CLKBUFX3 U28847 ( .A(n34311), .Y(n41818) );
  CLKBUFX3 U28848 ( .A(n34319), .Y(n41817) );
  CLKBUFX3 U28849 ( .A(n34303), .Y(n41819) );
  CLKBUFX3 U28850 ( .A(n34295), .Y(n41820) );
  CLKBUFX3 U28851 ( .A(n34279), .Y(n41822) );
  CLKBUFX3 U28852 ( .A(n34287), .Y(n41821) );
  CLKBUFX3 U28853 ( .A(n34271), .Y(n41823) );
  CLKBUFX3 U28854 ( .A(n34255), .Y(n41825) );
  CLKBUFX3 U28855 ( .A(n34263), .Y(n41824) );
  CLKBUFX3 U28856 ( .A(n34247), .Y(n41826) );
  CLKBUFX3 U28857 ( .A(n34239), .Y(n41827) );
  CLKBUFX3 U28858 ( .A(n34223), .Y(n41829) );
  CLKBUFX3 U28859 ( .A(n34231), .Y(n41828) );
  CLKBUFX3 U28860 ( .A(n34215), .Y(n41830) );
  CLKBUFX3 U28861 ( .A(n34199), .Y(n41832) );
  CLKBUFX3 U28862 ( .A(n34207), .Y(n41831) );
  CLKBUFX3 U28863 ( .A(n34191), .Y(n41833) );
  CLKBUFX3 U28864 ( .A(n34175), .Y(n41835) );
  CLKBUFX3 U28865 ( .A(n34183), .Y(n41834) );
  CLKBUFX3 U28866 ( .A(n34167), .Y(n41836) );
  CLKBUFX3 U28867 ( .A(n34159), .Y(n41837) );
  CLKBUFX3 U28868 ( .A(n34151), .Y(n41838) );
  CLKBUFX3 U28869 ( .A(n34143), .Y(n41839) );
  CLKBUFX3 U28870 ( .A(n34135), .Y(n41840) );
  CLKBUFX3 U28871 ( .A(n34127), .Y(n41841) );
  CLKBUFX3 U28872 ( .A(n34119), .Y(n41842) );
  CLKBUFX3 U28873 ( .A(n34111), .Y(n41843) );
  CLKBUFX3 U28874 ( .A(n34015), .Y(n41855) );
  CLKBUFX3 U28875 ( .A(n33943), .Y(n41864) );
  CLKBUFX3 U28876 ( .A(n33879), .Y(n41872) );
  CLKBUFX3 U28877 ( .A(n33887), .Y(n41871) );
  CLKBUFX3 U28878 ( .A(n33551), .Y(n41913) );
  CLKBUFX3 U28879 ( .A(n33543), .Y(n41914) );
  CLKBUFX3 U28880 ( .A(n33559), .Y(n41912) );
  CLKBUFX3 U28881 ( .A(n34387), .Y(n42067) );
  CLKBUFX3 U28882 ( .A(n34379), .Y(n42068) );
  CLKBUFX3 U28883 ( .A(net218696), .Y(n40116) );
  CLKBUFX3 U28884 ( .A(n34371), .Y(n42069) );
  CLKBUFX3 U28885 ( .A(n34363), .Y(n42070) );
  CLKBUFX3 U28886 ( .A(n34355), .Y(n42071) );
  CLKBUFX3 U28887 ( .A(n34347), .Y(n42072) );
  CLKBUFX3 U28888 ( .A(net218700), .Y(n40114) );
  CLKBUFX3 U28889 ( .A(net218374), .Y(net262608) );
  CLKBUFX3 U28890 ( .A(net218176), .Y(n40173) );
  CLKBUFX3 U28891 ( .A(n34331), .Y(n42074) );
  CLKBUFX3 U28892 ( .A(n34323), .Y(n42075) );
  CLKBUFX3 U28893 ( .A(net218702), .Y(n40113) );
  CLKBUFX3 U28894 ( .A(net218376), .Y(net262627) );
  CLKBUFX3 U28895 ( .A(n34315), .Y(n42076) );
  CLKBUFX3 U28896 ( .A(net218704), .Y(n40112) );
  CLKBUFX3 U28897 ( .A(net218378), .Y(net262646) );
  CLKBUFX3 U28898 ( .A(n34307), .Y(n42077) );
  CLKBUFX3 U28899 ( .A(n34299), .Y(n42078) );
  CLKBUFX3 U28900 ( .A(n34291), .Y(n42079) );
  CLKBUFX3 U28901 ( .A(net218352), .Y(net262399) );
  CLKBUFX3 U28902 ( .A(n34283), .Y(n42080) );
  CLKBUFX3 U28903 ( .A(net218676), .Y(n40122) );
  CLKBUFX3 U28904 ( .A(n34275), .Y(n42081) );
  CLKBUFX3 U28905 ( .A(net221922), .Y(net266423) );
  CLKBUFX3 U28906 ( .A(net218354), .Y(net262418) );
  CLKBUFX3 U28907 ( .A(net217146), .Y(n40301) );
  CLKBUFX3 U28908 ( .A(n34267), .Y(n42082) );
  CLKBUFX3 U28909 ( .A(net218678), .Y(n40121) );
  CLKBUFX3 U28910 ( .A(net218178), .Y(n40172) );
  CLKBUFX3 U28911 ( .A(n34259), .Y(n42083) );
  CLKBUFX3 U28912 ( .A(net218356), .Y(net262437) );
  CLKBUFX3 U28913 ( .A(n34251), .Y(n42084) );
  CLKBUFX3 U28914 ( .A(net218680), .Y(n40120) );
  CLKBUFX3 U28915 ( .A(n34243), .Y(n42085) );
  CLKBUFX3 U28916 ( .A(net218358), .Y(net262456) );
  CLKBUFX3 U28917 ( .A(n34235), .Y(n42086) );
  CLKBUFX3 U28918 ( .A(n34227), .Y(n42087) );
  CLKBUFX3 U28919 ( .A(net218684), .Y(n40119) );
  CLKBUFX3 U28920 ( .A(n34219), .Y(n42088) );
  CLKBUFX3 U28921 ( .A(net218360), .Y(net262475) );
  CLKBUFX3 U28922 ( .A(n34211), .Y(n42089) );
  CLKBUFX3 U28923 ( .A(n34203), .Y(n42090) );
  CLKBUFX3 U28924 ( .A(net221924), .Y(net266444) );
  CLKBUFX3 U28925 ( .A(n34195), .Y(n42091) );
  CLKBUFX3 U28926 ( .A(net217148), .Y(n40300) );
  CLKBUFX3 U28927 ( .A(net218688), .Y(n40118) );
  CLKBUFX3 U28928 ( .A(n34187), .Y(n42092) );
  CLKBUFX3 U28929 ( .A(n34179), .Y(n42093) );
  CLKBUFX3 U28930 ( .A(n34171), .Y(n42094) );
  BUFX4 U28931 ( .A(net218394), .Y(net262798) );
  CLKBUFX3 U28932 ( .A(n34115), .Y(n42101) );
  CLKBUFX3 U28933 ( .A(n34099), .Y(n42103) );
  CLKBUFX3 U28934 ( .A(n34107), .Y(n42102) );
  CLKBUFX3 U28935 ( .A(n34091), .Y(n42104) );
  CLKINVX1 U28936 ( .A(n43020), .Y(n42805) );
  CLKBUFX3 U28937 ( .A(net218708), .Y(n40111) );
  CLKBUFX3 U28938 ( .A(net218380), .Y(net262665) );
  CLKBUFX3 U28939 ( .A(n34011), .Y(n42114) );
  CLKBUFX3 U28940 ( .A(net218346), .Y(net262342) );
  CLKBUFX3 U28941 ( .A(n33839), .Y(n41877) );
  CLKBUFX3 U28942 ( .A(n33863), .Y(n41874) );
  CLKBUFX3 U28943 ( .A(n33855), .Y(n41875) );
  CLKBUFX3 U28944 ( .A(n33871), .Y(n41873) );
  CLKBUFX3 U28945 ( .A(n33831), .Y(n41878) );
  CLKBUFX3 U28946 ( .A(n33735), .Y(n41890) );
  CLKINVX1 U28947 ( .A(n43017), .Y(n42753) );
  CLKBUFX3 U28948 ( .A(n33727), .Y(n41891) );
  CLKBUFX3 U28949 ( .A(n33719), .Y(n41892) );
  CLKBUFX3 U28950 ( .A(n33535), .Y(n41915) );
  CLKINVX1 U28951 ( .A(n43017), .Y(n42750) );
  CLKBUFX3 U28952 ( .A(n33527), .Y(n41916) );
  CLKBUFX3 U28953 ( .A(n33875), .Y(n42131) );
  CLKBUFX3 U28954 ( .A(n33867), .Y(n42132) );
  CLKBUFX3 U28955 ( .A(n33859), .Y(n42133) );
  CLKBUFX3 U28956 ( .A(n33851), .Y(n42134) );
  CLKBUFX3 U28957 ( .A(net218316), .Y(net262057) );
  CLKBUFX3 U28958 ( .A(n33843), .Y(n42135) );
  CLKBUFX3 U28959 ( .A(net218636), .Y(n40140) );
  CLKBUFX3 U28960 ( .A(net217158), .Y(n40295) );
  CLKBUFX3 U28961 ( .A(n33835), .Y(n42136) );
  CLKBUFX3 U28962 ( .A(net221910), .Y(net266297) );
  CLKBUFX3 U28963 ( .A(n33819), .Y(n42138) );
  CLKBUFX3 U28964 ( .A(n33827), .Y(n42137) );
  CLKBUFX3 U28965 ( .A(n33811), .Y(n42139) );
  CLKBUFX3 U28966 ( .A(net218640), .Y(n40139) );
  CLKBUFX3 U28967 ( .A(net218320), .Y(net262095) );
  CLKBUFX3 U28968 ( .A(n33731), .Y(n42149) );
  CLKBUFX3 U28969 ( .A(net218618), .Y(n40148) );
  CLKBUFX3 U28970 ( .A(n33723), .Y(n42150) );
  CLKBUFX3 U28971 ( .A(net218302), .Y(net261924) );
  CLKBUFX3 U28972 ( .A(n33715), .Y(n42151) );
  CLKBUFX3 U28973 ( .A(net218674), .Y(n40123) );
  CLKBUFX3 U28974 ( .A(net218350), .Y(net262380) );
  CLKBUFX3 U28975 ( .A(n33523), .Y(n42175) );
  CLKBUFX3 U28976 ( .A(net218330), .Y(net262190) );
  CLKBUFX3 U28977 ( .A(n34031), .Y(n41853) );
  CLKBUFX3 U28978 ( .A(n34055), .Y(n41850) );
  CLKBUFX3 U28979 ( .A(n34023), .Y(n41854) );
  CLKBUFX3 U28980 ( .A(n34039), .Y(n41852) );
  CLKBUFX3 U28981 ( .A(n34047), .Y(n41851) );
  CLKBUFX3 U28982 ( .A(net218736), .Y(n40101) );
  CLKBUFX3 U28983 ( .A(net218406), .Y(net262912) );
  CLKBUFX3 U28984 ( .A(n33999), .Y(n41857) );
  CLKBUFX3 U28985 ( .A(n34007), .Y(n41856) );
  CLKINVX1 U28986 ( .A(n43021), .Y(n42811) );
  CLKBUFX3 U28987 ( .A(n34035), .Y(n42111) );
  CLKBUFX3 U28988 ( .A(n34027), .Y(n42112) );
  CLKBUFX3 U28989 ( .A(n34019), .Y(n42113) );
  CLKBUFX3 U28990 ( .A(net218738), .Y(n40100) );
  CLKBUFX3 U28991 ( .A(net218408), .Y(net262931) );
  CLKBUFX3 U28992 ( .A(n34003), .Y(n42115) );
  CLKBUFX3 U28993 ( .A(n34079), .Y(n41847) );
  CLKBUFX3 U28994 ( .A(n34071), .Y(n41848) );
  CLKBUFX3 U28995 ( .A(n34063), .Y(n41849) );
  CLKBUFX3 U28996 ( .A(n34103), .Y(n41844) );
  CLKBUFX3 U28997 ( .A(n34095), .Y(n41845) );
  CLKBUFX3 U28998 ( .A(n34087), .Y(n41846) );
  CLKBUFX3 U28999 ( .A(n33967), .Y(n41861) );
  CLKBUFX3 U29000 ( .A(n33959), .Y(n41862) );
  CLKBUFX3 U29001 ( .A(n33975), .Y(n41860) );
  CLKBUFX3 U29002 ( .A(n33983), .Y(n41859) );
  CLKBUFX3 U29003 ( .A(n33991), .Y(n41858) );
  CLKBUFX3 U29004 ( .A(n33903), .Y(n41869) );
  CLKBUFX3 U29005 ( .A(n33919), .Y(n41867) );
  CLKBUFX3 U29006 ( .A(n33927), .Y(n41866) );
  CLKBUFX3 U29007 ( .A(n33935), .Y(n41865) );
  CLKBUFX3 U29008 ( .A(n33895), .Y(n41870) );
  CLKBUFX3 U29009 ( .A(net218720), .Y(n40107) );
  CLKBUFX3 U29010 ( .A(n33759), .Y(n41887) );
  CLKBUFX3 U29011 ( .A(n33751), .Y(n41888) );
  CLKBUFX3 U29012 ( .A(n33743), .Y(n41889) );
  CLKBUFX3 U29013 ( .A(n33775), .Y(n41885) );
  CLKBUFX3 U29014 ( .A(n33767), .Y(n41886) );
  CLKBUFX3 U29015 ( .A(n33783), .Y(n41884) );
  CLKBUFX3 U29016 ( .A(n33711), .Y(n41893) );
  CLKBUFX3 U29017 ( .A(net218620), .Y(n40147) );
  CLKBUFX3 U29018 ( .A(n33703), .Y(n41894) );
  CLKBUFX3 U29019 ( .A(n33695), .Y(n41895) );
  CLKBUFX3 U29020 ( .A(n33687), .Y(n41896) );
  BUFX4 U29021 ( .A(net217164), .Y(n40292) );
  CLKBUFX3 U29022 ( .A(n33679), .Y(n41897) );
  CLKBUFX3 U29023 ( .A(n33671), .Y(n41898) );
  CLKBUFX3 U29024 ( .A(n33663), .Y(n41899) );
  CLKBUFX3 U29025 ( .A(n33647), .Y(n41901) );
  CLKBUFX3 U29026 ( .A(n33655), .Y(n41900) );
  CLKBUFX3 U29027 ( .A(n33639), .Y(n41902) );
  CLKBUFX3 U29028 ( .A(n33631), .Y(n41903) );
  CLKINVX1 U29029 ( .A(n43009), .Y(n42737) );
  CLKBUFX3 U29030 ( .A(n33607), .Y(n41906) );
  CLKBUFX3 U29031 ( .A(n33615), .Y(n41905) );
  CLKBUFX3 U29032 ( .A(n33623), .Y(n41904) );
  CLKBUFX3 U29033 ( .A(n33599), .Y(n41907) );
  CLKBUFX3 U29034 ( .A(n33591), .Y(n41908) );
  CLKBUFX3 U29035 ( .A(n33583), .Y(n41909) );
  CLKBUFX3 U29036 ( .A(n33503), .Y(n41919) );
  CLKBUFX3 U29037 ( .A(n33511), .Y(n41918) );
  CLKBUFX3 U29038 ( .A(n33519), .Y(n41917) );
  CLKBUFX3 U29039 ( .A(n33495), .Y(n41920) );
  CLKBUFX3 U29040 ( .A(net218324), .Y(net262133) );
  CLKINVX1 U29041 ( .A(n43019), .Y(n42784) );
  CLKBUFX3 U29042 ( .A(n33463), .Y(n41924) );
  CLKBUFX3 U29043 ( .A(n33471), .Y(n41923) );
  CLKBUFX3 U29044 ( .A(n33487), .Y(n41921) );
  CLKBUFX3 U29045 ( .A(n33479), .Y(n41922) );
  CLKBUFX3 U29046 ( .A(net218648), .Y(n40135) );
  CLKBUFX3 U29047 ( .A(n34139), .Y(n42098) );
  CLKBUFX3 U29048 ( .A(n34131), .Y(n42099) );
  CLKBUFX3 U29049 ( .A(n34123), .Y(n42100) );
  CLKBUFX3 U29050 ( .A(net217150), .Y(n40299) );
  CLKBUFX3 U29051 ( .A(net218182), .Y(n40170) );
  CLKBUFX3 U29052 ( .A(n34163), .Y(n42095) );
  CLKBUFX3 U29053 ( .A(net221926), .Y(net266465) );
  CLKBUFX3 U29054 ( .A(n34147), .Y(n42097) );
  CLKBUFX3 U29055 ( .A(n34155), .Y(n42096) );
  CLKBUFX3 U29056 ( .A(net218724), .Y(n40105) );
  CLKBUFX3 U29057 ( .A(net218396), .Y(net262817) );
  CLKBUFX3 U29058 ( .A(n34059), .Y(n42108) );
  CLKBUFX3 U29059 ( .A(n34051), .Y(n42109) );
  CLKBUFX3 U29060 ( .A(n34043), .Y(n42110) );
  CLKBUFX3 U29061 ( .A(net218184), .Y(n40169) );
  CLKBUFX3 U29062 ( .A(n34067), .Y(n42107) );
  CLKBUFX3 U29063 ( .A(n34075), .Y(n42106) );
  CLKBUFX3 U29064 ( .A(n34083), .Y(n42105) );
  CLKBUFX3 U29065 ( .A(net221928), .Y(net266486) );
  CLKBUFX3 U29066 ( .A(n33995), .Y(n42116) );
  CLKBUFX3 U29067 ( .A(net218186), .Y(n40168) );
  CLKBUFX3 U29068 ( .A(n33987), .Y(n42117) );
  CLKBUFX3 U29069 ( .A(net217154), .Y(n40297) );
  CLKBUFX3 U29070 ( .A(n33979), .Y(n42118) );
  CLKBUFX3 U29071 ( .A(n33971), .Y(n42119) );
  CLKBUFX3 U29072 ( .A(net218716), .Y(n40108) );
  CLKBUFX3 U29073 ( .A(net218388), .Y(net262741) );
  CLKBUFX3 U29074 ( .A(n33963), .Y(n42120) );
  CLKBUFX3 U29075 ( .A(net221930), .Y(net266507) );
  CLKBUFX3 U29076 ( .A(net218188), .Y(n40167) );
  CLKBUFX3 U29077 ( .A(n33955), .Y(n42121) );
  CLKBUFX3 U29078 ( .A(n33939), .Y(n42123) );
  CLKBUFX3 U29079 ( .A(net221932), .Y(net266528) );
  CLKBUFX3 U29080 ( .A(n33931), .Y(n42124) );
  CLKBUFX3 U29081 ( .A(net218722), .Y(n40106) );
  CLKBUFX3 U29082 ( .A(net218392), .Y(net262779) );
  CLKBUFX3 U29083 ( .A(n33899), .Y(n42128) );
  CLKBUFX3 U29084 ( .A(n33891), .Y(n42129) );
  CLKBUFX3 U29085 ( .A(net218164), .Y(n40179) );
  CLKBUFX3 U29086 ( .A(n33907), .Y(n42127) );
  CLKBUFX3 U29087 ( .A(net217156), .Y(n40296) );
  CLKBUFX3 U29088 ( .A(n33915), .Y(n42126) );
  CLKBUFX3 U29089 ( .A(n33923), .Y(n42125) );
  CLKBUFX3 U29090 ( .A(net218162), .Y(n40180) );
  CLKBUFX3 U29091 ( .A(n33803), .Y(n42140) );
  CLKBUFX3 U29092 ( .A(n33795), .Y(n42141) );
  CLKBUFX3 U29093 ( .A(net218642), .Y(n40138) );
  CLKBUFX3 U29094 ( .A(net218322), .Y(net262114) );
  CLKBUFX3 U29095 ( .A(n33787), .Y(n42142) );
  CLKBUFX3 U29096 ( .A(n33755), .Y(n42146) );
  CLKBUFX3 U29097 ( .A(n33747), .Y(n42147) );
  CLKBUFX3 U29098 ( .A(n33739), .Y(n42148) );
  CLKBUFX3 U29099 ( .A(net217160), .Y(n40294) );
  CLKBUFX3 U29100 ( .A(net218160), .Y(n40181) );
  CLKBUFX3 U29101 ( .A(n33779), .Y(n42143) );
  CLKBUFX3 U29102 ( .A(n33771), .Y(n42144) );
  CLKBUFX3 U29103 ( .A(n33763), .Y(n42145) );
  CLKBUFX3 U29104 ( .A(n33707), .Y(n42152) );
  CLKBUFX3 U29105 ( .A(n33699), .Y(n42153) );
  CLKBUFX3 U29106 ( .A(net218622), .Y(n40146) );
  CLKBUFX3 U29107 ( .A(net218304), .Y(net261943) );
  CLKBUFX3 U29108 ( .A(net217162), .Y(n40293) );
  CLKBUFX3 U29109 ( .A(n33691), .Y(n42154) );
  CLKBUFX3 U29110 ( .A(net221906), .Y(net266255) );
  CLKBUFX3 U29111 ( .A(n33683), .Y(n42155) );
  CLKBUFX3 U29112 ( .A(net221908), .Y(net266276) );
  CLKBUFX3 U29113 ( .A(net218624), .Y(n40145) );
  CLKBUFX3 U29114 ( .A(n33675), .Y(n42156) );
  CLKBUFX3 U29115 ( .A(net218308), .Y(net261981) );
  CLKBUFX3 U29116 ( .A(n33667), .Y(n42157) );
  CLKINVX1 U29117 ( .A(n43018), .Y(n42763) );
  CLKBUFX3 U29118 ( .A(n33659), .Y(n42158) );
  CLKBUFX3 U29119 ( .A(n33651), .Y(n42159) );
  CLKBUFX3 U29120 ( .A(n33643), .Y(n42160) );
  CLKBUFX3 U29121 ( .A(net221912), .Y(net266318) );
  CLKBUFX3 U29122 ( .A(net218166), .Y(n40178) );
  CLKBUFX3 U29123 ( .A(n33627), .Y(n42162) );
  CLKBUFX3 U29124 ( .A(n33579), .Y(n42168) );
  CLKBUFX3 U29125 ( .A(n33619), .Y(n42163) );
  CLKBUFX3 U29126 ( .A(n33611), .Y(n42164) );
  CLKBUFX3 U29127 ( .A(n33603), .Y(n42165) );
  CLKBUFX3 U29128 ( .A(n33595), .Y(n42166) );
  CLKBUFX3 U29129 ( .A(n33587), .Y(n42167) );
  CLKBUFX3 U29130 ( .A(net218664), .Y(n40128) );
  CLKBUFX3 U29131 ( .A(net218342), .Y(net262304) );
  CLKINVX1 U29132 ( .A(n43010), .Y(n42738) );
  CLKBUFX3 U29133 ( .A(n33539), .Y(n42173) );
  CLKBUFX3 U29134 ( .A(n33547), .Y(n42172) );
  CLKBUFX3 U29135 ( .A(n33531), .Y(n42174) );
  CLKBUFX3 U29136 ( .A(n33563), .Y(n42170) );
  CLKBUFX3 U29137 ( .A(n33555), .Y(n42171) );
  CLKBUFX3 U29138 ( .A(n33571), .Y(n42169) );
  CLKBUFX3 U29139 ( .A(net221914), .Y(net266339) );
  CLKBUFX3 U29140 ( .A(net217128), .Y(n40309) );
  CLKBUFX3 U29141 ( .A(net218670), .Y(n40125) );
  CLKBUFX3 U29142 ( .A(net218348), .Y(net262361) );
  CLKBUFX3 U29143 ( .A(n33507), .Y(n42177) );
  CLKBUFX3 U29144 ( .A(n33515), .Y(n42176) );
  CLKBUFX3 U29145 ( .A(net218170), .Y(n40176) );
  CLKBUFX3 U29146 ( .A(n33499), .Y(n42178) );
  CLKBUFX3 U29147 ( .A(n33491), .Y(n42179) );
  CLKBUFX3 U29148 ( .A(net218326), .Y(net262152) );
  CLKBUFX3 U29149 ( .A(n33459), .Y(n42183) );
  CLKBUFX3 U29150 ( .A(net221916), .Y(net266360) );
  CLKBUFX3 U29151 ( .A(net217126), .Y(n40310) );
  CLKBUFX3 U29152 ( .A(n33467), .Y(n42182) );
  CLKBUFX3 U29153 ( .A(n33483), .Y(n42180) );
  CLKBUFX3 U29154 ( .A(n33475), .Y(n42181) );
  CLKBUFX3 U29155 ( .A(net218650), .Y(n40134) );
  CLKBUFX3 U29156 ( .A(net218328), .Y(net262171) );
  CLKBUFX3 U29157 ( .A(n33447), .Y(n41926) );
  CLKBUFX3 U29158 ( .A(n33439), .Y(n41927) );
  CLKBUFX3 U29159 ( .A(n33455), .Y(n41925) );
  CLKBUFX3 U29160 ( .A(n33431), .Y(n41928) );
  CLKBUFX3 U29161 ( .A(net218334), .Y(net262228) );
  CLKBUFX3 U29162 ( .A(n33407), .Y(n41931) );
  CLKBUFX3 U29163 ( .A(n33423), .Y(n41929) );
  CLKBUFX3 U29164 ( .A(n33415), .Y(n41930) );
  CLKBUFX3 U29165 ( .A(net221944), .Y(net266654) );
  CLKBUFX3 U29166 ( .A(n33399), .Y(n41932) );
  CLKBUFX3 U29167 ( .A(n33391), .Y(n41933) );
  CLKBUFX3 U29168 ( .A(n33383), .Y(n41934) );
  CLKBUFX3 U29169 ( .A(n33375), .Y(n41935) );
  CLKBUFX3 U29170 ( .A(n33367), .Y(n41936) );
  CLKBUFX3 U29171 ( .A(n33319), .Y(n41942) );
  CLKBUFX3 U29172 ( .A(n33327), .Y(n41941) );
  CLKBUFX3 U29173 ( .A(n33359), .Y(n41937) );
  CLKBUFX3 U29174 ( .A(n33351), .Y(n41938) );
  CLKBUFX3 U29175 ( .A(n33343), .Y(n41939) );
  CLKBUFX3 U29176 ( .A(n33335), .Y(n41940) );
  CLKBUFX3 U29177 ( .A(n33311), .Y(n41943) );
  CLKBUFX3 U29178 ( .A(n33443), .Y(n42185) );
  CLKBUFX3 U29179 ( .A(n33451), .Y(n42184) );
  CLKBUFX3 U29180 ( .A(n33435), .Y(n42186) );
  CLKBUFX3 U29181 ( .A(net218332), .Y(net262209) );
  CLKBUFX3 U29182 ( .A(n33427), .Y(n42187) );
  CLKBUFX3 U29183 ( .A(net217124), .Y(n40311) );
  CLKBUFX3 U29184 ( .A(net218172), .Y(n40175) );
  CLKBUFX3 U29185 ( .A(n33403), .Y(n42190) );
  CLKBUFX3 U29186 ( .A(n33419), .Y(n42188) );
  CLKBUFX3 U29187 ( .A(n33411), .Y(n42189) );
  CLKBUFX3 U29188 ( .A(net218336), .Y(net262247) );
  CLKBUFX3 U29189 ( .A(n33395), .Y(n42191) );
  CLKBUFX3 U29190 ( .A(n33387), .Y(n42192) );
  CLKBUFX3 U29191 ( .A(net218204), .Y(n40159) );
  CLKBUFX3 U29192 ( .A(n33379), .Y(n42193) );
  CLKBUFX3 U29193 ( .A(n33371), .Y(n42194) );
  CLKBUFX3 U29194 ( .A(n33363), .Y(n42195) );
  CLKBUFX3 U29195 ( .A(net217122), .Y(n40312) );
  CLKBUFX3 U29196 ( .A(n33355), .Y(n42196) );
  CLKBUFX3 U29197 ( .A(n33347), .Y(n42197) );
  CLKBUFX3 U29198 ( .A(n33339), .Y(n42198) );
  CLKBUFX3 U29199 ( .A(n33331), .Y(n42199) );
  CLKBUFX3 U29200 ( .A(n33323), .Y(n42200) );
  CLKBUFX3 U29201 ( .A(net221946), .Y(net266675) );
  CLKBUFX3 U29202 ( .A(n33315), .Y(n42201) );
  CLKBUFX3 U29203 ( .A(net218206), .Y(n40158) );
  CLKBUFX3 U29204 ( .A(n33307), .Y(n42202) );
  CLKBUFX3 U29205 ( .A(n33303), .Y(n41944) );
  CLKBUFX3 U29206 ( .A(n33255), .Y(n41950) );
  CLKBUFX3 U29207 ( .A(n33263), .Y(n41949) );
  CLKBUFX3 U29208 ( .A(n33295), .Y(n41945) );
  CLKBUFX3 U29209 ( .A(n33287), .Y(n41946) );
  CLKBUFX3 U29210 ( .A(n33279), .Y(n41947) );
  CLKBUFX3 U29211 ( .A(n33271), .Y(n41948) );
  CLKBUFX3 U29212 ( .A(n33299), .Y(n42203) );
  CLKBUFX3 U29213 ( .A(net218832), .Y(n40055) );
  CLKBUFX3 U29214 ( .A(n33251), .Y(n42209) );
  CLKBUFX3 U29215 ( .A(n33267), .Y(n42207) );
  CLKBUFX3 U29216 ( .A(n33259), .Y(n42208) );
  CLKBUFX3 U29217 ( .A(net218208), .Y(n40157) );
  CLKBUFX3 U29218 ( .A(net217132), .Y(n40308) );
  CLKBUFX3 U29219 ( .A(n33291), .Y(n42204) );
  CLKBUFX3 U29220 ( .A(net221948), .Y(net266696) );
  CLKBUFX3 U29221 ( .A(n33283), .Y(n42205) );
  CLKBUFX3 U29222 ( .A(n33275), .Y(n42206) );
  CLKBUFX3 U29223 ( .A(net221822), .Y(net265473) );
  INVX3 U29224 ( .A(n33908), .Y(n51412) );
  INVX3 U29225 ( .A(n33916), .Y(n51413) );
  CLKINVX1 U29226 ( .A(n40313), .Y(net217092) );
  CLKBUFX3 U29227 ( .A(net218012), .Y(n40245) );
  CLKINVX1 U29228 ( .A(net218148), .Y(net218012) );
  CLKBUFX3 U29229 ( .A(net221786), .Y(net265131) );
  CLKINVX1 U29230 ( .A(net221910), .Y(net221786) );
  CLKBUFX3 U29231 ( .A(net218626), .Y(n40144) );
  INVX3 U29232 ( .A(n33604), .Y(n51374) );
  CLKBUFX3 U29233 ( .A(net218344), .Y(net262323) );
  CLKBUFX3 U29234 ( .A(net217062), .Y(n40339) );
  CLKINVX1 U29235 ( .A(n40314), .Y(net217062) );
  CLKBUFX3 U29236 ( .A(net217982), .Y(n40260) );
  CLKINVX1 U29237 ( .A(net218146), .Y(net217982) );
  CLKBUFX3 U29238 ( .A(net221760), .Y(net264884) );
  CLKINVX1 U29239 ( .A(net221954), .Y(net221760) );
  INVX3 U29240 ( .A(n33900), .Y(n51411) );
  CLKINVX1 U29241 ( .A(net218150), .Y(net218054) );
  CLKBUFX3 U29242 ( .A(net218628), .Y(n40143) );
  CLKBUFX3 U29243 ( .A(net218310), .Y(net262000) );
  CLKBUFX3 U29244 ( .A(net221764), .Y(net264922) );
  CLKINVX1 U29245 ( .A(net221910), .Y(net221764) );
  CLKBUFX3 U29246 ( .A(net218660), .Y(n40129) );
  CLKBUFX3 U29247 ( .A(net218340), .Y(net262285) );
  INVX3 U29248 ( .A(n33892), .Y(n51410) );
  CLKBUFX3 U29249 ( .A(net217088), .Y(n40326) );
  CLKINVX1 U29250 ( .A(n40314), .Y(net217088) );
  CLKBUFX3 U29251 ( .A(net221820), .Y(net265454) );
  CLKBUFX3 U29252 ( .A(net218312), .Y(net262019) );
  CLKINVX1 U29253 ( .A(n43023), .Y(n42860) );
  CLKBUFX3 U29254 ( .A(net218404), .Y(net262893) );
  INVX3 U29255 ( .A(n34012), .Y(n51425) );
  CLKBUFX3 U29256 ( .A(net218710), .Y(n40110) );
  CLKINVX1 U29257 ( .A(n43021), .Y(n42810) );
  INVX3 U29258 ( .A(n33876), .Y(n51408) );
  CLKINVX1 U29259 ( .A(net218150), .Y(net218052) );
  CLKBUFX3 U29260 ( .A(net217086), .Y(n40327) );
  CLKINVX1 U29261 ( .A(n40314), .Y(net217086) );
  CLKBUFX3 U29262 ( .A(net221818), .Y(net265435) );
  CLKBUFX3 U29263 ( .A(net218632), .Y(n40142) );
  CLKBUFX3 U29264 ( .A(net218314), .Y(net262038) );
  INVX3 U29265 ( .A(n33828), .Y(n51402) );
  CLKINVX1 U29266 ( .A(net218150), .Y(net218046) );
  CLKBUFX3 U29267 ( .A(net217082), .Y(n40329) );
  CLKINVX1 U29268 ( .A(n40314), .Y(net217082) );
  CLKBUFX3 U29269 ( .A(net221814), .Y(net265397) );
  INVX3 U29270 ( .A(n33780), .Y(n51396) );
  CLKINVX1 U29271 ( .A(net218150), .Y(net218042) );
  CLKBUFX3 U29272 ( .A(net217078), .Y(n40331) );
  CLKINVX1 U29273 ( .A(n40314), .Y(net217078) );
  INVX3 U29274 ( .A(n33772), .Y(n51395) );
  CLKINVX1 U29275 ( .A(net218150), .Y(net218040) );
  CLKBUFX3 U29276 ( .A(net217076), .Y(n40332) );
  CLKINVX1 U29277 ( .A(n40314), .Y(net217076) );
  CLKBUFX3 U29278 ( .A(net221810), .Y(net265359) );
  CLKBUFX3 U29279 ( .A(net218612), .Y(n40151) );
  CLKBUFX3 U29280 ( .A(net218296), .Y(net261867) );
  CLKINVX1 U29281 ( .A(n43022), .Y(n42845) );
  INVX3 U29282 ( .A(n33748), .Y(n51392) );
  CLKBUFX3 U29283 ( .A(net217074), .Y(n40333) );
  CLKINVX1 U29284 ( .A(n40314), .Y(net217074) );
  CLKBUFX3 U29285 ( .A(net218038), .Y(n40233) );
  CLKBUFX3 U29286 ( .A(net221808), .Y(net265340) );
  CLKBUFX3 U29287 ( .A(net218616), .Y(n40149) );
  CLKBUFX3 U29288 ( .A(net218300), .Y(net261905) );
  INVX3 U29289 ( .A(n33644), .Y(n51379) );
  INVX3 U29290 ( .A(n33660), .Y(n51381) );
  CLKBUFX3 U29291 ( .A(net217066), .Y(n40337) );
  CLKINVX1 U29292 ( .A(n40314), .Y(net217066) );
  CLKBUFX3 U29293 ( .A(net217986), .Y(n40258) );
  CLKINVX1 U29294 ( .A(net218146), .Y(net217986) );
  CLKBUFX3 U29295 ( .A(net221766), .Y(net264941) );
  CLKINVX1 U29296 ( .A(net221908), .Y(net221766) );
  CLKBUFX3 U29297 ( .A(net218658), .Y(n40130) );
  CLKBUFX3 U29298 ( .A(net218338), .Y(net262266) );
  INVX3 U29299 ( .A(n34100), .Y(n51436) );
  INVX3 U29300 ( .A(n34092), .Y(n51435) );
  CLKBUFX3 U29301 ( .A(net217106), .Y(n40318) );
  CLKINVX1 U29302 ( .A(n40313), .Y(net217106) );
  CLKBUFX3 U29303 ( .A(net218030), .Y(n40236) );
  CLKINVX1 U29304 ( .A(net218148), .Y(net218030) );
  CLKBUFX3 U29305 ( .A(net221802), .Y(net265283) );
  CLKBUFX3 U29306 ( .A(net218732), .Y(n40102) );
  CLKBUFX3 U29307 ( .A(net218402), .Y(net262874) );
  CLKINVX1 U29308 ( .A(net218156), .Y(net218130) );
  INVX3 U29309 ( .A(n34120), .Y(n49513) );
  CLKINVX1 U29310 ( .A(net218150), .Y(net218038) );
  CLKBUFX3 U29311 ( .A(net221804), .Y(net265302) );
  CLKBUFX3 U29312 ( .A(net218730), .Y(n40103) );
  CLKBUFX3 U29313 ( .A(net218180), .Y(n40171) );
  CLKBUFX3 U29314 ( .A(net217152), .Y(n40298) );
  CLKBUFX3 U29315 ( .A(net218698), .Y(n40115) );
  CLKBUFX3 U29316 ( .A(net218372), .Y(net262589) );
  CLKBUFX3 U29317 ( .A(n34395), .Y(n42066) );
  CLKBUFX3 U29318 ( .A(n34403), .Y(n42065) );
  CLKBUFX3 U29319 ( .A(net218364), .Y(net262513) );
  CLKBUFX3 U29320 ( .A(net221918), .Y(net266381) );
  CLKBUFX3 U29321 ( .A(net217142), .Y(n40303) );
  CLKBUFX3 U29322 ( .A(net218366), .Y(net262532) );
  CLKBUFX3 U29323 ( .A(net217950), .Y(n40272) );
  CLKINVX1 U29324 ( .A(net218154), .Y(net217950) );
  CLKINVX1 U29325 ( .A(net266151), .Y(net221732) );
  CLKBUFX3 U29326 ( .A(net217956), .Y(n40269) );
  CLKBUFX3 U29327 ( .A(net217188), .Y(n40281) );
  BUFX4 U29328 ( .A(net221856), .Y(net265796) );
  CLKINVX1 U29329 ( .A(net266218), .Y(net221856) );
  CLKBUFX3 U29330 ( .A(net218792), .Y(n40074) );
  CLKBUFX3 U29331 ( .A(net217184), .Y(n40283) );
  CLKBUFX3 U29332 ( .A(net217182), .Y(n40284) );
  CLKINVX1 U29333 ( .A(net218156), .Y(net218116) );
  CLKBUFX3 U29334 ( .A(net218778), .Y(n40080) );
  CLKINVX1 U29335 ( .A(net218156), .Y(net218114) );
  CLKBUFX3 U29336 ( .A(net218398), .Y(net262836) );
  CLKINVX1 U29337 ( .A(net266151), .Y(net221726) );
  CLKBUFX3 U29338 ( .A(net217196), .Y(n40279) );
  CLKBUFX3 U29339 ( .A(net218752), .Y(n40093) );
  CLKBUFX3 U29340 ( .A(net218368), .Y(net262551) );
  CLKBUFX3 U29341 ( .A(net218728), .Y(n40104) );
  CLKBUFX3 U29342 ( .A(net218400), .Y(net262855) );
  CLKBUFX3 U29343 ( .A(net218064), .Y(n40220) );
  CLKINVX1 U29344 ( .A(net218152), .Y(net218064) );
  CLKBUFX3 U29345 ( .A(net218004), .Y(n40249) );
  CLKINVX1 U29346 ( .A(net218146), .Y(net218004) );
  CLKBUFX3 U29347 ( .A(net221780), .Y(net265074) );
  CLKINVX1 U29348 ( .A(net221914), .Y(net221780) );
  CLKINVX1 U29349 ( .A(n43018), .Y(n42769) );
  CLKBUFX3 U29350 ( .A(net218480), .Y(net263615) );
  CLKINVX1 U29351 ( .A(n40315), .Y(net217044) );
  INVX3 U29352 ( .A(n33388), .Y(n51347) );
  INVX3 U29353 ( .A(n33380), .Y(n51346) );
  CLKBUFX3 U29354 ( .A(net218482), .Y(net263634) );
  CLKBUFX3 U29355 ( .A(net218002), .Y(n40250) );
  CLKINVX1 U29356 ( .A(net218146), .Y(net218002) );
  CLKBUFX3 U29357 ( .A(net221778), .Y(net265055) );
  CLKINVX1 U29358 ( .A(net221954), .Y(net221778) );
  INVX3 U29359 ( .A(n34004), .Y(n51424) );
  CLKBUFX3 U29360 ( .A(net217098), .Y(n40322) );
  CLKBUFX3 U29361 ( .A(net218022), .Y(n40240) );
  CLKINVX1 U29362 ( .A(net218148), .Y(net218022) );
  CLKBUFX3 U29363 ( .A(net218384), .Y(net262703) );
  INVX3 U29364 ( .A(n33996), .Y(n51423) );
  CLKBUFX3 U29365 ( .A(net217096), .Y(n40323) );
  CLKBUFX3 U29366 ( .A(net218020), .Y(n40241) );
  CLKINVX1 U29367 ( .A(net218148), .Y(net218020) );
  CLKINVX1 U29368 ( .A(net221966), .Y(net221794) );
  CLKBUFX3 U29369 ( .A(net218712), .Y(n40109) );
  CLKBUFX3 U29370 ( .A(net218386), .Y(net262722) );
  CLKBUFX3 U29371 ( .A(net218490), .Y(net263710) );
  CLKINVX1 U29372 ( .A(net218146), .Y(net217994) );
  CLKBUFX3 U29373 ( .A(net217998), .Y(n40252) );
  CLKINVX1 U29374 ( .A(net218146), .Y(net217998) );
  CLKBUFX3 U29375 ( .A(net218486), .Y(net263672) );
  CLKINVX1 U29376 ( .A(n40315), .Y(net217042) );
  CLKBUFX3 U29377 ( .A(net218484), .Y(net263653) );
  CLKBUFX3 U29378 ( .A(net218000), .Y(n40251) );
  CLKINVX1 U29379 ( .A(net218146), .Y(net218000) );
  CLKINVX1 U29380 ( .A(net221966), .Y(net221776) );
  CLKINVX1 U29381 ( .A(n43019), .Y(n42775) );
  CLKBUFX3 U29382 ( .A(net221774), .Y(net265017) );
  CLKINVX1 U29383 ( .A(net221916), .Y(net221774) );
  CLKINVX1 U29384 ( .A(n40315), .Y(net217038) );
  CLKBUFX3 U29385 ( .A(net217996), .Y(n40253) );
  CLKINVX1 U29386 ( .A(net218146), .Y(net217996) );
  CLKBUFX3 U29387 ( .A(net221772), .Y(net264998) );
  CLKINVX1 U29388 ( .A(net221912), .Y(net221772) );
  CLKBUFX3 U29389 ( .A(net218488), .Y(net263691) );
  CLKINVX1 U29390 ( .A(n43019), .Y(n42779) );
  CLKBUFX3 U29391 ( .A(net218850), .Y(n40046) );
  CLKBUFX3 U29392 ( .A(n34367), .Y(n41812) );
  CLKBUFX3 U29393 ( .A(n34359), .Y(n41813) );
  CLKBUFX3 U29394 ( .A(net218174), .Y(n40174) );
  CLKBUFX3 U29395 ( .A(n34391), .Y(n41809) );
  CLKBUFX3 U29396 ( .A(net221920), .Y(net266402) );
  CLKBUFX3 U29397 ( .A(net217144), .Y(n40302) );
  CLKBUFX3 U29398 ( .A(n34375), .Y(n41811) );
  CLKBUFX3 U29399 ( .A(n34383), .Y(n41810) );
  CLKBUFX3 U29400 ( .A(net218694), .Y(n40117) );
  CLKBUFX3 U29401 ( .A(net218370), .Y(net262570) );
  CLKBUFX3 U29402 ( .A(net217022), .Y(n40357) );
  CLKINVX1 U29403 ( .A(n40316), .Y(net217022) );
  CLKBUFX3 U29404 ( .A(net218106), .Y(n40199) );
  CLKINVX1 U29405 ( .A(net218154), .Y(net218106) );
  CLKBUFX3 U29406 ( .A(net218852), .Y(n40045) );
  CLKBUFX3 U29407 ( .A(net218508), .Y(net263881) );
  CLKBUFX3 U29408 ( .A(net221864), .Y(net265872) );
  CLKINVX1 U29409 ( .A(net266235), .Y(net221864) );
  CLKBUFX3 U29410 ( .A(net218510), .Y(net263900) );
  CLKBUFX3 U29411 ( .A(net217020), .Y(n40358) );
  CLKBUFX3 U29412 ( .A(net218104), .Y(n40200) );
  CLKINVX1 U29413 ( .A(net218154), .Y(net218104) );
  CLKBUFX3 U29414 ( .A(net218854), .Y(n40044) );
  CLKBUFX3 U29415 ( .A(net218512), .Y(net263919) );
  CLKINVX1 U29416 ( .A(n40316), .Y(net217026) );
  CLKBUFX3 U29417 ( .A(net221866), .Y(net265891) );
  CLKINVX1 U29418 ( .A(net266235), .Y(net221866) );
  CLKBUFX3 U29419 ( .A(net218518), .Y(net263976) );
  CLKBUFX3 U29420 ( .A(net218520), .Y(net263995) );
  CLKBUFX3 U29421 ( .A(net217018), .Y(n40359) );
  CLKBUFX3 U29422 ( .A(net218102), .Y(n40201) );
  CLKINVX1 U29423 ( .A(net218154), .Y(net218102) );
  CLKBUFX3 U29424 ( .A(net221862), .Y(net265853) );
  CLKINVX1 U29425 ( .A(net266218), .Y(net221862) );
  CLKBUFX3 U29426 ( .A(net218856), .Y(n40043) );
  CLKBUFX3 U29427 ( .A(net218100), .Y(n40202) );
  CLKINVX1 U29428 ( .A(net218154), .Y(net218100) );
  CLKBUFX3 U29429 ( .A(net221860), .Y(net265834) );
  CLKINVX1 U29430 ( .A(net266218), .Y(net221860) );
  CLKBUFX3 U29431 ( .A(net217016), .Y(n40360) );
  CLKBUFX3 U29432 ( .A(net218098), .Y(n40203) );
  CLKINVX1 U29433 ( .A(net218154), .Y(net218098) );
  CLKBUFX3 U29434 ( .A(net221858), .Y(net265815) );
  CLKINVX1 U29435 ( .A(net266218), .Y(net221858) );
  CLKBUFX3 U29436 ( .A(net218860), .Y(n40042) );
  CLKBUFX3 U29437 ( .A(net218516), .Y(net263957) );
  CLKBUFX3 U29438 ( .A(net217012), .Y(n40361) );
  CLKBUFX3 U29439 ( .A(net218834), .Y(n40054) );
  CLKBUFX3 U29440 ( .A(net218494), .Y(net263748) );
  CLKBUFX3 U29441 ( .A(net218132), .Y(n40186) );
  CLKBUFX3 U29442 ( .A(net221886), .Y(net266081) );
  CLKINVX1 U29443 ( .A(net266235), .Y(net221886) );
  CLKBUFX3 U29444 ( .A(net218840), .Y(n40051) );
  CLKBUFX3 U29445 ( .A(net217008), .Y(n40363) );
  CLKINVX1 U29446 ( .A(n40316), .Y(net217008) );
  CLKBUFX3 U29447 ( .A(net218136), .Y(n40185) );
  CLKINVX1 U29448 ( .A(n40182), .Y(net218136) );
  CLKBUFX3 U29449 ( .A(net221890), .Y(net266119) );
  CLKINVX1 U29450 ( .A(net266235), .Y(net221890) );
  CLKBUFX3 U29451 ( .A(net217010), .Y(n40362) );
  CLKBUFX3 U29452 ( .A(net218110), .Y(n40197) );
  CLKBUFX3 U29453 ( .A(net221888), .Y(net266100) );
  CLKINVX1 U29454 ( .A(net266235), .Y(net221888) );
  CLKBUFX3 U29455 ( .A(net218838), .Y(n40052) );
  CLKBUFX3 U29456 ( .A(net218496), .Y(net263767) );
  INVX12 U29457 ( .A(n41196), .Y(codeword[3]) );
  OAI21XL U29458 ( .A0(n40516), .A1(n40633), .B0(n40754), .Y(n40462) );
  AOI21X1 U29459 ( .A0(n40758), .A1(n40752), .B0(n36932), .Y(n40464) );
  NAND4BX1 U29460 ( .AN(n39475), .B(net208565), .C(n39476), .D(n39477), .Y(
        n34513) );
  NOR3BXL U29461 ( .AN(n39696), .B(net218294), .C(n39697), .Y(n39475) );
  NAND3BX1 U29462 ( .AN(net218610), .B(n40000), .C(n40020), .Y(n39477) );
  AOI211X1 U29463 ( .A0(n39875), .A1(n40004), .B0(n39774), .C0(n37526), .Y(
        n39476) );
  INVX20 U29464 ( .A(n37597), .Y(n37598) );
  NOR4X1 U29465 ( .A(n44980), .B(n44979), .C(n44978), .D(n44977), .Y(n44981)
         );
  XOR2X1 U29466 ( .A(n42069), .B(n36889), .Y(n44978) );
  OAI31X1 U29467 ( .A0(n11061), .A1(net209203), .A2(net151644), .B0(n11064),
        .Y(n11059) );
  INVXL U29468 ( .A(n42638), .Y(n41388) );
  CLKBUFX3 U29469 ( .A(n34458), .Y(n42499) );
  CLKBUFX3 U29470 ( .A(net217048), .Y(n40346) );
  CLKBUFX3 U29471 ( .A(net217054), .Y(n40343) );
  CLKBUFX3 U29472 ( .A(net217058), .Y(n40341) );
  CLKBUFX3 U29473 ( .A(net218128), .Y(n40188) );
  CLKBUFX3 U29474 ( .A(net218126), .Y(n40189) );
  CLKBUFX3 U29475 ( .A(net218108), .Y(n40198) );
  CLKBUFX3 U29476 ( .A(net218256), .Y(net218150) );
  CLKINVX1 U29477 ( .A(net218150), .Y(net218034) );
  CLKBUFX3 U29478 ( .A(net218034), .Y(n40235) );
  CLKINVX1 U29479 ( .A(net218156), .Y(net218124) );
  BUFX4 U29480 ( .A(net221776), .Y(net265036) );
  BUFX4 U29481 ( .A(net221794), .Y(net265207) );
  BUFX4 U29482 ( .A(net221768), .Y(net264960) );
  CLKBUFX3 U29483 ( .A(net217038), .Y(n40350) );
  CLKBUFX3 U29484 ( .A(net217042), .Y(n40349) );
  CLKBUFX3 U29485 ( .A(net217044), .Y(n40348) );
  CLKBUFX3 U29486 ( .A(net217120), .Y(n40313) );
  CLKINVX1 U29487 ( .A(n40313), .Y(net217096) );
  CLKINVX1 U29488 ( .A(n40313), .Y(net217098) );
  CLKINVX1 U29489 ( .A(n40313), .Y(net217102) );
  CLKBUFX3 U29490 ( .A(net218666), .Y(n40127) );
  CLKBUFX3 U29491 ( .A(net218864), .Y(n40040) );
  CLKBUFX3 U29492 ( .A(net218830), .Y(n40056) );
  CLKBUFX3 U29493 ( .A(net218836), .Y(n40053) );
  CLKBUFX3 U29494 ( .A(net218114), .Y(n40195) );
  CLKBUFX3 U29495 ( .A(net218116), .Y(n40194) );
  CLKBUFX3 U29496 ( .A(net218112), .Y(n40196) );
  CLKBUFX3 U29497 ( .A(net218158), .Y(n40182) );
  CLKINVX1 U29498 ( .A(net218156), .Y(net218110) );
  CLKINVX1 U29499 ( .A(net218156), .Y(net218132) );
  CLKBUFX3 U29500 ( .A(n42474), .Y(n42472) );
  CLKBUFX6 U29501 ( .A(net221788), .Y(net265150) );
  BUFX4 U29502 ( .A(net218440), .Y(net263235) );
  BUFX4 U29503 ( .A(net218446), .Y(net263292) );
  CLKBUFX3 U29504 ( .A(net218438), .Y(net263216) );
  CLKBUFX6 U29505 ( .A(net216968), .Y(n40382) );
  CLKBUFX3 U29506 ( .A(net216966), .Y(n40383) );
  CLKINVX1 U29507 ( .A(net217242), .Y(net216968) );
  CLKBUFX3 U29508 ( .A(net218774), .Y(n40082) );
  CLKBUFX3 U29509 ( .A(net218794), .Y(n40073) );
  CLKBUFX3 U29510 ( .A(net218776), .Y(n40081) );
  BUFX4 U29511 ( .A(net221762), .Y(net264903) );
  BUFX4 U29512 ( .A(net221756), .Y(net264846) );
  CLKBUFX3 U29513 ( .A(net218672), .Y(n40124) );
  CLKBUFX3 U29514 ( .A(net218654), .Y(n40132) );
  CLKBUFX3 U29515 ( .A(net218656), .Y(n40131) );
  BUFX4 U29516 ( .A(net218796), .Y(n40072) );
  CLKBUFX3 U29517 ( .A(net218254), .Y(net218154) );
  CLKBUFX3 U29518 ( .A(net218168), .Y(n40177) );
  BUFX4 U29519 ( .A(n42468), .Y(n42465) );
  INVX3 U29520 ( .A(net219346), .Y(net219314) );
  INVX3 U29521 ( .A(net219472), .Y(net219466) );
  INVX6 U29522 ( .A(net219478), .Y(net219450) );
  BUFX4 U29523 ( .A(n42650), .Y(n42663) );
  INVX4 U29524 ( .A(n42716), .Y(n42706) );
  INVX4 U29525 ( .A(n42679), .Y(n42670) );
  BUFX4 U29526 ( .A(net216978), .Y(n40377) );
  CLKBUFX3 U29527 ( .A(net217034), .Y(n40351) );
  CLKBUFX3 U29528 ( .A(net217046), .Y(n40347) );
  CLKBUFX3 U29529 ( .A(net217114), .Y(n40316) );
  CLKINVX1 U29530 ( .A(n40316), .Y(net217020) );
  CLKINVX1 U29531 ( .A(n40316), .Y(net217016) );
  CLKINVX1 U29532 ( .A(n40316), .Y(net217018) );
  BUFX4 U29533 ( .A(net218824), .Y(n40058) );
  CLKBUFX3 U29534 ( .A(net218754), .Y(n40092) );
  CLKBUFX3 U29535 ( .A(net218800), .Y(n40070) );
  CLKBUFX3 U29536 ( .A(net218842), .Y(n40050) );
  CLKBUFX3 U29537 ( .A(net218844), .Y(n40049) );
  INVX4 U29538 ( .A(n42714), .Y(n42705) );
  CLKBUFX3 U29539 ( .A(n42511), .Y(n42527) );
  CLKBUFX3 U29540 ( .A(net217004), .Y(n40364) );
  CLKBUFX3 U29541 ( .A(net216984), .Y(n40374) );
  CLKBUFX3 U29542 ( .A(net216998), .Y(n40367) );
  CLKBUFX3 U29543 ( .A(net217112), .Y(n40317) );
  CLKINVX1 U29544 ( .A(n40317), .Y(net217000) );
  CLKBUFX3 U29545 ( .A(net217000), .Y(n40366) );
  CLKINVX1 U29546 ( .A(n40317), .Y(net216982) );
  CLKBUFX3 U29547 ( .A(net218770), .Y(n40084) );
  CLKBUFX3 U29548 ( .A(net218768), .Y(n40085) );
  CLKBUFX3 U29549 ( .A(net218756), .Y(n40091) );
  CLKBUFX3 U29550 ( .A(net218018), .Y(n40242) );
  CLKBUFX3 U29551 ( .A(net218048), .Y(n40228) );
  CLKBUFX3 U29552 ( .A(net218052), .Y(n40226) );
  CLKBUFX3 U29553 ( .A(net218122), .Y(n40191) );
  CLKINVX1 U29554 ( .A(net266201), .Y(net221802) );
  CLKINVX1 U29555 ( .A(net266201), .Y(net221810) );
  CLKINVX1 U29556 ( .A(net266201), .Y(net221804) );
  CLKBUFX3 U29557 ( .A(n42599), .Y(n42598) );
  INVX4 U29558 ( .A(n42621), .Y(n42618) );
  CLKBUFX6 U29559 ( .A(net217174), .Y(n40287) );
  BUFX4 U29560 ( .A(net218804), .Y(n40068) );
  CLKBUFX3 U29561 ( .A(net218828), .Y(n40057) );
  CLKBUFX3 U29562 ( .A(net217994), .Y(n40254) );
  CLKBUFX3 U29563 ( .A(net218054), .Y(n40225) );
  CLKBUFX3 U29564 ( .A(net218060), .Y(n40222) );
  CLKBUFX3 U29565 ( .A(net218046), .Y(n40229) );
  CLKBUFX3 U29566 ( .A(n42476), .Y(n42468) );
  BUFX4 U29567 ( .A(net221790), .Y(net265169) );
  BUFX4 U29568 ( .A(net221798), .Y(net265245) );
  INVX3 U29569 ( .A(n42556), .Y(n42549) );
  INVX4 U29570 ( .A(n42713), .Y(n42704) );
  INVX3 U29571 ( .A(n42585), .Y(n42575) );
  INVX6 U29572 ( .A(n42510), .Y(n42500) );
  INVX6 U29573 ( .A(n42686), .Y(n42681) );
  CLKBUFX3 U29574 ( .A(n34452), .Y(n42557) );
  BUFX4 U29575 ( .A(net217136), .Y(n40306) );
  BUFX4 U29576 ( .A(net217170), .Y(n40289) );
  CLKBUFX3 U29577 ( .A(net218862), .Y(n40041) );
  CLKBUFX3 U29578 ( .A(net218822), .Y(n40059) );
  CLKBUFX3 U29579 ( .A(net218820), .Y(n40060) );
  CLKINVX1 U29580 ( .A(n40183), .Y(net217968) );
  CLKBUFX3 U29581 ( .A(net218006), .Y(n40248) );
  CLKBUFX3 U29582 ( .A(net218016), .Y(n40243) );
  CLKBUFX3 U29583 ( .A(net218040), .Y(n40232) );
  BUFX4 U29584 ( .A(net221828), .Y(net265530) );
  BUFX4 U29585 ( .A(net221826), .Y(net265511) );
  BUFX4 U29586 ( .A(net221816), .Y(net265416) );
  BUFX4 U29587 ( .A(net221824), .Y(net265492) );
  CLKBUFX3 U29588 ( .A(n42703), .Y(n41384) );
  INVX4 U29589 ( .A(n42677), .Y(n42675) );
  INVX6 U29590 ( .A(n42713), .Y(n42711) );
  INVX3 U29591 ( .A(n42714), .Y(n41642) );
  INVX6 U29592 ( .A(n42585), .Y(n42579) );
  CLKINVX1 U29593 ( .A(n42688), .Y(n42680) );
  CLKINVX1 U29594 ( .A(net217224), .Y(net216970) );
  BUFX4 U29595 ( .A(net216970), .Y(n40381) );
  CLKBUFX3 U29596 ( .A(net218762), .Y(n40088) );
  CLKBUFX3 U29597 ( .A(net218848), .Y(n40047) );
  CLKBUFX3 U29598 ( .A(net218764), .Y(n40087) );
  CLKINVX1 U29599 ( .A(n40183), .Y(net217962) );
  CLKBUFX3 U29600 ( .A(net218050), .Y(n40227) );
  CLKBUFX3 U29601 ( .A(net218042), .Y(n40231) );
  CLKBUFX3 U29602 ( .A(net218044), .Y(n40230) );
  INVX4 U29603 ( .A(n42572), .Y(n42560) );
  CLKBUFX3 U29604 ( .A(n34474), .Y(n42458) );
  CLKBUFX3 U29605 ( .A(net221902), .Y(net266218) );
  CLKINVX1 U29606 ( .A(net266218), .Y(net221854) );
  CLKINVX1 U29607 ( .A(net266201), .Y(net221800) );
  CLKINVX1 U29608 ( .A(net266201), .Y(net221806) );
  CLKINVX1 U29609 ( .A(net266201), .Y(net221830) );
  CLKBUFX3 U29610 ( .A(n42598), .Y(n42595) );
  INVX3 U29611 ( .A(net219492), .Y(net219460) );
  BUFX4 U29612 ( .A(net217118), .Y(n40314) );
  CLKBUFX3 U29613 ( .A(net218668), .Y(n40126) );
  CLKBUFX3 U29614 ( .A(net218646), .Y(n40136) );
  CLKBUFX3 U29615 ( .A(net218644), .Y(n40137) );
  CLKBUFX3 U29616 ( .A(net218810), .Y(n40065) );
  CLKBUFX3 U29617 ( .A(net217938), .Y(n40275) );
  INVX6 U29618 ( .A(n42510), .Y(n42505) );
  BUFX4 U29619 ( .A(net221850), .Y(net265739) );
  BUFX4 U29620 ( .A(net221854), .Y(net265777) );
  BUFX4 U29621 ( .A(net221844), .Y(net265682) );
  INVX4 U29622 ( .A(n42645), .Y(n42641) );
  INVX3 U29623 ( .A(n36927), .Y(n42550) );
  INVX4 U29624 ( .A(n41308), .Y(n41309) );
  CLKBUFX3 U29625 ( .A(n42531), .Y(n42516) );
  CLKBUFX3 U29626 ( .A(net218634), .Y(n40141) );
  CLKBUFX3 U29627 ( .A(net218652), .Y(n40133) );
  CLKBUFX3 U29628 ( .A(net218816), .Y(n40062) );
  CLKBUFX3 U29629 ( .A(net218802), .Y(n40069) );
  CLKBUFX3 U29630 ( .A(net218812), .Y(n40064) );
  CLKINVX1 U29631 ( .A(n40177), .Y(net217930) );
  CLKBUFX3 U29632 ( .A(net218014), .Y(n40244) );
  CLKBUFX3 U29633 ( .A(net218010), .Y(n40246) );
  CLKBUFX3 U29634 ( .A(net218036), .Y(n40234) );
  INVX6 U29635 ( .A(n42570), .Y(n42569) );
  CLKBUFX3 U29636 ( .A(net221904), .Y(net266235) );
  CLKINVX1 U29637 ( .A(net266235), .Y(net221880) );
  CLKINVX1 U29638 ( .A(net266218), .Y(net221848) );
  CLKINVX1 U29639 ( .A(net266218), .Y(net221852) );
  CLKINVX1 U29640 ( .A(net266218), .Y(net221834) );
  INVX6 U29641 ( .A(n41289), .Y(n41296) );
  AND2X2 U29642 ( .A(n36928), .B(n41736), .Y(n41789) );
  INVX3 U29643 ( .A(n34465), .Y(n41315) );
  INVX6 U29644 ( .A(n41315), .Y(n41318) );
  INVX4 U29645 ( .A(n41315), .Y(n41317) );
  INVX4 U29646 ( .A(n41326), .Y(n41328) );
  INVX4 U29647 ( .A(n42727), .Y(n42721) );
  CLKINVX1 U29648 ( .A(n42727), .Y(n42722) );
  CLKBUFX3 U29649 ( .A(net218760), .Y(n40089) );
  CLKBUFX3 U29650 ( .A(net218748), .Y(n40095) );
  BUFX4 U29651 ( .A(net218766), .Y(n40086) );
  CLKBUFX3 U29652 ( .A(net218808), .Y(n40066) );
  CLKBUFX3 U29653 ( .A(net218818), .Y(n40061) );
  CLKBUFX3 U29654 ( .A(net218806), .Y(n40067) );
  CLKBUFX6 U29655 ( .A(net217218), .Y(net217178) );
  CLKINVX1 U29656 ( .A(n40178), .Y(net217936) );
  CLKBUFX3 U29657 ( .A(net217946), .Y(n40273) );
  CLKBUFX3 U29658 ( .A(net217934), .Y(n40276) );
  INVX4 U29659 ( .A(n42573), .Y(n42558) );
  CLKBUFX3 U29660 ( .A(net218452), .Y(net263349) );
  CLKBUFX3 U29661 ( .A(net218462), .Y(net263444) );
  CLKBUFX3 U29662 ( .A(net221894), .Y(net266151) );
  INVX6 U29663 ( .A(net221962), .Y(net221892) );
  CLKBUFX6 U29664 ( .A(n34453), .Y(n41321) );
  NAND2BX2 U29665 ( .AN(n_cell_301249_net267385), .B(net216337), .Y(
        n_cell_303546_net275987) );
  INVX3 U29666 ( .A(n42713), .Y(n42712) );
  INVX6 U29667 ( .A(n41315), .Y(n41316) );
  INVX6 U29668 ( .A(n41298), .Y(n41305) );
  INVX6 U29669 ( .A(n41326), .Y(n41331) );
  CLKBUFX3 U29670 ( .A(n42649), .Y(n42666) );
  CLKBUFX3 U29671 ( .A(net218786), .Y(n40077) );
  CLKBUFX3 U29672 ( .A(net218780), .Y(n40079) );
  CLKBUFX3 U29673 ( .A(net218846), .Y(n40048) );
  CLKBUFX3 U29674 ( .A(net218814), .Y(n40063) );
  INVX3 U29675 ( .A(net219484), .Y(net258207) );
  CLKBUFX3 U29676 ( .A(net218144), .Y(n40183) );
  CLKBUFX3 U29677 ( .A(net218120), .Y(n40192) );
  INVX4 U29678 ( .A(n42571), .Y(n42568) );
  CLKBUFX3 U29679 ( .A(n42480), .Y(n42479) );
  CLKBUFX3 U29680 ( .A(net221726), .Y(net264607) );
  CLKBUFX3 U29681 ( .A(net221722), .Y(net264577) );
  CLKBUFX3 U29682 ( .A(net221732), .Y(net264652) );
  AND2X2 U29683 ( .A(n41736), .B(n41199), .Y(n41790) );
  NAND2BX2 U29684 ( .AN(n_cell_301249_net267141), .B(net211788), .Y(
        n_cell_303546_net275956) );
  CLKBUFX6 U29685 ( .A(n36873), .Y(n41325) );
  NAND2BX2 U29686 ( .AN(n_cell_301249_net267117), .B(net213552), .Y(
        n_cell_303546_net275923) );
  NAND2BX2 U29687 ( .AN(n40779), .B(net212826), .Y(n10904) );
  NAND2X1 U29688 ( .A(n37013), .B(net216166), .Y(n11917) );
  NAND2X1 U29689 ( .A(n37122), .B(net216274), .Y(n11932) );
  INVX3 U29690 ( .A(n42545), .Y(n42538) );
  CLKINVX1 U29691 ( .A(n34436), .Y(n42716) );
  NAND2BX1 U29692 ( .AN(n_cell_301249_net267628), .B(net213487), .Y(n12392) );
  NAND2BX1 U29693 ( .AN(n40434), .B(n_cell_301249_net267903), .Y(n11568) );
  INVX3 U29694 ( .A(n41315), .Y(n41314) );
  INVX6 U29695 ( .A(n41315), .Y(n41311) );
  INVX6 U29696 ( .A(n41298), .Y(n41303) );
  INVX6 U29697 ( .A(n41326), .Y(n41327) );
  INVX3 U29698 ( .A(n41289), .Y(n41290) );
  INVX6 U29699 ( .A(n41289), .Y(n41291) );
  INVX4 U29700 ( .A(n41289), .Y(n41292) );
  CLKBUFX3 U29701 ( .A(net218758), .Y(n40090) );
  CLKBUFX3 U29702 ( .A(net218798), .Y(n40071) );
  NOR2X1 U29703 ( .A(n37239), .B(net171535), .Y(n36926) );
  NAND3X2 U29704 ( .A(net216291), .B(net216290), .C(n_cell_301249_net267447),
        .Y(n40411) );
  CLKINVX1 U29705 ( .A(net218232), .Y(net217940) );
  CLKBUFX3 U29706 ( .A(net217940), .Y(n40274) );
  CLKBUFX3 U29707 ( .A(net217960), .Y(n40268) );
  CLKBUFX3 U29708 ( .A(net217932), .Y(n40277) );
  NOR2X1 U29709 ( .A(net260384), .B(net171380), .Y(n36928) );
  INVX3 U29710 ( .A(n41648), .Y(n41287) );
  INVX4 U29711 ( .A(n42585), .Y(n42577) );
  NOR2X1 U29712 ( .A(net209402), .B(n40457), .Y(n36929) );
  NAND2BX1 U29713 ( .AN(n_cell_301249_net267846), .B(net212073), .Y(n39342) );
  AO21X1 U29714 ( .A0(n39548), .A1(n36929), .B0(n40755), .Y(n36932) );
  BUFX4 U29715 ( .A(n42472), .Y(n42466) );
  NAND4X1 U29716 ( .A(n43275), .B(n43274), .C(n43273), .D(n43272), .Y(
        net214730) );
  NAND2BX1 U29717 ( .AN(n_cell_301249_net267135), .B(net211783), .Y(n11291) );
  CLKINVX1 U29718 ( .A(net266151), .Y(net221720) );
  CLKBUFX3 U29719 ( .A(net221736), .Y(net264682) );
  CLKINVX1 U29720 ( .A(net266151), .Y(net221736) );
  INVX3 U29721 ( .A(n11282), .Y(n_cell_303546_net277530) );
  AND4X1 U29722 ( .A(n45054), .B(n45053), .C(n45052), .D(n45051), .Y(n36934)
         );
  NAND2X2 U29723 ( .A(n41736), .B(n9747), .Y(n36935) );
  AND2X2 U29724 ( .A(n47982), .B(n47980), .Y(n36936) );
  OR4X1 U29725 ( .A(n27520), .B(n27521), .C(n27522), .D(n27523), .Y(n36937) );
  OR4X1 U29726 ( .A(n27309), .B(n27310), .C(n27311), .D(n27312), .Y(n36938) );
  OR4X1 U29727 ( .A(n45327), .B(n45326), .C(n45325), .D(n45324), .Y(n36940) );
  CLKINVX1 U29728 ( .A(net210047), .Y(net171535) );
  NOR4X1 U29729 ( .A(n45089), .B(n45088), .C(n45087), .D(n45086), .Y(n36941)
         );
  CLKINVX1 U29730 ( .A(net209249), .Y(net171486) );
  AND4X1 U29731 ( .A(n46708), .B(n46707), .C(n46706), .D(n46705), .Y(n36942)
         );
  AND4X1 U29732 ( .A(n46808), .B(n46807), .C(n46806), .D(n46805), .Y(n36943)
         );
  AND4X1 U29733 ( .A(n47188), .B(n47187), .C(n47186), .D(n47185), .Y(n36944)
         );
  AND4X1 U29734 ( .A(n47946), .B(n47945), .C(n47944), .D(n47943), .Y(n36945)
         );
  NAND2BX1 U29735 ( .AN(n_cell_301249_net267373), .B(net216283), .Y(n12804) );
  NAND2BX1 U29736 ( .AN(n_cell_301249_net267484), .B(net212038), .Y(n12848) );
  NAND4X1 U29737 ( .A(n45989), .B(n45988), .C(n45987), .D(n45986), .Y(n11034)
         );
  AND4X1 U29738 ( .A(n47247), .B(n47246), .C(n47245), .D(n47244), .Y(n36948)
         );
  NAND4X1 U29739 ( .A(n45822), .B(n45821), .C(n45820), .D(n45819), .Y(n12388)
         );
  XOR2X1 U29740 ( .A(n33770), .B(n42562), .Y(n36949) );
  XOR2X1 U29741 ( .A(n36846), .B(n33986), .Y(n36950) );
  XOR2X1 U29742 ( .A(n36844), .B(n33954), .Y(n36951) );
  OR4X1 U29743 ( .A(n30369), .B(n30370), .C(n30371), .D(n30372), .Y(n36952) );
  OR4X1 U29744 ( .A(n26827), .B(n26828), .C(n26829), .D(n26830), .Y(n36953) );
  OR4X1 U29745 ( .A(n29406), .B(n29407), .C(n29408), .D(n29409), .Y(n36954) );
  OR4X1 U29746 ( .A(n30339), .B(n30340), .C(n30341), .D(n30342), .Y(n36955) );
  OR4X1 U29747 ( .A(n30429), .B(n30430), .C(n30431), .D(n30432), .Y(n36956) );
  OR4X1 U29748 ( .A(n31724), .B(n31725), .C(n31726), .D(n31727), .Y(n36957) );
  OR4X1 U29749 ( .A(n31664), .B(n31665), .C(n31666), .D(n31667), .Y(n36958) );
  OR4X1 U29750 ( .A(n31814), .B(n31815), .C(n31816), .D(n31817), .Y(n36959) );
  OR4X1 U29751 ( .A(n30882), .B(n30883), .C(n30884), .D(n30885), .Y(n36960) );
  OR4X1 U29752 ( .A(n30702), .B(n30703), .C(n30704), .D(n30705), .Y(n36961) );
  OR4X1 U29753 ( .A(n29565), .B(n29566), .C(n29567), .D(n29568), .Y(n36962) );
  OR4X1 U29754 ( .A(n26526), .B(n26527), .C(n26528), .D(n26529), .Y(n36963) );
  OR4X1 U29755 ( .A(n29776), .B(n29777), .C(n29778), .D(n29779), .Y(n36964) );
  OR4X1 U29756 ( .A(n30641), .B(n30642), .C(n30643), .D(n30644), .Y(n36965) );
  OR4X1 U29757 ( .A(n30551), .B(n30552), .C(n30553), .D(n30554), .Y(n36966) );
  OR4X1 U29758 ( .A(n29527), .B(n29528), .C(n29529), .D(n29530), .Y(n36967) );
  OR4X1 U29759 ( .A(n29715), .B(n29716), .C(n29717), .D(n29718), .Y(n36968) );
  OR4X1 U29760 ( .A(n29655), .B(n29656), .C(n29657), .D(n29658), .Y(n36969) );
  OR4X1 U29761 ( .A(n30461), .B(n30462), .C(n30463), .D(n30464), .Y(n36970) );
  OR4X1 U29762 ( .A(n30671), .B(n30672), .C(n30673), .D(n30674), .Y(n36971) );
  OR4X1 U29763 ( .A(n30491), .B(n30492), .C(n30493), .D(n30494), .Y(n36972) );
  OR4X1 U29764 ( .A(n30762), .B(n30763), .C(n30764), .D(n30765), .Y(n36973) );
  OR4X1 U29765 ( .A(n29486), .B(n29485), .C(n29484), .D(n29483), .Y(n36974) );
  OR4X1 U29766 ( .A(n27381), .B(n27380), .C(n27379), .D(n27378), .Y(n36975) );
  OR4X1 U29767 ( .A(n27320), .B(n27319), .C(n27318), .D(n27317), .Y(n36976) );
  OR4X1 U29768 ( .A(n27350), .B(n27349), .C(n27348), .D(n27347), .Y(n36977) );
  OR4X1 U29769 ( .A(n30822), .B(n30823), .C(n30824), .D(n30825), .Y(n36978) );
  OR4X1 U29770 ( .A(n30852), .B(n30853), .C(n30854), .D(n30855), .Y(n36979) );
  OR4X1 U29771 ( .A(n30732), .B(n30733), .C(n30734), .D(n30735), .Y(n36980) );
  OR4X1 U29772 ( .A(n27400), .B(n27401), .C(n27402), .D(n27403), .Y(n36981) );
  OR4X1 U29773 ( .A(n25805), .B(n25806), .C(n25807), .D(n25808), .Y(n36982) );
  OR4X1 U29774 ( .A(n26887), .B(n26888), .C(n26889), .D(n26890), .Y(n36983) );
  OR4X1 U29775 ( .A(n26948), .B(n26949), .C(n26950), .D(n26951), .Y(n36984) );
  OR4X1 U29776 ( .A(n46238), .B(n46237), .C(n46236), .D(n46235), .Y(n36985) );
  OR4X1 U29777 ( .A(n25827), .B(n25828), .C(n25829), .D(n25830), .Y(n36986) );
  OR4X1 U29778 ( .A(n26007), .B(n26008), .C(n26009), .D(n26010), .Y(n36987) );
  OR4X1 U29779 ( .A(n25977), .B(n25978), .C(n25979), .D(n25980), .Y(n36988) );
  OR4X1 U29780 ( .A(n29918), .B(n29919), .C(n29920), .D(n29921), .Y(n36989) );
  OR4X1 U29781 ( .A(n29978), .B(n29979), .C(n29980), .D(n29981), .Y(n36990) );
  OR4X1 U29782 ( .A(n30038), .B(n30039), .C(n30040), .D(n30041), .Y(n36991) );
  OR4X1 U29783 ( .A(n30128), .B(n30129), .C(n30130), .D(n30131), .Y(n36992) );
  OR4X1 U29784 ( .A(n30098), .B(n30099), .C(n30100), .D(n30101), .Y(n36993) );
  OR4X1 U29785 ( .A(n25703), .B(n25704), .C(n25705), .D(n25706), .Y(n36994) );
  OR4X1 U29786 ( .A(n29290), .B(n29291), .C(n29292), .D(n29293), .Y(n36995) );
  XOR2X1 U29787 ( .A(n36837), .B(n34066), .Y(n36996) );
  XOR2X1 U29788 ( .A(n36844), .B(n33978), .Y(n36997) );
  XOR2X1 U29789 ( .A(n33962), .B(n42562), .Y(n36998) );
  XOR2X1 U29790 ( .A(n34074), .B(n42569), .Y(n36999) );
  CLKINVX1 U29791 ( .A(n42714), .Y(n42709) );
  XOR2X1 U29792 ( .A(n36858), .B(n34248), .Y(n37000) );
  XOR2X1 U29793 ( .A(n36860), .B(n34272), .Y(n37001) );
  OR4X1 U29794 ( .A(n30403), .B(n30404), .C(n30405), .D(n30406), .Y(n37002) );
  OR4X1 U29795 ( .A(n26033), .B(n26034), .C(n26035), .D(n26036), .Y(n37003) );
  OR4X1 U29796 ( .A(n26243), .B(n26244), .C(n26245), .D(n26246), .Y(n37004) );
  OR4X1 U29797 ( .A(n26213), .B(n26214), .C(n26215), .D(n26216), .Y(n37005) );
  INVX3 U29798 ( .A(n41326), .Y(n41329) );
  INVX6 U29799 ( .A(n41326), .Y(n41330) );
  OR4X1 U29800 ( .A(n26161), .B(n26162), .C(n26163), .D(n26164), .Y(n37006) );
  OR2X1 U29801 ( .A(n31865), .B(n31864), .Y(n37007) );
  OR2X1 U29802 ( .A(n28044), .B(n28043), .Y(n37008) );
  INVX6 U29803 ( .A(n41288), .Y(n41294) );
  INVX4 U29804 ( .A(n41298), .Y(n41304) );
  INVX4 U29805 ( .A(n41298), .Y(n41301) );
  INVX6 U29806 ( .A(n41298), .Y(n41302) );
  OR4X1 U29807 ( .A(n28061), .B(n28062), .C(n28063), .D(n28064), .Y(n37009) );
  OR4X1 U29808 ( .A(n27181), .B(n27182), .C(n27183), .D(n27184), .Y(n37010) );
  OR4X1 U29809 ( .A(n25917), .B(n25918), .C(n25919), .D(n25920), .Y(n37011) );
  INVX3 U29810 ( .A(n42677), .Y(n42676) );
  AO21X1 U29811 ( .A0(n48549), .A1(n10996), .B0(net209151), .Y(n37012) );
  AND2X2 U29812 ( .A(n40956), .B(net216167), .Y(n37013) );
  AO21X1 U29813 ( .A0(n48400), .A1(n10336), .B0(net171328), .Y(n37014) );
  NAND2BX2 U29814 ( .AN(n_cell_301249_net267123), .B(net213527), .Y(
        n_cell_303546_net275959) );
  NAND3X2 U29815 ( .A(net216309), .B(net216308), .C(n_cell_301249_net267441),
        .Y(n40415) );
  NAND3X2 U29816 ( .A(net216444), .B(net216443), .C(n_cell_301249_net267233),
        .Y(n39470) );
  NAND2BX2 U29817 ( .AN(n40782), .B(net216508), .Y(n11961) );
  NAND3X2 U29818 ( .A(net216253), .B(n_cell_301249_net267595), .C(net216254),
        .Y(n40418) );
  NAND3X1 U29819 ( .A(n13017), .B(n11360), .C(n12922), .Y(n10025) );
  INVX3 U29820 ( .A(n42645), .Y(n42643) );
  INVX3 U29821 ( .A(net258261), .Y(net219336) );
  NAND2BX2 U29822 ( .AN(n_cell_301249_net267619), .B(net216238), .Y(n11924) );
  NOR2X1 U29823 ( .A(net151766), .B(n37350), .Y(n37016) );
  CLKBUFX3 U29824 ( .A(n42649), .Y(n42648) );
  CLKBUFX3 U29825 ( .A(n42649), .Y(n42647) );
  CLKINVX1 U29826 ( .A(n40316), .Y(net217108) );
  CLKBUFX3 U29827 ( .A(net216996), .Y(n40368) );
  CLKINVX1 U29828 ( .A(net218152), .Y(net218074) );
  CLKINVX1 U29829 ( .A(net218146), .Y(net217988) );
  CLKINVX1 U29830 ( .A(net218156), .Y(net218118) );
  CLKINVX1 U29831 ( .A(n40183), .Y(net217954) );
  NOR2X1 U29832 ( .A(net210620), .B(net210587), .Y(n37018) );
  XOR2X1 U29833 ( .A(n32530), .B(n42564), .Y(n37021) );
  XOR2X1 U29834 ( .A(n32882), .B(n42568), .Y(n37022) );
  XOR2X1 U29835 ( .A(n32954), .B(n42567), .Y(n37023) );
  XOR2X1 U29836 ( .A(n32946), .B(n42567), .Y(n37024) );
  XOR2X1 U29837 ( .A(n36837), .B(n32674), .Y(n37025) );
  XOR2X1 U29838 ( .A(n36734), .B(n34018), .Y(n37026) );
  XOR2X1 U29839 ( .A(n36735), .B(n34074), .Y(n37027) );
  XOR2X1 U29840 ( .A(n36735), .B(n32634), .Y(n37028) );
  XOR2X1 U29841 ( .A(n36841), .B(n32978), .Y(n37029) );
  XOR2X1 U29842 ( .A(n36839), .B(n33066), .Y(n37030) );
  XOR2X1 U29843 ( .A(n36733), .B(n34026), .Y(n37031) );
  XOR2X1 U29844 ( .A(n36841), .B(n32954), .Y(n37032) );
  XOR2X1 U29845 ( .A(n36843), .B(n32962), .Y(n37033) );
  XOR2X1 U29846 ( .A(n36846), .B(n33058), .Y(n37034) );
  XOR2X1 U29847 ( .A(n36838), .B(n32994), .Y(n37035) );
  XOR2X1 U29848 ( .A(n36846), .B(n33746), .Y(n37036) );
  XOR2X1 U29849 ( .A(n36847), .B(n32970), .Y(n37037) );
  XOR2X1 U29850 ( .A(n36841), .B(n32914), .Y(n37038) );
  XOR2X1 U29851 ( .A(n36840), .B(n32770), .Y(n37039) );
  XOR2X1 U29852 ( .A(n36845), .B(n32946), .Y(n37040) );
  XOR2X1 U29853 ( .A(n36844), .B(n32930), .Y(n37041) );
  XOR2X1 U29854 ( .A(n36764), .B(n32617), .Y(n37042) );
  XOR2X1 U29855 ( .A(n36846), .B(n32722), .Y(n37043) );
  XOR2X1 U29856 ( .A(n36733), .B(n32954), .Y(n37044) );
  XOR2X1 U29857 ( .A(n36734), .B(n32946), .Y(n37045) );
  OR4X1 U29858 ( .A(n26466), .B(n26467), .C(n26468), .D(n26469), .Y(n37046) );
  OR4X1 U29859 ( .A(n29685), .B(n29686), .C(n29687), .D(n29688), .Y(n37047) );
  OR4X1 U29860 ( .A(n29746), .B(n29747), .C(n29748), .D(n29749), .Y(n37048) );
  OR4X1 U29861 ( .A(n29606), .B(n29605), .C(n29604), .D(n29603), .Y(n37049) );
  OR4X1 U29862 ( .A(n29516), .B(n29515), .C(n29514), .D(n29513), .Y(n37050) );
  OR4X1 U29863 ( .A(n29817), .B(n29816), .C(n29815), .D(n29814), .Y(n37051) );
  OR4X1 U29864 ( .A(n29787), .B(n29786), .C(n29785), .D(n29784), .Y(n37052) );
  OR4X1 U29865 ( .A(n29727), .B(n29726), .C(n29725), .D(n29724), .Y(n37053) );
  OR4X1 U29866 ( .A(n29546), .B(n29545), .C(n29544), .D(n29543), .Y(n37054) );
  OR4X1 U29867 ( .A(n23036), .B(n23035), .C(n23034), .D(n23033), .Y(n37055) );
  OR4X1 U29868 ( .A(n23026), .B(n23025), .C(n23024), .D(n23023), .Y(n37056) );
  OR4X1 U29869 ( .A(n23156), .B(n23155), .C(n23154), .D(n23153), .Y(n37057) );
  OR4X1 U29870 ( .A(n24139), .B(n24138), .C(n24137), .D(n24136), .Y(n37058) );
  OR4X1 U29871 ( .A(n23126), .B(n23125), .C(n23124), .D(n23123), .Y(n37059) );
  OR4X1 U29872 ( .A(n30358), .B(n30357), .C(n30356), .D(n30355), .Y(n37060) );
  OR4X1 U29873 ( .A(n30418), .B(n30417), .C(n30416), .D(n30415), .Y(n37061) );
  OR4X1 U29874 ( .A(n30388), .B(n30387), .C(n30386), .D(n30385), .Y(n37062) );
  OR4X1 U29875 ( .A(n21656), .B(n21655), .C(n21654), .D(n21653), .Y(n37063) );
  OR4X1 U29876 ( .A(n30480), .B(n30479), .C(n30478), .D(n30477), .Y(n37064) );
  OR4X1 U29877 ( .A(n20114), .B(n20113), .C(n20112), .D(n20111), .Y(n37065) );
  OR4X1 U29878 ( .A(n29858), .B(n29859), .C(n29860), .D(n29861), .Y(n37066) );
  OR4X1 U29879 ( .A(n29888), .B(n29889), .C(n29890), .D(n29891), .Y(n37067) );
  OR4X1 U29880 ( .A(n29828), .B(n29829), .C(n29830), .D(n29831), .Y(n37068) );
  OR4X1 U29881 ( .A(n30008), .B(n30009), .C(n30010), .D(n30011), .Y(n37069) );
  OR4X1 U29882 ( .A(n30158), .B(n30159), .C(n30160), .D(n30161), .Y(n37070) );
  OR4X1 U29883 ( .A(n21880), .B(n21879), .C(n21878), .D(n21877), .Y(n37071) );
  OR4X1 U29884 ( .A(n21890), .B(n21889), .C(n21888), .D(n21887), .Y(n37072) );
  OR4X1 U29885 ( .A(n29847), .B(n29846), .C(n29845), .D(n29844), .Y(n37073) );
  XOR2X1 U29886 ( .A(n36734), .B(n34002), .Y(n37074) );
  XOR2X1 U29887 ( .A(n36847), .B(n32666), .Y(n37075) );
  XOR2X1 U29888 ( .A(n36846), .B(n32810), .Y(n37076) );
  XOR2X1 U29889 ( .A(n36839), .B(n33682), .Y(n37077) );
  XOR2X1 U29890 ( .A(n36844), .B(n33762), .Y(n37078) );
  XOR2X1 U29891 ( .A(n36841), .B(n33754), .Y(n37079) );
  XOR2X1 U29892 ( .A(n36736), .B(n34066), .Y(n37080) );
  XOR2X1 U29893 ( .A(n36734), .B(n34010), .Y(n37081) );
  XOR2X1 U29894 ( .A(n36844), .B(n33770), .Y(n37082) );
  XOR2X1 U29895 ( .A(n36837), .B(n32882), .Y(n37083) );
  XOR2X1 U29896 ( .A(n36839), .B(n32890), .Y(n37084) );
  XOR2X1 U29897 ( .A(n36838), .B(n32594), .Y(n37085) );
  XOR2X1 U29898 ( .A(n36846), .B(n32602), .Y(n37086) );
  XOR2X1 U29899 ( .A(n36837), .B(n32898), .Y(n37087) );
  XOR2X1 U29900 ( .A(n36841), .B(n32618), .Y(n37088) );
  XOR2X1 U29901 ( .A(n36838), .B(n32826), .Y(n37089) );
  XOR2X1 U29902 ( .A(n36839), .B(n32906), .Y(n37090) );
  XOR2X1 U29903 ( .A(n36840), .B(n33050), .Y(n37091) );
  XOR2X1 U29904 ( .A(n36837), .B(n32626), .Y(n37092) );
  XOR2X1 U29905 ( .A(n36847), .B(n32834), .Y(n37093) );
  XOR2X1 U29906 ( .A(n36839), .B(n32794), .Y(n37094) );
  XOR2X1 U29907 ( .A(n36846), .B(n32866), .Y(n37095) );
  XOR2X1 U29908 ( .A(n36846), .B(n32642), .Y(n37096) );
  XOR2X1 U29909 ( .A(n36843), .B(n32634), .Y(n37097) );
  XOR2X1 U29910 ( .A(n33042), .B(n42565), .Y(n37098) );
  XOR2X1 U29911 ( .A(n33074), .B(n42568), .Y(n37099) );
  XOR2X1 U29912 ( .A(n33762), .B(n42562), .Y(n37100) );
  XOR2X1 U29913 ( .A(n33474), .B(n41630), .Y(n37101) );
  XOR2X1 U29914 ( .A(n33754), .B(n42562), .Y(n37102) );
  XOR2X1 U29915 ( .A(n33730), .B(n42562), .Y(n37103) );
  XOR2X1 U29916 ( .A(n33722), .B(n42562), .Y(n37104) );
  XOR2X1 U29917 ( .A(n33738), .B(n42562), .Y(n37105) );
  XOR2X1 U29918 ( .A(n33634), .B(n42569), .Y(n37106) );
  XOR2X1 U29919 ( .A(n33882), .B(n42568), .Y(n37107) );
  XOR2X1 U29920 ( .A(n33874), .B(n42568), .Y(n37108) );
  XOR2X1 U29921 ( .A(n33106), .B(n36725), .Y(n37109) );
  OR4X1 U29922 ( .A(n30253), .B(n30254), .C(n30255), .D(n30256), .Y(n37110) );
  OR4X1 U29923 ( .A(n26432), .B(n26433), .C(n26434), .D(n26435), .Y(n37111) );
  OR4X1 U29924 ( .A(n26183), .B(n26184), .C(n26185), .D(n26186), .Y(n37112) );
  OR4X1 U29925 ( .A(n26333), .B(n26334), .C(n26335), .D(n26336), .Y(n37113) );
  OR2X1 U29926 ( .A(n31986), .B(n31985), .Y(n37114) );
  OR2X1 U29927 ( .A(n30723), .B(n30722), .Y(n37115) );
  OR2X1 U29928 ( .A(n21405), .B(n21404), .Y(n37116) );
  OR2X1 U29929 ( .A(n30783), .B(n30782), .Y(n37117) );
  OR2X1 U29930 ( .A(n30753), .B(n30752), .Y(n37118) );
  OR2X1 U29931 ( .A(n20845), .B(n20843), .Y(n37119) );
  AND2X2 U29932 ( .A(n12207), .B(n12210), .Y(n37120) );
  AND3X2 U29933 ( .A(net216312), .B(net216311), .C(net216313), .Y(n37121) );
  AND3X2 U29934 ( .A(net216276), .B(net216275), .C(net216277), .Y(n37122) );
  AND3X2 U29935 ( .A(n10939), .B(n39542), .C(n10941), .Y(n37123) );
  AND2X2 U29936 ( .A(n40966), .B(net216365), .Y(n37124) );
  CLKINVX1 U29937 ( .A(n_cell_303546_net275956), .Y(n39677) );
  AND3X2 U29938 ( .A(net209572), .B(net209595), .C(n39460), .Y(n37125) );
  XOR2X1 U29939 ( .A(n32546), .B(n42564), .Y(n37127) );
  XOR2X1 U29940 ( .A(n32410), .B(n42562), .Y(n37128) );
  XOR2X1 U29941 ( .A(n36735), .B(n33290), .Y(n37129) );
  XOR2X1 U29942 ( .A(n36733), .B(n32562), .Y(n37130) );
  XOR2X1 U29943 ( .A(n36733), .B(n32594), .Y(n37131) );
  XOR2X1 U29944 ( .A(n36841), .B(n32746), .Y(n37132) );
  XOR2X1 U29945 ( .A(n36736), .B(n33274), .Y(n37133) );
  XOR2X1 U29946 ( .A(n36735), .B(n33002), .Y(n37134) );
  XOR2X1 U29947 ( .A(n36839), .B(n32450), .Y(n37135) );
  XOR2X1 U29948 ( .A(n36840), .B(n32474), .Y(n37136) );
  XOR2X1 U29949 ( .A(n36736), .B(n32570), .Y(n37137) );
  XOR2X1 U29950 ( .A(n36735), .B(n32514), .Y(n37138) );
  XOR2X1 U29951 ( .A(n36735), .B(n32754), .Y(n37139) );
  XOR2X1 U29952 ( .A(n36839), .B(n32402), .Y(n37140) );
  XOR2X1 U29953 ( .A(n36847), .B(n32410), .Y(n37141) );
  XOR2X1 U29954 ( .A(n36764), .B(n32585), .Y(n37142) );
  XOR2X1 U29955 ( .A(n36838), .B(n32738), .Y(n37143) );
  XOR2X1 U29956 ( .A(n36734), .B(n32994), .Y(n37144) );
  XOR2X1 U29957 ( .A(n36733), .B(n32922), .Y(n37145) );
  XOR2X1 U29958 ( .A(n36733), .B(n32914), .Y(n37146) );
  XOR2X1 U29959 ( .A(n36733), .B(n32482), .Y(n37147) );
  XOR2X1 U29960 ( .A(n36733), .B(n32938), .Y(n37148) );
  XOR2X1 U29961 ( .A(n36735), .B(n32930), .Y(n37149) );
  BUFX4 U29962 ( .A(n42465), .Y(n42459) );
  OR4X1 U29963 ( .A(n21646), .B(n21645), .C(n21644), .D(n21643), .Y(n37150) );
  OR4X1 U29964 ( .A(n20905), .B(n20904), .C(n20903), .D(n20902), .Y(n37151) );
  OR4X1 U29965 ( .A(n20463), .B(n20462), .C(n20461), .D(n20460), .Y(n37152) );
  OR4X1 U29966 ( .A(n20063), .B(n20062), .C(n20061), .D(n20060), .Y(n37153) );
  OR4X1 U29967 ( .A(n20452), .B(n20451), .C(n20450), .D(n20449), .Y(n37154) );
  OR4X1 U29968 ( .A(n21829), .B(n21828), .C(n21827), .D(n21826), .Y(n37155) );
  OR4X1 U29969 ( .A(n26544), .B(n26545), .C(n26546), .D(n26547), .Y(n37156) );
  OR4X1 U29970 ( .A(n21849), .B(n21848), .C(n21847), .D(n21846), .Y(n37157) );
  OR4X1 U29971 ( .A(n20831), .B(n20830), .C(n20829), .D(n20828), .Y(n37158) );
  XOR2X1 U29972 ( .A(n36735), .B(n33266), .Y(n37159) );
  XOR2X1 U29973 ( .A(n36845), .B(n32802), .Y(n37160) );
  XOR2X1 U29974 ( .A(n36839), .B(n32818), .Y(n37161) );
  XOR2X1 U29975 ( .A(n36837), .B(n32546), .Y(n37162) );
  XOR2X1 U29976 ( .A(n36845), .B(n32538), .Y(n37163) );
  XOR2X1 U29977 ( .A(n36843), .B(n32658), .Y(n37164) );
  XOR2X1 U29978 ( .A(n36734), .B(n33466), .Y(n37165) );
  XOR2X1 U29979 ( .A(n36840), .B(n32530), .Y(n37166) );
  XOR2X1 U29980 ( .A(n36838), .B(n33706), .Y(n37167) );
  XOR2X1 U29981 ( .A(n36845), .B(n33698), .Y(n37168) );
  XOR2X1 U29982 ( .A(n36846), .B(n32842), .Y(n37169) );
  XOR2X1 U29983 ( .A(n36843), .B(n32786), .Y(n37170) );
  XOR2X1 U29984 ( .A(n36840), .B(n33002), .Y(n37171) );
  BUFX4 U29985 ( .A(n42478), .Y(n42490) );
  NAND4X1 U29986 ( .A(n43204), .B(n43203), .C(n43202), .D(n43201), .Y(
        net214729) );
  NAND4BX1 U29987 ( .AN(n41672), .B(n44577), .C(n44576), .D(n44575), .Y(n12549) );
  CLKINVX1 U29988 ( .A(n12549), .Y(net171314) );
  OR2X1 U29989 ( .A(n21790), .B(n21788), .Y(n37172) );
  OR2X1 U29990 ( .A(n20035), .B(n20034), .Y(n37173) );
  OR2X1 U29991 ( .A(n20025), .B(n20024), .Y(n37174) );
  OR2X1 U29992 ( .A(n21811), .B(n21810), .Y(n37175) );
  OR2X1 U29993 ( .A(n20496), .B(n20495), .Y(n37176) );
  OR2X1 U29994 ( .A(n20813), .B(n20811), .Y(n37177) );
  OR2X1 U29995 ( .A(n20823), .B(n20822), .Y(n37178) );
  CLKINVX1 U29996 ( .A(n11265), .Y(n39343) );
  INVX3 U29997 ( .A(n10206), .Y(net151584) );
  CLKINVX1 U29998 ( .A(n11942), .Y(n39605) );
  CLKINVX1 U29999 ( .A(n11959), .Y(n39555) );
  CLKINVX1 U30000 ( .A(n10974), .Y(n39483) );
  OR2X1 U30001 ( .A(net151509), .B(net151503), .Y(n37179) );
  XOR2X1 U30002 ( .A(n36734), .B(n32418), .Y(n37180) );
  NAND2BX1 U30003 ( .AN(n40446), .B(net210368), .Y(n12826) );
  CLKINVX1 U30004 ( .A(n12826), .Y(net151809) );
  CLKINVX1 U30005 ( .A(n11568), .Y(net171280) );
  NAND2BX1 U30006 ( .AN(n_cell_301249_net267397), .B(net216319), .Y(n10480) );
  NAND2BX1 U30007 ( .AN(n_cell_301249_net267391), .B(net212154), .Y(n12165) );
  CLKINVX1 U30008 ( .A(n12165), .Y(net151542) );
  AND3X2 U30009 ( .A(net259641), .B(net259645), .C(net151275), .Y(n37181) );
  NOR2X4 U30010 ( .A(n19334), .B(n50145), .Y(n37182) );
  NAND2X4 U30011 ( .A(n19411), .B(n41796), .Y(n37183) );
  CLKBUFX3 U30012 ( .A(net221740), .Y(net264712) );
  CLKBUFX3 U30013 ( .A(net221744), .Y(net264742) );
  CLKINVX1 U30014 ( .A(net266151), .Y(net221730) );
  CLKINVX1 U30015 ( .A(net266151), .Y(net221718) );
  CLKINVX1 U30016 ( .A(net266151), .Y(net221734) );
  CLKBUFX3 U30017 ( .A(n34130), .Y(n42063) );
  AND2X2 U30018 ( .A(n44841), .B(n44840), .Y(n37196) );
  AND3X2 U30019 ( .A(n44869), .B(n44872), .C(n44870), .Y(n37197) );
  OR4X1 U30020 ( .A(n45323), .B(n45322), .C(n45321), .D(n45320), .Y(n37198) );
  NAND4X1 U30021 ( .A(n44814), .B(n44813), .C(n44812), .D(n44811), .Y(
        net210650) );
  CLKINVX1 U30022 ( .A(net211197), .Y(net171489) );
  AND4X1 U30023 ( .A(n47242), .B(n47241), .C(n47240), .D(n47239), .Y(n37199)
         );
  NAND2BX1 U30024 ( .AN(n39425), .B(net213342), .Y(n10869) );
  CLKINVX1 U30025 ( .A(n10869), .Y(n39953) );
  CLKBUFX3 U30026 ( .A(n34399), .Y(n41808) );
  CLKBUFX3 U30027 ( .A(n34411), .Y(n42064) );
  CLKBUFX3 U30028 ( .A(n34339), .Y(n42073) );
  CLKBUFX3 U30029 ( .A(n33567), .Y(n41911) );
  AND3X2 U30030 ( .A(n46339), .B(n46340), .C(n46341), .Y(n37204) );
  NAND4X1 U30031 ( .A(n44090), .B(n44089), .C(n44088), .D(n44087), .Y(
        net210643) );
  CLKINVX1 U30032 ( .A(net210643), .Y(n39479) );
  AND4X1 U30033 ( .A(n47227), .B(n47226), .C(n47225), .D(n47224), .Y(n37205)
         );
  NAND4X1 U30034 ( .A(n45807), .B(n45806), .C(n45805), .D(n45804), .Y(n11075)
         );
  CLKINVX1 U30035 ( .A(n11075), .Y(n39491) );
  OR3X2 U30036 ( .A(n43892), .B(n43893), .C(n43890), .Y(n37206) );
  OR2X1 U30037 ( .A(n26794), .B(n26793), .Y(n37207) );
  AND3X2 U30038 ( .A(n43838), .B(n43839), .C(n43840), .Y(n37208) );
  XNOR2X1 U30039 ( .A(n41868), .B(n42515), .Y(n37209) );
  XNOR2X1 U30040 ( .A(n41882), .B(n42522), .Y(n37210) );
  OR4X1 U30041 ( .A(n46382), .B(n46381), .C(n46380), .D(n46379), .Y(n37211) );
  OR4X1 U30042 ( .A(n29402), .B(n29403), .C(n29404), .D(n29405), .Y(n37212) );
  OR4X1 U30043 ( .A(n27305), .B(n27306), .C(n27307), .D(n27308), .Y(n37213) );
  OR4X1 U30044 ( .A(n27516), .B(n27517), .C(n27518), .D(n27519), .Y(n37214) );
  OR4X1 U30045 ( .A(n27396), .B(n27397), .C(n27398), .D(n27399), .Y(n37215) );
  OR4X1 U30046 ( .A(n31660), .B(n31661), .C(n31662), .D(n31663), .Y(n37216) );
  AND2X2 U30047 ( .A(n45688), .B(n45689), .Y(n37217) );
  NAND3X1 U30048 ( .A(n39297), .B(net215225), .C(net215222), .Y(n10554) );
  CLKINVX1 U30049 ( .A(n10554), .Y(n39806) );
  OR4X1 U30050 ( .A(n27155), .B(n27156), .C(n27157), .D(n27158), .Y(n37218) );
  OR4X1 U30051 ( .A(n27365), .B(n27366), .C(n27367), .D(n27368), .Y(n37219) );
  OR4X1 U30052 ( .A(n28027), .B(n28028), .C(n28029), .D(n28030), .Y(n37220) );
  OA21XL U30053 ( .A0(n48155), .A1(n48154), .B0(n48153), .Y(n37221) );
  OR2X1 U30054 ( .A(n27383), .B(n27382), .Y(n37222) );
  OR2X1 U30055 ( .A(n27202), .B(n27201), .Y(n37223) );
  OR2X1 U30056 ( .A(n27322), .B(n27321), .Y(n37224) );
  OR2X1 U30057 ( .A(n27352), .B(n27351), .Y(n37225) );
  OR2X1 U30058 ( .A(n46385), .B(n46384), .Y(n37226) );
  OR2X1 U30059 ( .A(n28074), .B(n28073), .Y(n37227) );
  OR2X1 U30060 ( .A(n46234), .B(n46233), .Y(n37228) );
  OR2X1 U30061 ( .A(n46465), .B(n46464), .Y(n37229) );
  OR4X1 U30062 ( .A(n29294), .B(n29295), .C(n29296), .D(n29297), .Y(n37230) );
  OR4X1 U30063 ( .A(n28057), .B(n28058), .C(n28059), .D(n28060), .Y(n37231) );
  OR4X1 U30064 ( .A(n27177), .B(n27178), .C(n27179), .D(n27180), .Y(n37232) );
  INVX6 U30065 ( .A(n41326), .Y(n41332) );
  AO21X1 U30066 ( .A0(n47724), .A1(n47723), .B0(net210680), .Y(n37233) );
  INVX3 U30067 ( .A(n41289), .Y(n41295) );
  INVX6 U30068 ( .A(n41288), .Y(n41293) );
  OR4X1 U30069 ( .A(n45097), .B(n45096), .C(n45095), .D(n45094), .Y(n37234) );
  INVX6 U30070 ( .A(n41298), .Y(n41300) );
  INVX4 U30071 ( .A(n41298), .Y(n41299) );
  AND2X2 U30072 ( .A(n44964), .B(n44963), .Y(n37235) );
  OR4X1 U30073 ( .A(n27546), .B(n27547), .C(n27548), .D(n27549), .Y(n37236) );
  NOR2X1 U30074 ( .A(n46248), .B(n46247), .Y(n37237) );
  NOR2X1 U30075 ( .A(n12951), .B(n37205), .Y(n11418) );
  NAND2BX2 U30076 ( .AN(n39305), .B(net215822), .Y(n39304) );
  CLKINVX1 U30077 ( .A(net258261), .Y(net219324) );
  NAND4X1 U30078 ( .A(n45817), .B(n45816), .C(n45815), .D(n45814), .Y(n11073)
         );
  OR2X1 U30079 ( .A(n39912), .B(net151426), .Y(n37239) );
  AND4X1 U30080 ( .A(n46778), .B(n46777), .C(n46776), .D(n46775), .Y(n37240)
         );
  NAND2X2 U30081 ( .A(n41736), .B(net260384), .Y(n37241) );
  CLKBUFX3 U30082 ( .A(n33947), .Y(n42122) );
  CLKBUFX3 U30083 ( .A(n33635), .Y(n42161) );
  CLKBUFX3 U30084 ( .A(n33951), .Y(n41863) );
  CLKBUFX3 U30085 ( .A(n33847), .Y(n41876) );
  CLKBUFX3 U30086 ( .A(n33883), .Y(n42130) );
  NAND4X1 U30087 ( .A(n44560), .B(n44559), .C(n44558), .D(n44557), .Y(n12703)
         );
  CLKINVX1 U30088 ( .A(n12703), .Y(n39561) );
  NAND4X1 U30089 ( .A(n46713), .B(n46712), .C(n46711), .D(n46710), .Y(n13018)
         );
  CLKINVX1 U30090 ( .A(n13018), .Y(n39631) );
  NAND4X1 U30091 ( .A(n43549), .B(n43548), .C(n43547), .D(n43546), .Y(n11848)
         );
  CLKINVX1 U30092 ( .A(n11848), .Y(net209659) );
  NAND2BX1 U30093 ( .AN(n40440), .B(net211623), .Y(net209996) );
  INVX3 U30094 ( .A(net209996), .Y(n40710) );
  NAND4X1 U30095 ( .A(n43740), .B(n43739), .C(n43738), .D(n43737), .Y(n12017)
         );
  CLKINVX1 U30096 ( .A(n12017), .Y(n39560) );
  NAND2BX1 U30097 ( .AN(n39377), .B(net211651), .Y(n10752) );
  CLKINVX1 U30098 ( .A(n10752), .Y(n39900) );
  NAND4X1 U30099 ( .A(net215465), .B(net215466), .C(net215467), .D(net215468),
        .Y(n10394) );
  XNOR2X1 U30100 ( .A(n41867), .B(n42515), .Y(n37254) );
  NAND4X1 U30101 ( .A(n46097), .B(n46096), .C(n46095), .D(n46094), .Y(n11200)
         );
  CLKINVX1 U30102 ( .A(n11388), .Y(n39636) );
  AND3X2 U30103 ( .A(n43674), .B(n43675), .C(n43676), .Y(n37255) );
  NAND4X1 U30104 ( .A(n43628), .B(n43627), .C(n43626), .D(n43625), .Y(n12535)
         );
  OR4X1 U30105 ( .A(n26658), .B(n26657), .C(n26656), .D(n26655), .Y(n37256) );
  OR4X1 U30106 ( .A(n30691), .B(n30690), .C(n30689), .D(n30688), .Y(n37257) );
  OR4X1 U30107 ( .A(n30208), .B(n30207), .C(n30206), .D(n30205), .Y(n37258) );
  OR4X1 U30108 ( .A(n29557), .B(n29558), .C(n29559), .D(n29560), .Y(n37259) );
  OR4X1 U30109 ( .A(n26823), .B(n26824), .C(n26825), .D(n26826), .Y(n37260) );
  OR4X1 U30110 ( .A(n26944), .B(n26945), .C(n26946), .D(n26947), .Y(n37261) );
  OR4X1 U30111 ( .A(n30698), .B(n30699), .C(n30700), .D(n30701), .Y(n37262) );
  OR4X1 U30112 ( .A(n30728), .B(n30729), .C(n30730), .D(n30731), .Y(n37263) );
  OR4X1 U30113 ( .A(n30758), .B(n30759), .C(n30760), .D(n30761), .Y(n37264) );
  OR4X1 U30114 ( .A(n29772), .B(n29773), .C(n29774), .D(n29775), .Y(n37265) );
  OR4X1 U30115 ( .A(n30365), .B(n30366), .C(n30367), .D(n30368), .Y(n37266) );
  OR4X1 U30116 ( .A(n30335), .B(n30336), .C(n30337), .D(n30338), .Y(n37267) );
  OR4X1 U30117 ( .A(n30425), .B(n30426), .C(n30427), .D(n30428), .Y(n37268) );
  OR4X1 U30118 ( .A(n29711), .B(n29712), .C(n29713), .D(n29714), .Y(n37269) );
  OR4X1 U30119 ( .A(n29681), .B(n29682), .C(n29683), .D(n29684), .Y(n37270) );
  OR4X1 U30120 ( .A(n29742), .B(n29743), .C(n29744), .D(n29745), .Y(n37271) );
  OR4X1 U30121 ( .A(n29531), .B(n29532), .C(n29533), .D(n29534), .Y(n37272) );
  OR4X1 U30122 ( .A(n30457), .B(n30458), .C(n30459), .D(n30460), .Y(n37273) );
  OR4X1 U30123 ( .A(n30637), .B(n30638), .C(n30639), .D(n30640), .Y(n37274) );
  OR4X1 U30124 ( .A(n30547), .B(n30548), .C(n30549), .D(n30550), .Y(n37275) );
  OR4X1 U30125 ( .A(n29651), .B(n29652), .C(n29653), .D(n29654), .Y(n37276) );
  OR4X1 U30126 ( .A(n31720), .B(n31721), .C(n31722), .D(n31723), .Y(n37277) );
  OR4X1 U30127 ( .A(n31810), .B(n31811), .C(n31812), .D(n31813), .Y(n37278) );
  OR4X1 U30128 ( .A(n30878), .B(n30879), .C(n30880), .D(n30881), .Y(n37279) );
  OR4X1 U30129 ( .A(n30667), .B(n30668), .C(n30669), .D(n30670), .Y(n37280) );
  OR4X1 U30130 ( .A(n30487), .B(n30488), .C(n30489), .D(n30490), .Y(n37281) );
  OR4X1 U30131 ( .A(n30818), .B(n30819), .C(n30820), .D(n30821), .Y(n37282) );
  OR4X1 U30132 ( .A(n30848), .B(n30849), .C(n30850), .D(n30851), .Y(n37283) );
  OR4X1 U30133 ( .A(n25823), .B(n25824), .C(n25825), .D(n25826), .Y(n37284) );
  OR4X1 U30134 ( .A(n29892), .B(n29893), .C(n29894), .D(n29895), .Y(n37285) );
  OR4X1 U30135 ( .A(n29832), .B(n29833), .C(n29834), .D(n29835), .Y(n37286) );
  OR4X1 U30136 ( .A(n25913), .B(n25914), .C(n25915), .D(n25916), .Y(n37287) );
  OR4X1 U30137 ( .A(n26462), .B(n26463), .C(n26464), .D(n26465), .Y(n37288) );
  OR4X1 U30138 ( .A(n26522), .B(n26523), .C(n26524), .D(n26525), .Y(n37289) );
  OR4X1 U30139 ( .A(n26003), .B(n26004), .C(n26005), .D(n26006), .Y(n37290) );
  OR4X1 U30140 ( .A(n25973), .B(n25974), .C(n25975), .D(n25976), .Y(n37291) );
  OR4X1 U30141 ( .A(n29922), .B(n29923), .C(n29924), .D(n29925), .Y(n37292) );
  OR4X1 U30142 ( .A(n29982), .B(n29983), .C(n29984), .D(n29985), .Y(n37293) );
  OR4X1 U30143 ( .A(n30034), .B(n30035), .C(n30036), .D(n30037), .Y(n37294) );
  OR4X1 U30144 ( .A(n30004), .B(n30005), .C(n30006), .D(n30007), .Y(n37295) );
  OR4X1 U30145 ( .A(n30124), .B(n30125), .C(n30126), .D(n30127), .Y(n37296) );
  OR4X1 U30146 ( .A(n30094), .B(n30095), .C(n30096), .D(n30097), .Y(n37297) );
  OR4X1 U30147 ( .A(n30154), .B(n30155), .C(n30156), .D(n30157), .Y(n37298) );
  AND2X2 U30148 ( .A(n44498), .B(n44497), .Y(n37299) );
  NAND4X1 U30149 ( .A(n47138), .B(n47137), .C(n47136), .D(n47135), .Y(n11416)
         );
  XOR2X1 U30150 ( .A(n36734), .B(n33962), .Y(n37300) );
  CLKINVX1 U30151 ( .A(n12278), .Y(net151458) );
  XOR2X1 U30152 ( .A(n34066), .B(n42569), .Y(n37301) );
  OR4X1 U30153 ( .A(n26974), .B(n26975), .C(n26976), .D(n26977), .Y(n37302) );
  OR4X1 U30154 ( .A(n27094), .B(n27095), .C(n27096), .D(n27097), .Y(n37303) );
  OR4X1 U30155 ( .A(n26914), .B(n26915), .C(n26916), .D(n26917), .Y(n37304) );
  OR4X1 U30156 ( .A(n29591), .B(n29592), .C(n29593), .D(n29594), .Y(n37305) );
  OR4X1 U30157 ( .A(n31156), .B(n31157), .C(n31158), .D(n31159), .Y(n37306) );
  OR4X1 U30158 ( .A(n26153), .B(n26154), .C(n26155), .D(n26156), .Y(n37307) );
  OR2X1 U30159 ( .A(n26870), .B(n26869), .Y(n37308) );
  OR2X1 U30160 ( .A(n25007), .B(n25006), .Y(n37309) );
  OR2X1 U30161 ( .A(n26810), .B(n26809), .Y(n37310) );
  OR2X1 U30162 ( .A(n29277), .B(n29276), .Y(n37311) );
  OR2X1 U30163 ( .A(n32016), .B(n32015), .Y(n37312) );
  OR2X1 U30164 ( .A(n29247), .B(n29246), .Y(n37313) );
  OR2X1 U30165 ( .A(n26901), .B(n26900), .Y(n37314) );
  OR2X1 U30166 ( .A(n23738), .B(n23737), .Y(n37315) );
  OR2X1 U30167 ( .A(n26931), .B(n26930), .Y(n37316) );
  OR2X1 U30168 ( .A(n23839), .B(n23838), .Y(n37317) );
  OR2X1 U30169 ( .A(n23128), .B(n23127), .Y(n37318) );
  OR2X1 U30170 ( .A(n28345), .B(n28344), .Y(n37319) );
  OR2X1 U30171 ( .A(n26961), .B(n26960), .Y(n37320) );
  OR2X1 U30172 ( .A(n30662), .B(n30661), .Y(n37321) );
  OR2X1 U30173 ( .A(n30420), .B(n30419), .Y(n37322) );
  OR2X1 U30174 ( .A(n30632), .B(n30631), .Y(n37323) );
  OR2X1 U30175 ( .A(n29488), .B(n29487), .Y(n37324) );
  OR2X1 U30176 ( .A(n20271), .B(n20270), .Y(n37325) );
  OR2X1 U30177 ( .A(n20281), .B(n20280), .Y(n37326) );
  OR2X1 U30178 ( .A(n20229), .B(n20228), .Y(n37327) );
  OR2X1 U30179 ( .A(n20239), .B(n20238), .Y(n37328) );
  OR2X1 U30180 ( .A(n20249), .B(n20248), .Y(n37329) );
  OR2X1 U30181 ( .A(n20260), .B(n20258), .Y(n37330) );
  OR2X1 U30182 ( .A(n29548), .B(n29547), .Y(n37331) );
  OR4X1 U30183 ( .A(n26883), .B(n26884), .C(n26885), .D(n26886), .Y(n37332) );
  OR2X1 U30184 ( .A(n26840), .B(n26839), .Y(n37333) );
  OR2X1 U30185 ( .A(n23748), .B(n23747), .Y(n37334) );
  NAND2BX1 U30186 ( .AN(n_cell_301249_net267948), .B(net215060), .Y(n11906) );
  CLKINVX1 U30187 ( .A(n11906), .Y(n_cell_303546_net277854) );
  OR2X1 U30188 ( .A(n23768), .B(n23767), .Y(n37335) );
  OR2X1 U30189 ( .A(net259665), .B(n43545), .Y(n37336) );
  OR2X1 U30190 ( .A(n39444), .B(n43463), .Y(n37337) );
  NAND2BX1 U30191 ( .AN(n_cell_301249_net267275), .B(net212174), .Y(n11282) );
  CLKINVX1 U30192 ( .A(n40315), .Y(net217056) );
  CLKINVX1 U30193 ( .A(n40316), .Y(net217032) );
  CLKINVX1 U30194 ( .A(n40316), .Y(net217028) );
  CLKINVX1 U30195 ( .A(n40316), .Y(net217030) );
  AND3X2 U30196 ( .A(net216267), .B(net216266), .C(net216268), .Y(n37338) );
  AND3X2 U30197 ( .A(net216258), .B(net216257), .C(net216259), .Y(n37339) );
  AND3X2 U30198 ( .A(net215080), .B(net215079), .C(net215081), .Y(n37340) );
  AND3X2 U30199 ( .A(net215071), .B(net215070), .C(net215072), .Y(n37341) );
  CLKBUFX3 U30200 ( .A(net218782), .Y(n40078) );
  AND2X2 U30201 ( .A(n10612), .B(n10613), .Y(n37342) );
  CLKINVX1 U30202 ( .A(n11049), .Y(n39520) );
  CLKBUFX3 U30203 ( .A(net209103), .Y(net260830) );
  NAND3X2 U30204 ( .A(net214767), .B(n_cell_301249_net267786), .C(net214766),
        .Y(n_cell_303546_net276365) );
  NAND4X1 U30205 ( .A(n11365), .B(n11366), .C(n11510), .D(n11509), .Y(n10026)
         );
  OR2X1 U30206 ( .A(net171542), .B(net238789), .Y(n37343) );
  NAND2BX2 U30207 ( .AN(n_cell_301249_net267966), .B(net211608), .Y(n39341) );
  NAND2BX1 U30208 ( .AN(n39346), .B(net210497), .Y(n10662) );
  CLKINVX1 U30209 ( .A(n10662), .Y(n39916) );
  NAND3BX1 U30210 ( .AN(n47731), .B(n48305), .C(n47727), .Y(net210392) );
  OR2X1 U30211 ( .A(n37240), .B(net171532), .Y(n37344) );
  CLKINVX1 U30212 ( .A(n40177), .Y(net217952) );
  CLKINVX1 U30213 ( .A(n40183), .Y(net217964) );
  CLKINVX1 U30214 ( .A(n40176), .Y(net217942) );
  CLKINVX1 U30215 ( .A(n40183), .Y(net217956) );
  OR2X1 U30216 ( .A(n47774), .B(n47772), .Y(net210416) );
  NAND3X2 U30217 ( .A(net216226), .B(n_cell_301249_net267589), .C(net216225),
        .Y(n40422) );
  NAND2BX2 U30218 ( .AN(n_cell_301249_net268023), .B(net213225), .Y(n10928) );
  NAND2BX2 U30219 ( .AN(n_cell_301249_net267706), .B(net213618), .Y(n10947) );
  NOR4X1 U30220 ( .A(net171546), .B(net171547), .C(net151721), .D(net151720),
        .Y(n37345) );
  AND3X2 U30221 ( .A(net260830), .B(net211602), .C(n39543), .Y(n37346) );
  NAND2BX2 U30222 ( .AN(n_cell_301249_net267562), .B(net213462), .Y(n10957) );
  NOR2X1 U30223 ( .A(net171152), .B(net171153), .Y(n37347) );
  NOR4X1 U30224 ( .A(net171439), .B(net151767), .C(net151772), .D(net171437),
        .Y(n37348) );
  NOR3X1 U30225 ( .A(net171252), .B(net151757), .C(n39575), .Y(n37349) );
  NAND4X1 U30226 ( .A(n45752), .B(n45751), .C(n45750), .D(n45749), .Y(n11094)
         );
  OR3X2 U30227 ( .A(net151769), .B(net171544), .C(net171545), .Y(n37350) );
  OR2X1 U30228 ( .A(net151790), .B(net151793), .Y(n37351) );
  OR2X1 U30229 ( .A(net151550), .B(net151555), .Y(n37352) );
  OR2X1 U30230 ( .A(n37011), .B(n37287), .Y(n37353) );
  OR2X1 U30231 ( .A(n37343), .B(net151806), .Y(n37354) );
  OR4X1 U30232 ( .A(net171408), .B(net151571), .C(net151566), .D(net171406),
        .Y(n39537) );
  CLKINVX1 U30233 ( .A(n12799), .Y(net171127) );
  CLKINVX1 U30234 ( .A(n12388), .Y(net171448) );
  CLKINVX1 U30235 ( .A(n12085), .Y(net209844) );
  CLKINVX1 U30236 ( .A(n11015), .Y(n39485) );
  NAND2BX1 U30237 ( .AN(n39383), .B(net211997), .Y(n10755) );
  CLKINVX1 U30238 ( .A(n10755), .Y(n39908) );
  CLKINVX1 U30239 ( .A(n12665), .Y(n39335) );
  CLKINVX1 U30240 ( .A(n12280), .Y(n39488) );
  NAND2BX1 U30241 ( .AN(n39328), .B(net215912), .Y(n10529) );
  CLKINVX1 U30242 ( .A(n10529), .Y(n39815) );
  NAND4X1 U30243 ( .A(n44479), .B(n44478), .C(n44477), .D(n44476), .Y(n12518)
         );
  CLKINVX1 U30244 ( .A(n12518), .Y(net209509) );
  CLKINVX1 U30245 ( .A(n11066), .Y(net209203) );
  XOR2X1 U30246 ( .A(n51338), .B(n41305), .Y(n37355) );
  NAND3X1 U30247 ( .A(net215294), .B(net215295), .C(n39468), .Y(n10422) );
  CLKINVX1 U30248 ( .A(n12251), .Y(net151494) );
  NAND4X1 U30249 ( .A(n46874), .B(n46873), .C(n46872), .D(n46871), .Y(n11516)
         );
  CLKINVX1 U30250 ( .A(n11516), .Y(n39628) );
  NAND4X1 U30251 ( .A(n44511), .B(n44510), .C(n44509), .D(n44508), .Y(n11717)
         );
  XOR2X1 U30252 ( .A(n32738), .B(n42560), .Y(n37356) );
  XOR2X1 U30253 ( .A(n32674), .B(n42560), .Y(n37357) );
  XOR2X1 U30254 ( .A(n32434), .B(n42565), .Y(n37358) );
  XOR2X1 U30255 ( .A(n32538), .B(n42564), .Y(n37359) );
  XOR2X1 U30256 ( .A(n32722), .B(n42560), .Y(n37360) );
  XOR2X1 U30257 ( .A(n32482), .B(n42563), .Y(n37361) );
  XOR2X1 U30258 ( .A(n32474), .B(n42563), .Y(n37362) );
  XOR2X1 U30259 ( .A(n32466), .B(n42563), .Y(n37363) );
  NAND4X1 U30260 ( .A(n44255), .B(n44254), .C(n44253), .D(n44252), .Y(n11731)
         );
  CLKINVX1 U30261 ( .A(n11731), .Y(net209513) );
  NAND4X1 U30262 ( .A(n43731), .B(n43730), .C(n43729), .D(n43728), .Y(n12016)
         );
  NAND4X1 U30263 ( .A(n45721), .B(n45720), .C(n45719), .D(n45718), .Y(n12387)
         );
  NAND4X1 U30264 ( .A(n45802), .B(n45801), .C(n45800), .D(n45799), .Y(n11074)
         );
  OR4X1 U30265 ( .A(n22673), .B(n22672), .C(n22671), .D(n22670), .Y(n37364) );
  OR4X1 U30266 ( .A(n22092), .B(n22091), .C(n22090), .D(n22089), .Y(n37365) );
  OR4X1 U30267 ( .A(n24233), .B(n24232), .C(n24231), .D(n24230), .Y(n37366) );
  OR4X1 U30268 ( .A(n25711), .B(n25712), .C(n25713), .D(n25714), .Y(n37367) );
  OR4X1 U30269 ( .A(n21272), .B(n21271), .C(n21270), .D(n21269), .Y(n37368) );
  OR4X1 U30270 ( .A(n24223), .B(n24222), .C(n24221), .D(n24220), .Y(n37369) );
  OR4X1 U30271 ( .A(n21252), .B(n21251), .C(n21250), .D(n21249), .Y(n37370) );
  OR4X1 U30272 ( .A(n21282), .B(n21281), .C(n21280), .D(n21279), .Y(n37371) );
  OR4X1 U30273 ( .A(n21262), .B(n21261), .C(n21260), .D(n21259), .Y(n37372) );
  OR4X1 U30274 ( .A(n21222), .B(n21221), .C(n21220), .D(n21219), .Y(n37373) );
  OR4X1 U30275 ( .A(n21212), .B(n21211), .C(n21210), .D(n21209), .Y(n37374) );
  OR4X1 U30276 ( .A(n21676), .B(n21675), .C(n21674), .D(n21673), .Y(n37375) );
  OR4X1 U30277 ( .A(n20895), .B(n20894), .C(n20893), .D(n20892), .Y(n37376) );
  OR4X1 U30278 ( .A(n24545), .B(n24544), .C(n24543), .D(n24542), .Y(n37377) );
  OR4X1 U30279 ( .A(n21951), .B(n21950), .C(n21949), .D(n21948), .Y(n37378) );
  OR4X1 U30280 ( .A(n22031), .B(n22030), .C(n22029), .D(n22028), .Y(n37379) );
  OR4X1 U30281 ( .A(n26552), .B(n26553), .C(n26554), .D(n26555), .Y(n37380) );
  OR4X1 U30282 ( .A(n25801), .B(n25802), .C(n25803), .D(n25804), .Y(n37381) );
  OR4X1 U30283 ( .A(n29862), .B(n29863), .C(n29864), .D(n29865), .Y(n37382) );
  CLKINVX1 U30284 ( .A(n39657), .Y(n10033) );
  OR2X1 U30285 ( .A(net151857), .B(n39658), .Y(n39657) );
  XOR2X1 U30286 ( .A(n36735), .B(n33106), .Y(n37383) );
  XOR2X1 U30287 ( .A(n36735), .B(n33034), .Y(n37384) );
  XOR2X1 U30288 ( .A(n36736), .B(n32658), .Y(n37385) );
  XOR2X1 U30289 ( .A(n36736), .B(n32674), .Y(n37386) );
  XOR2X1 U30290 ( .A(n36733), .B(n32730), .Y(n37387) );
  XOR2X1 U30291 ( .A(n33130), .B(n36725), .Y(n37388) );
  XOR2X1 U30292 ( .A(n33034), .B(n42569), .Y(n37389) );
  XOR2X1 U30293 ( .A(n33018), .B(n42569), .Y(n37390) );
  XOR2X1 U30294 ( .A(n33026), .B(n42569), .Y(n37391) );
  XOR2X1 U30295 ( .A(n33274), .B(n42568), .Y(n37392) );
  NAND4BX1 U30296 ( .AN(n37305), .B(net216201), .C(net216198), .D(net216199),
        .Y(n11585) );
  CLKINVX1 U30297 ( .A(n11585), .Y(n_cell_301249_net269635) );
  NAND4X1 U30298 ( .A(n43638), .B(n43637), .C(n43636), .D(n43635), .Y(n12583)
         );
  NAND2BX2 U30299 ( .AN(n41199), .B(net266255), .Y(net209402) );
  NAND4BX1 U30300 ( .AN(n41666), .B(n44609), .C(n44608), .D(n44607), .Y(n11742) );
  NAND4BX1 U30301 ( .AN(n41670), .B(n44574), .C(n44573), .D(n44572), .Y(n11778) );
  CLKINVX1 U30302 ( .A(n11778), .Y(net209638) );
  CLKBUFX3 U30303 ( .A(n42479), .Y(n42483) );
  OR4X1 U30304 ( .A(n26612), .B(n26613), .C(n26614), .D(n26615), .Y(n37393) );
  OR4X1 U30305 ( .A(n26041), .B(n26042), .C(n26043), .D(n26044), .Y(n37394) );
  OR4X1 U30306 ( .A(n26191), .B(n26192), .C(n26193), .D(n26194), .Y(n37395) );
  OR4X1 U30307 ( .A(n26251), .B(n26252), .C(n26253), .D(n26254), .Y(n37396) );
  OR4X1 U30308 ( .A(n26221), .B(n26222), .C(n26223), .D(n26224), .Y(n37397) );
  OR4X1 U30309 ( .A(n26341), .B(n26342), .C(n26343), .D(n26344), .Y(n37398) );
  OR4X1 U30310 ( .A(n26424), .B(n26425), .C(n26426), .D(n26427), .Y(n37399) );
  OR2X1 U30311 ( .A(n22084), .B(n22082), .Y(n37400) );
  OR2X1 U30312 ( .A(n21749), .B(n21748), .Y(n37401) );
  OR2X1 U30313 ( .A(n21779), .B(n21778), .Y(n37402) );
  OR2X1 U30314 ( .A(n21688), .B(n21687), .Y(n37403) );
  OR2X1 U30315 ( .A(n21769), .B(n21768), .Y(n37404) );
  OR2X1 U30316 ( .A(n24152), .B(n24151), .Y(n37405) );
  OR2X1 U30317 ( .A(n20045), .B(n20044), .Y(n37406) );
  OR2X1 U30318 ( .A(n23038), .B(n23037), .Y(n37407) );
  OR2X1 U30319 ( .A(n24142), .B(n24140), .Y(n37408) );
  OR2X1 U30320 ( .A(n24173), .B(n24171), .Y(n37409) );
  OR2X1 U30321 ( .A(n20939), .B(n20938), .Y(n37410) );
  OR2X1 U30322 ( .A(n19972), .B(n19971), .Y(n37411) );
  OR2X1 U30323 ( .A(n23158), .B(n23157), .Y(n37412) );
  OR2X1 U30324 ( .A(n32316), .B(n32315), .Y(n37413) );
  OR2X1 U30325 ( .A(n22645), .B(n22644), .Y(n37414) );
  OR2X1 U30326 ( .A(n22665), .B(n22664), .Y(n37415) );
  OR2X1 U30327 ( .A(n22655), .B(n22654), .Y(n37416) );
  OR2X1 U30328 ( .A(n30482), .B(n30481), .Y(n37417) );
  OR2X1 U30329 ( .A(n22634), .B(n22633), .Y(n37418) );
  OR2X1 U30330 ( .A(n22624), .B(n22623), .Y(n37419) );
  OR2X1 U30331 ( .A(n22614), .B(n22613), .Y(n37420) );
  OR2X1 U30332 ( .A(n26539), .B(n26538), .Y(n37421) );
  OR2X1 U30333 ( .A(n20929), .B(n20927), .Y(n37422) );
  OR2X1 U30334 ( .A(n25758), .B(n25757), .Y(n37423) );
  OR2X1 U30335 ( .A(n25698), .B(n25697), .Y(n37424) );
  OR2X1 U30336 ( .A(n32256), .B(n32255), .Y(n37425) );
  OR2X1 U30337 ( .A(n30390), .B(n30389), .Y(n37426) );
  OR2X1 U30338 ( .A(n30360), .B(n30359), .Y(n37427) );
  OR2X1 U30339 ( .A(n22553), .B(n22552), .Y(n37428) );
  OR2X1 U30340 ( .A(n22533), .B(n22532), .Y(n37429) );
  OR2X1 U30341 ( .A(n22543), .B(n22542), .Y(n37430) );
  OR2X1 U30342 ( .A(n22513), .B(n22512), .Y(n37431) );
  OR2X1 U30343 ( .A(n22503), .B(n22502), .Y(n37432) );
  OR2X1 U30344 ( .A(n22523), .B(n22522), .Y(n37433) );
  OR2X1 U30345 ( .A(n29518), .B(n29517), .Y(n37434) );
  OR2X1 U30346 ( .A(n24355), .B(n24354), .Y(n37435) );
  OR2X1 U30347 ( .A(n23028), .B(n23027), .Y(n37436) );
  OR2X1 U30348 ( .A(n24162), .B(n24161), .Y(n37437) );
  OR2X1 U30349 ( .A(n24090), .B(n24089), .Y(n37438) );
  OR2X1 U30350 ( .A(n24080), .B(n24079), .Y(n37439) );
  OR2X1 U30351 ( .A(n24070), .B(n24069), .Y(n37440) );
  OR2X1 U30352 ( .A(n20865), .B(n20864), .Y(n37441) );
  OR2X1 U30353 ( .A(n20876), .B(n20874), .Y(n37442) );
  OR2X1 U30354 ( .A(n20855), .B(n20854), .Y(n37443) );
  OR2X1 U30355 ( .A(n20887), .B(n20886), .Y(n37444) );
  OR2X1 U30356 ( .A(n21699), .B(n21698), .Y(n37445) );
  OR2X1 U30357 ( .A(n24305), .B(n24304), .Y(n37446) );
  OR2X1 U30358 ( .A(n24345), .B(n24344), .Y(n37447) );
  OR2X1 U30359 ( .A(n24619), .B(n24618), .Y(n37448) );
  OR2X1 U30360 ( .A(n24265), .B(n24264), .Y(n37449) );
  OR2X1 U30361 ( .A(n24407), .B(n24406), .Y(n37450) );
  OR2X1 U30362 ( .A(n30240), .B(n30239), .Y(n37451) );
  OR2X1 U30363 ( .A(n29608), .B(n29607), .Y(n37452) );
  OR2X1 U30364 ( .A(n24437), .B(n24436), .Y(n37453) );
  OR2X1 U30365 ( .A(n24447), .B(n24446), .Y(n37454) );
  OR2X1 U30366 ( .A(n24569), .B(n24568), .Y(n37455) );
  OR2X1 U30367 ( .A(n24599), .B(n24598), .Y(n37456) );
  OR2X1 U30368 ( .A(n24589), .B(n24588), .Y(n37457) );
  OR2X1 U30369 ( .A(n24365), .B(n24364), .Y(n37458) );
  OR2X1 U30370 ( .A(n24417), .B(n24416), .Y(n37459) );
  OR2X1 U30371 ( .A(n24457), .B(n24456), .Y(n37460) );
  OR2X1 U30372 ( .A(n29819), .B(n29818), .Y(n37461) );
  OR2X1 U30373 ( .A(n29789), .B(n29788), .Y(n37462) );
  OR2X1 U30374 ( .A(n29849), .B(n29848), .Y(n37463) );
  OR2X1 U30375 ( .A(n24325), .B(n24324), .Y(n37464) );
  OR2X1 U30376 ( .A(n29729), .B(n29728), .Y(n37465) );
  XOR2X1 U30377 ( .A(n33266), .B(n42559), .Y(n37466) );
  NAND4X1 U30378 ( .A(n43222), .B(n43221), .C(n43220), .D(n43219), .Y(n12493)
         );
  NAND4X1 U30379 ( .A(n44059), .B(n44058), .C(n44057), .D(n44056), .Y(
        net209589) );
  CLKINVX1 U30380 ( .A(net209589), .Y(net209570) );
  OR2X1 U30381 ( .A(n24020), .B(n24019), .Y(n37467) );
  NAND2X1 U30382 ( .A(n37338), .B(net216265), .Y(n11933) );
  NAND4X1 U30383 ( .A(n43302), .B(n43301), .C(n43300), .D(n43299), .Y(n11668)
         );
  CLKINVX1 U30384 ( .A(n11668), .Y(net209479) );
  AND3X2 U30385 ( .A(net209927), .B(net209884), .C(net209893), .Y(n37469) );
  NAND4X1 U30386 ( .A(n44132), .B(n44131), .C(n44130), .D(n44129), .Y(
        net209868) );
  CLKINVX1 U30387 ( .A(net209868), .Y(net209885) );
  AND2X2 U30388 ( .A(n39745), .B(n39746), .Y(n37470) );
  AND2X2 U30389 ( .A(n40635), .B(net171523), .Y(n37471) );
  NAND4X1 U30390 ( .A(n47040), .B(n47039), .C(n47038), .D(n47037), .Y(n11132)
         );
  AND2X2 U30391 ( .A(n41149), .B(net213535), .Y(n37472) );
  AND2X2 U30392 ( .A(n40955), .B(net214991), .Y(n37473) );
  AND2X2 U30393 ( .A(n41015), .B(net215135), .Y(n37474) );
  OA21XL U30394 ( .A0(n39644), .A1(n39647), .B0(n39894), .Y(n37475) );
  CLKINVX1 U30395 ( .A(n12796), .Y(net171313) );
  CLKINVX1 U30396 ( .A(n11607), .Y(n_cell_301249_net269488) );
  CLKINVX1 U30397 ( .A(n12887), .Y(n39626) );
  NAND4X1 U30398 ( .A(n43744), .B(n43743), .C(n43742), .D(n43741), .Y(n11693)
         );
  NAND4X1 U30399 ( .A(n43280), .B(n43279), .C(n43278), .D(n43277), .Y(n12686)
         );
  CLKINVX1 U30400 ( .A(n12686), .Y(n39557) );
  CLKINVX1 U30401 ( .A(n11977), .Y(n39289) );
  XOR2X1 U30402 ( .A(n32442), .B(n36736), .Y(n37476) );
  XOR2X1 U30403 ( .A(n36734), .B(n32546), .Y(n37477) );
  XOR2X1 U30404 ( .A(n36734), .B(n32506), .Y(n37478) );
  XOR2X1 U30405 ( .A(n36733), .B(n32498), .Y(n37479) );
  XOR2X1 U30406 ( .A(n36735), .B(n32530), .Y(n37480) );
  XOR2X1 U30407 ( .A(n36735), .B(n32426), .Y(n37481) );
  XOR2X1 U30408 ( .A(n36734), .B(n32762), .Y(n37482) );
  XOR2X1 U30409 ( .A(n36736), .B(n32538), .Y(n37483) );
  XOR2X1 U30410 ( .A(n36734), .B(n32490), .Y(n37484) );
  XOR2X1 U30411 ( .A(n36735), .B(n32978), .Y(n37485) );
  NAND4X1 U30412 ( .A(n46039), .B(n46038), .C(n46037), .D(n46036), .Y(n12390)
         );
  CLKINVX1 U30413 ( .A(n12390), .Y(n39487) );
  XOR2X1 U30414 ( .A(n36749), .B(n32716), .Y(n37486) );
  XOR2X1 U30415 ( .A(n32449), .B(n36771), .Y(n37487) );
  NAND4BX2 U30416 ( .AN(n37306), .B(net216597), .C(net216594), .D(net216595),
        .Y(n10341) );
  OR4X1 U30417 ( .A(n20073), .B(n20072), .C(n20071), .D(n20070), .Y(n37488) );
  OR4X1 U30418 ( .A(n20504), .B(n20503), .C(n20502), .D(n20501), .Y(n37489) );
  XOR2X1 U30419 ( .A(n36736), .B(n32778), .Y(n37490) );
  XOR2X1 U30420 ( .A(n36771), .B(n32577), .Y(n37491) );
  XOR2X1 U30421 ( .A(n36771), .B(n32641), .Y(n37492) );
  OR2X1 U30422 ( .A(n23331), .B(n23330), .Y(n37493) );
  OR2X1 U30423 ( .A(n23626), .B(n23625), .Y(n37494) );
  OR2X1 U30424 ( .A(n23666), .B(n23665), .Y(n37495) );
  OR2X1 U30425 ( .A(n23656), .B(n23655), .Y(n37496) );
  OR2X1 U30426 ( .A(n24517), .B(n24516), .Y(n37497) );
  OR2X1 U30427 ( .A(n24315), .B(n24314), .Y(n37498) );
  OR2X1 U30428 ( .A(n24507), .B(n24506), .Y(n37499) );
  OR2X1 U30429 ( .A(n24537), .B(n24536), .Y(n37500) );
  OR2X1 U30430 ( .A(n24579), .B(n24578), .Y(n37501) );
  OR2X1 U30431 ( .A(n24559), .B(n24557), .Y(n37502) );
  OR2X1 U30432 ( .A(n24295), .B(n24294), .Y(n37503) );
  OR2X1 U30433 ( .A(n24375), .B(n24374), .Y(n37504) );
  OR2X1 U30434 ( .A(n24497), .B(n24496), .Y(n37505) );
  OR2X1 U30435 ( .A(n24467), .B(n24466), .Y(n37506) );
  OR2X1 U30436 ( .A(n24487), .B(n24486), .Y(n37507) );
  OR2X1 U30437 ( .A(n24477), .B(n24476), .Y(n37508) );
  AND2X2 U30438 ( .A(net212214), .B(net209924), .Y(n37509) );
  NAND2BX1 U30439 ( .AN(n39356), .B(net211256), .Y(n10710) );
  CLKINVX1 U30440 ( .A(n10710), .Y(net210238) );
  NAND2BX1 U30441 ( .AN(n39376), .B(net211641), .Y(n10753) );
  CLKINVX1 U30442 ( .A(n10753), .Y(net151737) );
  NAND2BX1 U30443 ( .AN(n39382), .B(net211992), .Y(n10756) );
  CLKINVX1 U30444 ( .A(n10756), .Y(net151481) );
  NAND2X1 U30445 ( .A(n12329), .B(n12324), .Y(n10861) );
  CLKINVX1 U30446 ( .A(n10861), .Y(net151599) );
  NAND2BX1 U30447 ( .AN(n39370), .B(net210772), .Y(net210526) );
  NAND2BX1 U30448 ( .AN(n39367), .B(net211513), .Y(n10733) );
  NAND2BX1 U30449 ( .AN(n39412), .B(net213362), .Y(n10879) );
  NAND2BX1 U30450 ( .AN(n39379), .B(net211348), .Y(n10689) );
  CLKINVX1 U30451 ( .A(n10689), .Y(net171548) );
  OR2X1 U30452 ( .A(n36945), .B(net259841), .Y(n37510) );
  OA21XL U30453 ( .A0(n39567), .A1(n39568), .B0(n39791), .Y(n37511) );
  NAND2X1 U30454 ( .A(net210148), .B(net210234), .Y(n10040) );
  NAND2BX1 U30455 ( .AN(net210673), .B(n36947), .Y(net210481) );
  OA21XL U30456 ( .A0(n39533), .A1(n10219), .B0(net151557), .Y(n37512) );
  OR2X1 U30457 ( .A(n39498), .B(net210543), .Y(n37513) );
  NAND2X1 U30458 ( .A(n37237), .B(net210702), .Y(net209287) );
  CLKINVX1 U30459 ( .A(net209287), .Y(net209302) );
  OR2X1 U30460 ( .A(net210544), .B(n39946), .Y(n37514) );
  NAND3X1 U30461 ( .A(n39337), .B(net216817), .C(net216814), .Y(n10504) );
  NAND2BX1 U30462 ( .AN(n39390), .B(net212901), .Y(n10274) );
  CLKINVX1 U30463 ( .A(n10274), .Y(n39987) );
  CLKINVX1 U30464 ( .A(n11985), .Y(net209760) );
  NAND2X1 U30465 ( .A(n40788), .B(net216490), .Y(n11959) );
  NAND2BX1 U30466 ( .AN(n39387), .B(net212866), .Y(n10807) );
  NAND2BX1 U30467 ( .AN(n_cell_301249_net267822), .B(net213603), .Y(n10939) );
  CLKINVX1 U30468 ( .A(n10939), .Y(n_cell_301249_net269836) );
  NAND4BBX1 U30469 ( .AN(n37006), .BN(n37307), .C(net215095), .D(net215093),
        .Y(n11576) );
  CLKINVX1 U30470 ( .A(n11576), .Y(n39701) );
  NAND3X1 U30471 ( .A(net216497), .B(net216498), .C(n40786), .Y(n11622) );
  CLKINVX1 U30472 ( .A(n11622), .Y(n39702) );
  OR2X1 U30473 ( .A(net171105), .B(net171103), .Y(n37515) );
  NAND2BX1 U30474 ( .AN(n_cell_301249_net267885), .B(net212094), .Y(n10760) );
  CLKINVX1 U30475 ( .A(n10760), .Y(n39927) );
  NAND2BX1 U30476 ( .AN(n_cell_301249_net267840), .B(net212099), .Y(n10761) );
  CLKINVX1 U30477 ( .A(n10761), .Y(n39929) );
  NAND2BX1 U30478 ( .AN(n_cell_301249_net266944), .B(net212831), .Y(n10905) );
  CLKINVX1 U30479 ( .A(n10905), .Y(n39991) );
  NAND3X1 U30480 ( .A(net216403), .B(net216400), .C(n_cell_301249_net267165),
        .Y(n10487) );
  NAND2X1 U30481 ( .A(n40797), .B(net212124), .Y(n11272) );
  CLKINVX1 U30482 ( .A(n11272), .Y(net151550) );
  NAND2BX1 U30483 ( .AN(n_cell_301249_net267490), .B(net212119), .Y(n10646) );
  CLKINVX1 U30484 ( .A(n10646), .Y(n39923) );
  NAND4BX1 U30485 ( .AN(n37219), .B(net215369), .C(net215366), .D(net215367),
        .Y(n10382) );
  NAND2BX1 U30486 ( .AN(n40436), .B(net210353), .Y(n12834) );
  NAND2X1 U30487 ( .A(n39391), .B(net212911), .Y(n10273) );
  CLKINVX1 U30488 ( .A(n10273), .Y(net209155) );
  NAND2BX1 U30489 ( .AN(n_cell_301249_net267855), .B(net211618), .Y(n10638) );
  CLKINVX1 U30490 ( .A(n10638), .Y(n_cell_303546_net277804) );
  NAND2BX1 U30491 ( .AN(n_cell_301249_net266916), .B(net216868), .Y(n10502) );
  CLKINVX1 U30492 ( .A(n10502), .Y(net209746) );
  NAND2BX1 U30493 ( .AN(n_cell_301249_net267409), .B(net212129), .Y(n11274) );
  CLKINVX1 U30494 ( .A(n11274), .Y(n39621) );
  NAND2X1 U30495 ( .A(n37340), .B(net215078), .Y(n12807) );
  CLKINVX1 U30496 ( .A(n12807), .Y(n39550) );
  NAND2BX1 U30497 ( .AN(n_cell_301249_net268223), .B(net211443), .Y(n10626) );
  CLKINVX1 U30498 ( .A(n10626), .Y(n39934) );
  NAND2BX1 U30499 ( .AN(n_cell_301249_net267225), .B(net211778), .Y(n10657) );
  NAND2BX1 U30500 ( .AN(n_cell_301249_net268103), .B(net211591), .Y(n10631) );
  CLKINVX1 U30501 ( .A(n10631), .Y(n_cell_303546_net277822) );
  NAND2BX1 U30502 ( .AN(n_cell_301249_net268166), .B(net211433), .Y(n10624) );
  CLKINVX1 U30503 ( .A(n10624), .Y(n_cell_301249_net269755) );
  NAND2BX1 U30504 ( .AN(n40790), .B(net213542), .Y(n10982) );
  NAND2BX1 U30505 ( .AN(n_cell_301249_net267213), .B(net211768), .Y(n10659) );
  CLKINVX1 U30506 ( .A(n10659), .Y(n_cell_303546_net277772) );
  NAND2BX1 U30507 ( .AN(n_cell_301249_net267207), .B(net211773), .Y(n10658) );
  CLKINVX1 U30508 ( .A(n10658), .Y(n_cell_301249_net269701) );
  NAND2BX1 U30509 ( .AN(n40429), .B(net212053), .Y(net210007) );
  INVX3 U30510 ( .A(net210007), .Y(net171528) );
  NAND3X1 U30511 ( .A(net216358), .B(net216355), .C(n_cell_301249_net267308),
        .Y(n11942) );
  NAND2BX1 U30512 ( .AN(n39389), .B(net212906), .Y(n10272) );
  CLKINVX1 U30513 ( .A(n10272), .Y(net171474) );
  NAND2BX1 U30514 ( .AN(n40789), .B(net216499), .Y(n11958) );
  CLKINVX1 U30515 ( .A(n11958), .Y(n39556) );
  NAND2BX1 U30516 ( .AN(n_cell_301249_net267646), .B(net212043), .Y(n11262) );
  CLKINVX1 U30517 ( .A(n11262), .Y(net171530) );
  NAND2BX1 U30518 ( .AN(n40423), .B(net212078), .Y(n12212) );
  INVX3 U30519 ( .A(n12212), .Y(net151586) );
  NAND2BX1 U30520 ( .AN(n_cell_301249_net267343), .B(net212144), .Y(n12856) );
  CLKINVX1 U30521 ( .A(n12856), .Y(n_cell_301249_net269714) );
  NAND2BX1 U30522 ( .AN(n_cell_301249_net267349), .B(net212159), .Y(n11281) );
  CLKINVX1 U30523 ( .A(n11281), .Y(net171525) );
  NAND2BX1 U30524 ( .AN(n_cell_301249_net267269), .B(net212169), .Y(n11283) );
  CLKINVX1 U30525 ( .A(n11283), .Y(n39623) );
  NAND2X1 U30526 ( .A(n12671), .B(n12668), .Y(n10518) );
  NAND2BX1 U30527 ( .AN(n_cell_301249_net267694), .B(net214678), .Y(n10470) );
  CLKINVX1 U30528 ( .A(n10470), .Y(n39833) );
  NAND2BX1 U30529 ( .AN(n_cell_301249_net267574), .B(net212017), .Y(n11265) );
  NAND2BX1 U30530 ( .AN(n40420), .B(net212022), .Y(n12221) );
  CLKINVX1 U30531 ( .A(n12221), .Y(net151571) );
  NAND2BX1 U30532 ( .AN(n40442), .B(net213582), .Y(net209099) );
  CLKINVX1 U30533 ( .A(net209099), .Y(net171392) );
  NAND2BX1 U30534 ( .AN(n_cell_301249_net268355), .B(net211167), .Y(n10613) );
  CLKINVX1 U30535 ( .A(n10613), .Y(n_cell_301249_net269763) );
  NAND2BX1 U30536 ( .AN(n_cell_301249_net268172), .B(net211448), .Y(n10622) );
  CLKINVX1 U30537 ( .A(n10622), .Y(n39935) );
  NAND4BX1 U30538 ( .AN(n37303), .B(net215315), .C(net215312), .D(net215313),
        .Y(n10424) );
  NAND2BX1 U30539 ( .AN(n_cell_301249_net268044), .B(net211579), .Y(n10629) );
  CLKINVX1 U30540 ( .A(n10629), .Y(n_cell_301249_net269746) );
  NAND2BX1 U30541 ( .AN(n39296), .B(net215213), .Y(n10555) );
  NAND2BX1 U30542 ( .AN(n40417), .B(net213477), .Y(net209124) );
  CLKINVX1 U30543 ( .A(net209124), .Y(net171408) );
  NAND2BX1 U30544 ( .AN(n40445), .B(net211603), .Y(net209992) );
  NAND2BX1 U30545 ( .AN(n_cell_301249_net267415), .B(net212134), .Y(n11273) );
  CLKINVX1 U30546 ( .A(n11273), .Y(n39622) );
  NAND2BX1 U30547 ( .AN(n_cell_301249_net267257), .B(net213557), .Y(n10974) );
  NAND2BX1 U30548 ( .AN(n40454), .B(net211463), .Y(n13026) );
  CLKINVX1 U30549 ( .A(n13026), .Y(n39619) );
  NAND3X1 U30550 ( .A(net215433), .B(net215434), .C(n39302), .Y(n10585) );
  CLKINVX1 U30551 ( .A(n10585), .Y(net171234) );
  NAND3X1 U30552 ( .A(n11054), .B(n11057), .C(n39397), .Y(n10239) );
  NAND2BX1 U30553 ( .AN(n40416), .B(net212048), .Y(n12219) );
  CLKINVX1 U30554 ( .A(n12219), .Y(net151566) );
  NAND2BX1 U30555 ( .AN(n39336), .B(net216805), .Y(n10505) );
  NAND2BX1 U30556 ( .AN(n39327), .B(net215903), .Y(n10530) );
  OR2X1 U30557 ( .A(net209753), .B(n40970), .Y(n37516) );
  AO21X1 U30558 ( .A0(n41094), .A1(n11521), .B0(n41096), .Y(n37517) );
  AO21X1 U30559 ( .A0(n_cell_301249_net269746), .A1(n10630), .B0(n40717), .Y(
        n37518) );
  CLKINVX1 U30560 ( .A(n11932), .Y(n39552) );
  CLKINVX1 U30561 ( .A(n12392), .Y(n_cell_303546_net277738) );
  CLKINVX1 U30562 ( .A(n10806), .Y(net171477) );
  NAND2BX2 U30563 ( .AN(n39388), .B(net212871), .Y(n10806) );
  OR2X1 U30564 ( .A(n9999), .B(net171530), .Y(n37519) );
  CLKINVX1 U30565 ( .A(n11934), .Y(n_cell_301249_net269571) );
  CLKINVX1 U30566 ( .A(n12166), .Y(n_cell_301249_net269583) );
  CLKINVX1 U30567 ( .A(n12803), .Y(n_cell_301249_net269568) );
  CLKINVX1 U30568 ( .A(n_cell_303546_net275934), .Y(net151283) );
  CLKINVX1 U30569 ( .A(n10904), .Y(n39532) );
  CLKINVX1 U30570 ( .A(n12186), .Y(net151767) );
  CLKINVX1 U30571 ( .A(n_cell_303546_net276178), .Y(n39551) );
  CLKINVX1 U30572 ( .A(n11994), .Y(net209768) );
  CLKINVX1 U30573 ( .A(n10205), .Y(net171414) );
  CLKINVX1 U30574 ( .A(n_cell_303546_net275923), .Y(n_cell_301249_net269797)
         );
  INVX3 U30575 ( .A(n10906), .Y(net171480) );
  CLKINVX1 U30576 ( .A(n10501), .Y(net171108) );
  CLKINVX1 U30577 ( .A(n_cell_303546_net276009), .Y(n_cell_301249_net269711)
         );
  CLKINVX1 U30578 ( .A(n10801), .Y(net151532) );
  CLKINVX1 U30579 ( .A(n11519), .Y(net210034) );
  CLKBUFX3 U30580 ( .A(n11954), .Y(net260247) );
  CLKBUFX3 U30581 ( .A(n10426), .Y(net259641) );
  NAND2X1 U30582 ( .A(n19412), .B(n41796), .Y(n19292) );
  NOR2X2 U30583 ( .A(n19278), .B(n50145), .Y(n37520) );
  NAND2X1 U30584 ( .A(n19281), .B(n41796), .Y(n37525) );
  CLKINVX1 U30585 ( .A(n12591), .Y(n39699) );
  NAND3X1 U30586 ( .A(n40798), .B(net214777), .C(net214774), .Y(n11586) );
  INVX3 U30587 ( .A(n11586), .Y(net171315) );
  CLKINVX1 U30588 ( .A(n11613), .Y(net171158) );
  NAND3X1 U30589 ( .A(net216488), .B(net216489), .C(n40792), .Y(n11620) );
  CLKINVX1 U30590 ( .A(n11620), .Y(net151275) );
  NAND3X1 U30591 ( .A(net214984), .B(n40449), .C(net214985), .Y(n12408) );
  CLKINVX1 U30592 ( .A(n12408), .Y(net151380) );
  NAND2BX1 U30593 ( .AN(n_cell_301249_net267700), .B(net213623), .Y(n10946) );
  CLKINVX1 U30594 ( .A(n10946), .Y(n_cell_303546_net278017) );
  NAND2BX1 U30595 ( .AN(n_cell_301249_net267828), .B(net213613), .Y(n10938) );
  CLKINVX1 U30596 ( .A(n10938), .Y(n39482) );
  NAND2BX1 U30597 ( .AN(n_cell_301249_net268342), .B(net212557), .Y(net210556)
         );
  CLKINVX1 U30598 ( .A(net210556), .Y(n_cell_301249_net269853) );
  NAND2BX1 U30599 ( .AN(n_cell_301249_net268336), .B(net212552), .Y(net210555)
         );
  CLKINVX1 U30600 ( .A(net210555), .Y(n40001) );
  NAND2X1 U30601 ( .A(n37339), .B(net216256), .Y(n12167) );
  CLKINVX1 U30602 ( .A(n12167), .Y(n_cell_303546_net277942) );
  NAND2BX1 U30603 ( .AN(n_cell_301249_net267676), .B(net214672), .Y(n10469) );
  CLKINVX1 U30604 ( .A(n10469), .Y(n_cell_303546_net277936) );
  NAND2BX1 U30605 ( .AN(n_cell_301249_net267769), .B(net213608), .Y(n10940) );
  NAND2BX1 U30606 ( .AN(n_cell_301249_net267804), .B(net214688), .Y(n11915) );
  NAND2BX1 U30607 ( .AN(n_cell_301249_net268398), .B(net211187), .Y(n10614) );
  CLKINVX1 U30608 ( .A(n10614), .Y(n39937) );
  NAND3X1 U30609 ( .A(net214960), .B(net214958), .C(n_cell_301249_net267980),
        .Y(n10292) );
  CLKINVX1 U30610 ( .A(n10292), .Y(n_cell_301249_net269650) );
  NAND2BX1 U30611 ( .AN(n_cell_301249_net268380), .B(net213312), .Y(n10762) );
  CLKINVX1 U30612 ( .A(n10762), .Y(n40003) );
  NAND2BX1 U30613 ( .AN(n_cell_301249_net268386), .B(net212562), .Y(n10763) );
  CLKINVX1 U30614 ( .A(n10763), .Y(n40002) );
  NAND2BX1 U30615 ( .AN(n40421), .B(n_cell_301249_net267510), .Y(n11595) );
  CLKINVX1 U30616 ( .A(n11595), .Y(n_cell_301249_net269941) );
  NAND2X1 U30617 ( .A(n12449), .B(n12453), .Y(n10080) );
  CLKINVX1 U30618 ( .A(n10080), .Y(n_cell_301249_net269615) );
  NAND2BX1 U30619 ( .AN(n_cell_301249_net268217), .B(net211438), .Y(n10625) );
  CLKINVX1 U30620 ( .A(n10625), .Y(n_cell_301249_net269758) );
  NAND2BX1 U30621 ( .AN(n40460), .B(net211563), .Y(net209976) );
  CLKINVX1 U30622 ( .A(net209976), .Y(net171545) );
  NAND2BX1 U30623 ( .AN(n40451), .B(net215096), .Y(net209689) );
  CLKINVX1 U30624 ( .A(net209689), .Y(net171274) );
  NAND3X1 U30625 ( .A(net216191), .B(net216189), .C(n40427), .Y(n11870) );
  CLKINVX1 U30626 ( .A(n11870), .Y(net151304) );
  NAND2BX1 U30627 ( .AN(n40453), .B(net213220), .Y(n12604) );
  CLKINVX1 U30628 ( .A(n12604), .Y(net151786) );
  NAND2BX1 U30629 ( .AN(n40419), .B(n_cell_301249_net267516), .Y(n11594) );
  CLKINVX1 U30630 ( .A(n11594), .Y(n_cell_301249_net269943) );
  AND2X2 U30631 ( .A(net265207), .B(n51444), .Y(n37526) );
  CLKINVX1 U30632 ( .A(n11917), .Y(n_cell_303546_net277852) );
  AO21X1 U30633 ( .A0(n41183), .A1(n11228), .B0(n41184), .Y(n37527) );
  AND3X2 U30634 ( .A(net259641), .B(net259645), .C(n_cell_301249_net269950),
        .Y(n37528) );
  CLKINVX1 U30635 ( .A(n10927), .Y(n_cell_303546_net277759) );
  OR2X1 U30636 ( .A(n37336), .B(n_cell_301249_net267810), .Y(n10464) );
  CLKINVX1 U30637 ( .A(n10464), .Y(n_cell_301249_net269596) );
  OR2X1 U30638 ( .A(n10295), .B(net171280), .Y(n37529) );
  BUFX4 U30639 ( .A(net221956), .Y(net266780) );
  CLKINVX1 U30640 ( .A(n_cell_303546_net275987), .Y(n_cell_303546_net277834)
         );
  CLKBUFX3 U30641 ( .A(n12415), .Y(net260352) );
  CLKINVX1 U30642 ( .A(net260352), .Y(net151374) );
  CLKINVX1 U30643 ( .A(n39444), .Y(n_cell_303546_net277667) );
  CLKINVX1 U30644 ( .A(n10447), .Y(net171259) );
  CLKINVX1 U30645 ( .A(net209974), .Y(net171544) );
  NAND2X1 U30646 ( .A(n19523), .B(n41796), .Y(n19420) );
  NOR2X2 U30647 ( .A(n19335), .B(n50145), .Y(n37530) );
  NAND4X1 U30648 ( .A(net215148), .B(net215146), .C(net215147), .D(net215149),
        .Y(n11551) );
  CLKINVX1 U30649 ( .A(n11551), .Y(n39698) );
  NAND4X1 U30650 ( .A(net214735), .B(net214736), .C(net214737), .D(net214738),
        .Y(n11537) );
  NAND4X1 U30651 ( .A(net215203), .B(net215202), .C(net215200), .D(net215201),
        .Y(n11538) );
  NAND4X1 U30652 ( .A(net215164), .B(net215165), .C(net215166), .D(net215167),
        .Y(n11542) );
  CLKINVX1 U30653 ( .A(n11542), .Y(n_cell_303546_net277506) );
  CLKBUFX3 U30654 ( .A(n34136), .Y(n42058) );
  CLKBUFX3 U30655 ( .A(n34137), .Y(n42060) );
  CLKBUFX3 U30656 ( .A(n34129), .Y(n42061) );
  CLKBUFX3 U30657 ( .A(n34132), .Y(n41799) );
  CLKBUFX3 U30658 ( .A(n34141), .Y(n41801) );
  CLKBUFX3 U30659 ( .A(n34133), .Y(n41802) );
  CLKBUFX3 U30660 ( .A(n34142), .Y(n41804) );
  CLKBUFX3 U30661 ( .A(n34134), .Y(n41805) );
  CLKBUFX3 U30662 ( .A(n34413), .Y(n41800) );
  CLKBUFX3 U30663 ( .A(n34414), .Y(n41803) );
  CLKBUFX3 U30664 ( .A(n34416), .Y(n42057) );
  CLKBUFX3 U30665 ( .A(n34409), .Y(n42059) );
  CLKBUFX3 U30666 ( .A(n34410), .Y(n42062) );
  CLKBUFX3 U30667 ( .A(n34412), .Y(n41798) );
  NAND2X1 U30668 ( .A(n39731), .B(n11725), .Y(n39730) );
  AOI211X1 U30669 ( .A0(n11725), .A1(n11726), .B0(net209509), .C0(net151394),
        .Y(n11719) );
  NOR2X1 U30670 ( .A(n49502), .B(n49504), .Y(n11725) );
  NOR2X1 U30671 ( .A(n11149), .B(n47292), .Y(net211147) );
  XOR2X1 U30672 ( .A(n36746), .B(n34076), .Y(n47292) );
  NOR2X1 U30673 ( .A(n12751), .B(n45660), .Y(n45664) );
  XOR2X1 U30674 ( .A(n34017), .B(n36779), .Y(n45660) );
  NOR2X1 U30675 ( .A(n12089), .B(n45670), .Y(n45674) );
  XOR2X1 U30676 ( .A(n34041), .B(n36786), .Y(n45670) );
  NOR2X1 U30677 ( .A(n12747), .B(n45655), .Y(n45659) );
  XOR2X1 U30678 ( .A(n34009), .B(n36780), .Y(n45655) );
  XOR2X1 U30679 ( .A(n34033), .B(n36782), .Y(n45680) );
  NOR4X1 U30680 ( .A(n44148), .B(n44147), .C(n44146), .D(n44145), .Y(n44149)
         );
  XOR2X1 U30681 ( .A(n42090), .B(n36879), .Y(n44146) );
  XOR2X1 U30682 ( .A(n41813), .B(n42515), .Y(n44984) );
  XOR2X1 U30683 ( .A(n41825), .B(n42518), .Y(n44873) );
  NOR2X1 U30684 ( .A(n45336), .B(net209603), .Y(n45346) );
  XOR2X1 U30685 ( .A(n41824), .B(n42523), .Y(n45336) );
  NOR2X1 U30686 ( .A(n46522), .B(net210695), .Y(n46532) );
  XOR2X1 U30687 ( .A(n41317), .B(n41816), .Y(n46522) );
  XOR2X1 U30688 ( .A(n36754), .B(n41816), .Y(n47579) );
  NOR2X1 U30689 ( .A(n46343), .B(net209900), .Y(n46353) );
  XOR2X1 U30690 ( .A(n41316), .B(n41817), .Y(n46343) );
  NOR2X1 U30691 ( .A(n46221), .B(n48182), .Y(n46231) );
  XOR2X1 U30692 ( .A(n41316), .B(n41838), .Y(n46221) );
  NOR2X1 U30693 ( .A(n46390), .B(n48172), .Y(n46400) );
  XOR2X1 U30694 ( .A(n41313), .B(n41830), .Y(n46390) );
  XOR2X1 U30695 ( .A(n41313), .B(n41814), .Y(n46533) );
  INVX3 U30696 ( .A(n41308), .Y(n41313) );
  XOR2X1 U30697 ( .A(n41318), .B(n41822), .Y(n46365) );
  XOR2X1 U30698 ( .A(n41312), .B(n41825), .Y(n46456) );
  XOR2X1 U30699 ( .A(n41309), .B(n41813), .Y(n46489) );
  XOR2X1 U30700 ( .A(n41310), .B(n41833), .Y(n46232) );
  INVX3 U30701 ( .A(n41308), .Y(n41310) );
  XOR2X1 U30702 ( .A(n41312), .B(n41821), .Y(n46354) );
  INVX3 U30703 ( .A(n41315), .Y(n41312) );
  XOR2X1 U30704 ( .A(n36760), .B(n41820), .Y(n47325) );
  XOR2X1 U30705 ( .A(n36764), .B(n34089), .Y(n47286) );
  NOR2X1 U30706 ( .A(n46189), .B(n48133), .Y(n46193) );
  XOR2X1 U30707 ( .A(n34081), .B(n36780), .Y(n46189) );
  NAND3X1 U30708 ( .A(n11066), .B(n11065), .C(n11064), .Y(n10829) );
  AND2X2 U30709 ( .A(n48522), .B(n48521), .Y(n11064) );
  OR4X1 U30710 ( .A(net151491), .B(net151494), .C(net171459), .D(net171460),
        .Y(n39525) );
  OAI21XL U30711 ( .A0(net171459), .A1(n48539), .B0(n11024), .Y(n48540) );
  CLKINVX1 U30712 ( .A(n11023), .Y(net171459) );
  NAND3X1 U30713 ( .A(n12323), .B(n12385), .C(n11118), .Y(n10254) );
  AOI211X1 U30714 ( .A0(n11119), .A1(n11118), .B0(net171491), .C0(net171490),
        .Y(n11112) );
  AND2X2 U30715 ( .A(n12322), .B(n12326), .Y(n11118) );
  AND2X2 U30716 ( .A(n12915), .B(n12918), .Y(n11352) );
  CLKINVX1 U30717 ( .A(n10506), .Y(net171111) );
  CLKINVX1 U30718 ( .A(net213666), .Y(net210462) );
  OAI21XL U30719 ( .A0(net213666), .A1(n39714), .B0(n39842), .Y(n39717) );
  NAND4BX1 U30720 ( .AN(n48291), .B(n48293), .C(n48337), .D(n48335), .Y(
        net213666) );
  NAND2XL U30721 ( .A(net217946), .B(n49516), .Y(n48867) );
  XNOR2XL U30722 ( .A(n49516), .B(n42627), .Y(n27720) );
  NAND2BX1 U30723 ( .AN(net210417), .B(n40030), .Y(n40031) );
  CLKINVX1 U30724 ( .A(net210417), .Y(net210517) );
  OR2X1 U30725 ( .A(n47759), .B(n47771), .Y(net210417) );
  CLKINVX1 U30726 ( .A(net258320), .Y(n41196) );
  XOR2X1 U30727 ( .A(n9661), .B(n42592), .Y(n45236) );
  XOR2X1 U30728 ( .A(n9661), .B(net219468), .Y(n45267) );
  XOR2X1 U30729 ( .A(n9663), .B(n36893), .Y(n45272) );
  XNOR2X1 U30730 ( .A(n51200), .B(n41281), .Y(n29321) );
  XOR2X1 U30731 ( .A(n34429), .B(n42549), .Y(n45230) );
  XOR2X1 U30732 ( .A(n34430), .B(net219330), .Y(n45037) );
  XOR2X1 U30733 ( .A(n34430), .B(n42615), .Y(n45258) );
  XOR2X1 U30734 ( .A(n34432), .B(n34450), .Y(n45260) );
  XOR2X1 U30735 ( .A(n34432), .B(n36730), .Y(n45229) );
  XOR2X1 U30736 ( .A(n34426), .B(n41630), .Y(n45234) );
  XNOR2X1 U30737 ( .A(n50718), .B(n36856), .Y(n23125) );
  XNOR2X1 U30738 ( .A(n50939), .B(n36870), .Y(n28208) );
  XNOR2X1 U30739 ( .A(n50985), .B(n36870), .Y(n29350) );
  XNOR2X1 U30740 ( .A(n51223), .B(n42547), .Y(n27680) );
  XNOR2X1 U30741 ( .A(n50942), .B(net219310), .Y(n28148) );
  XNOR2X1 U30742 ( .A(n50977), .B(net219330), .Y(n29109) );
  XNOR2X1 U30743 ( .A(n50995), .B(net219310), .Y(n27185) );
  XOR2X1 U30744 ( .A(n41305), .B(n33692), .Y(n45638) );
  OA22XL U30745 ( .A0(net261924), .A1(n33684), .B0(n33692), .B1(n40147), .Y(
        n17029) );
  OA22XL U30746 ( .A0(net262741), .A1(n33940), .B0(n33948), .B1(n40108), .Y(
        n17797) );
  OA22XL U30747 ( .A0(net263216), .A1(n32466), .B0(n32474), .B1(n40083), .Y(
        n13375) );
  OA22XL U30748 ( .A0(net263805), .A1(n32930), .B0(n32938), .B1(n40050), .Y(
        n14767) );
  OA22XL U30749 ( .A0(net263748), .A1(n32978), .B0(n32986), .B1(n40053), .Y(
        n14911) );
  OA22XL U30750 ( .A0(net263767), .A1(n32956), .B0(n32964), .B1(n40052), .Y(
        n14845) );
  OA22XL U30751 ( .A0(net218478), .A1(n32948), .B0(n32956), .B1(n40051), .Y(
        n14821) );
  OA22XL U30752 ( .A0(net263159), .A1(n32780), .B0(n32788), .B1(n40087), .Y(
        n14317) );
  OA22XL U30753 ( .A0(net263140), .A1(n32788), .B0(n32796), .B1(n40087), .Y(
        n14341) );
  OA22XL U30754 ( .A0(net262969), .A1(n32700), .B0(n32708), .B1(n40098), .Y(
        n14077) );
  OA22XL U30755 ( .A0(net262969), .A1(n32692), .B0(n32700), .B1(n40097), .Y(
        n14053) );
  OA22XL U30756 ( .A0(net263368), .A1(n32578), .B0(n32586), .B1(n40075), .Y(
        n13711) );
  OA22XL U30757 ( .A0(net263178), .A1(n32754), .B0(n32762), .B1(n40085), .Y(
        n14239) );
  OA22XL U30758 ( .A0(net263178), .A1(n32762), .B0(n32770), .B1(n40086), .Y(
        n14263) );
  OA22XL U30759 ( .A0(net218354), .A1(n32474), .B0(n32482), .B1(n40084), .Y(
        n13399) );
  OA22XL U30760 ( .A0(net218432), .A1(n32938), .B0(n32946), .B1(n40051), .Y(
        n14791) );
  OA22XL U30761 ( .A0(net263368), .A1(n32570), .B0(n32578), .B1(n40075), .Y(
        n13687) );
  OA22XL U30762 ( .A0(net218496), .A1(n32514), .B0(n32522), .B1(n40071), .Y(
        n13519) );
  OA22XL U30763 ( .A0(net218348), .A1(n32410), .B0(n32418), .B1(n40080), .Y(
        n13207) );
  OA22XL U30764 ( .A0(net218310), .A1(n32402), .B0(n32410), .B1(n40079), .Y(
        n13183) );
  XNOR2X1 U30765 ( .A(n50952), .B(net219310), .Y(n25200) );
  OA22XL U30766 ( .A0(net263083), .A1(n32850), .B0(n32858), .B1(n40091), .Y(
        n14527) );
  XOR2X1 U30767 ( .A(n41302), .B(n34068), .Y(n46194) );
  OA22XL U30768 ( .A0(net263216), .A1(n32468), .B0(n32476), .B1(n40083), .Y(
        n13381) );
  OA22XL U30769 ( .A0(net263406), .A1(n32532), .B0(n32540), .B1(n40072), .Y(
        n13573) );
  OA22XL U30770 ( .A0(net218494), .A1(n32524), .B0(n32532), .B1(n40072), .Y(
        n13549) );
  OA22XL U30771 ( .A0(net218320), .A1(n32404), .B0(n32412), .B1(n40079), .Y(
        n13189) );
  OA22XL U30772 ( .A0(net263216), .A1(n32460), .B0(n32468), .B1(n40083), .Y(
        n13357) );
  XNOR2X1 U30773 ( .A(n36837), .B(n34090), .Y(n46182) );
  OA22XL U30774 ( .A0(net262190), .A1(n33428), .B0(n33436), .B1(n40133), .Y(
        n16261) );
  OA22XL U30775 ( .A0(net263824), .A1(n32916), .B0(n32924), .B1(n40049), .Y(
        n14725) );
  OA22XL U30776 ( .A0(net263007), .A1(n32660), .B0(n32668), .B1(n40095), .Y(
        n13957) );
  OA22XL U30777 ( .A0(net262171), .A1(n33444), .B0(n33452), .B1(n40134), .Y(
        n16309) );
  OA22XL U30778 ( .A0(net262190), .A1(n33436), .B0(n33444), .B1(n40134), .Y(
        n16285) );
  OA22XL U30779 ( .A0(net262209), .A1(n33420), .B0(n33428), .B1(n40133), .Y(
        n16237) );
  OA22XL U30780 ( .A0(net263805), .A1(n32924), .B0(n32932), .B1(n40050), .Y(
        n14749) );
  OA22XL U30781 ( .A0(net263824), .A1(n32908), .B0(n32916), .B1(n40049), .Y(
        n14701) );
  OAI211XL U30782 ( .A0(n32916), .A1(n42964), .B0(n14677), .C0(n14678), .Y(
        n35065) );
  OA22XL U30783 ( .A0(net263007), .A1(n32668), .B0(n32676), .B1(n40096), .Y(
        n13981) );
  OAI211XL U30784 ( .A0(n32660), .A1(n42871), .B0(n13909), .C0(n13910), .Y(
        n34809) );
  OA22XL U30785 ( .A0(net263748), .A1(n32986), .B0(n32994), .B1(n40054), .Y(
        n14935) );
  OA22XL U30786 ( .A0(net263216), .A1(n32458), .B0(n32466), .B1(n40083), .Y(
        n13351) );
  OA22XL U30787 ( .A0(net263235), .A1(n32450), .B0(n32458), .B1(n40082), .Y(
        n13327) );
  OA22XL U30788 ( .A0(net263767), .A1(n32970), .B0(n32978), .B1(n40053), .Y(
        n14887) );
  OAI211XL U30789 ( .A0(n32466), .A1(n42899), .B0(n13327), .C0(n13328), .Y(
        n34615) );
  OA22XL U30790 ( .A0(net263805), .A1(n32922), .B0(n32930), .B1(n40050), .Y(
        n14743) );
  OA22XL U30791 ( .A0(net263824), .A1(n32914), .B0(n32922), .B1(n40049), .Y(
        n14719) );
  OAI211XL U30792 ( .A0(n32930), .A1(n42962), .B0(n14719), .C0(n14720), .Y(
        n35079) );
  OAI211XL U30793 ( .A0(n32938), .A1(n42961), .B0(n14743), .C0(n14744), .Y(
        n35087) );
  OAI211XL U30794 ( .A0(n32402), .A1(n42908), .B0(n13135), .C0(n13136), .Y(
        n34551) );
  OA22XL U30795 ( .A0(net218396), .A1(n33986), .B0(n33994), .B1(n40110), .Y(
        n17935) );
  OA22XL U30796 ( .A0(net263368), .A1(n33058), .B0(n33066), .B1(n40141), .Y(
        n15151) );
  XOR2X1 U30797 ( .A(n41299), .B(n33988), .Y(n45693) );
  XNOR2X1 U30798 ( .A(n36843), .B(n34098), .Y(n46198) );
  OA22XL U30799 ( .A0(net262950), .A1(n32706), .B0(n32714), .B1(n40098), .Y(
        n14095) );
  OAI211XL U30800 ( .A0(n32978), .A1(n42987), .B0(n14863), .C0(n14864), .Y(
        n35127) );
  OA22XL U30801 ( .A0(net263026), .A1(n32634), .B0(n32642), .B1(n40094), .Y(
        n13879) );
  OA22XL U30802 ( .A0(net262209), .A1(n33410), .B0(n33418), .B1(n40132), .Y(
        n16207) );
  OA22XL U30803 ( .A0(net262950), .A1(n32714), .B0(n32722), .B1(n40099), .Y(
        n14119) );
  OA22XL U30804 ( .A0(net218308), .A1(n32522), .B0(n32530), .B1(n40072), .Y(
        n13543) );
  OAI211XL U30805 ( .A0(n32514), .A1(n42924), .B0(n13471), .C0(n13472), .Y(
        n34663) );
  OAI211XL U30806 ( .A0(n32754), .A1(n42890), .B0(n14191), .C0(n14192), .Y(
        n34903) );
  OA22XL U30807 ( .A0(net263064), .A1(n32858), .B0(n32866), .B1(n40092), .Y(
        n14551) );
  OAI211XL U30808 ( .A0(n32850), .A1(n42973), .B0(n14479), .C0(n14480), .Y(
        n34999) );
  OAI211XL U30809 ( .A0(n32762), .A1(n42889), .B0(n14215), .C0(n14216), .Y(
        n34911) );
  OAI211XL U30810 ( .A0(n32770), .A1(n42888), .B0(n14239), .C0(n14240), .Y(
        n34919) );
  OA22XL U30811 ( .A0(net263026), .A1(n32642), .B0(n32650), .B1(n40094), .Y(
        n13903) );
  OAI211XL U30812 ( .A0(n32474), .A1(n42898), .B0(n13351), .C0(n13352), .Y(
        n34623) );
  OAI211XL U30813 ( .A0(n32482), .A1(n42897), .B0(n13375), .C0(n13376), .Y(
        n34631) );
  OAI211XL U30814 ( .A0(n32410), .A1(n42907), .B0(n13159), .C0(n13160), .Y(
        n34559) );
  OA22XL U30815 ( .A0(net263007), .A1(n32652), .B0(n32660), .B1(n40095), .Y(
        n13933) );
  OA22XL U30816 ( .A0(net262247), .A1(n33386), .B0(n33394), .B1(n40131), .Y(
        n16135) );
  XOR2X1 U30817 ( .A(n41305), .B(n33964), .Y(n47036) );
  OAI211XL U30818 ( .A0(n33436), .A1(n42793), .B0(n16237), .C0(n16238), .Y(
        n35585) );
  OA22XL U30819 ( .A0(net262722), .A1(n33948), .B0(n33956), .B1(n40085), .Y(
        n17821) );
  OAI211XL U30820 ( .A0(n33538), .A1(n42746), .B0(n16543), .C0(n16544), .Y(
        n35687) );
  OAI211XL U30821 ( .A0(n32418), .A1(n42906), .B0(n13183), .C0(n13184), .Y(
        n34567) );
  XNOR2X1 U30822 ( .A(n36841), .B(n33498), .Y(n45811) );
  OAI211XL U30823 ( .A0(n32700), .A1(n42866), .B0(n14029), .C0(n14030), .Y(
        n34849) );
  OAI211XL U30824 ( .A0(n32692), .A1(n42867), .B0(n14005), .C0(n14006), .Y(
        n34841) );
  OAI211XL U30825 ( .A0(n32412), .A1(n42907), .B0(n13165), .C0(n13166), .Y(
        n34561) );
  OAI211XL U30826 ( .A0(n33410), .A1(n42797), .B0(n16159), .C0(n16160), .Y(
        n35559) );
  OA22XL U30827 ( .A0(net262304), .A1(n33578), .B0(n33586), .B1(n40128), .Y(
        n16711) );
  OAI211XL U30828 ( .A0(n33546), .A1(n42745), .B0(n16567), .C0(n16568), .Y(
        n35695) );
  OA22XL U30829 ( .A0(net218564), .A1(n33050), .B0(n33058), .B1(net218640),
        .Y(n15127) );
  OA22XL U30830 ( .A0(net262247), .A1(n33378), .B0(n33386), .B1(n40130), .Y(
        n16111) );
  OA22XL U30831 ( .A0(net262019), .A1(n33858), .B0(n33866), .B1(n40041), .Y(
        n17551) );
  OAI211XL U30832 ( .A0(n33714), .A1(n42753), .B0(n17071), .C0(n17072), .Y(
        n35863) );
  OA22XL U30833 ( .A0(net263881), .A1(n33106), .B0(n33114), .B1(n40045), .Y(
        n15295) );
  OAI211XL U30834 ( .A0(n32586), .A1(n42914), .B0(n13687), .C0(n13688), .Y(
        n34735) );
  XNOR2X1 U30835 ( .A(n36846), .B(n34082), .Y(n46192) );
  OA22XL U30836 ( .A0(net262855), .A1(n34082), .B0(n34090), .B1(n40103), .Y(
        n18223) );
  OA22XL U30837 ( .A0(net262855), .A1(n34074), .B0(n34082), .B1(n40103), .Y(
        n18199) );
  OAI211XL U30838 ( .A0(n32722), .A1(n42895), .B0(n14095), .C0(n14096), .Y(
        n34871) );
  OAI211XL U30839 ( .A0(n32706), .A1(n42865), .B0(n14047), .C0(n14048), .Y(
        n34855) );
  OAI211XL U30840 ( .A0(n32714), .A1(n42864), .B0(n14071), .C0(n14072), .Y(
        n34863) );
  OAI211XL U30841 ( .A0(n32570), .A1(n42916), .B0(n13639), .C0(n13640), .Y(
        n34719) );
  OA22XL U30842 ( .A0(net263045), .A1(n32626), .B0(n32634), .B1(n40093), .Y(
        n13855) );
  OA22XL U30843 ( .A0(net263045), .A1(n32618), .B0(n32626), .B1(n40093), .Y(
        n13831) );
  OAI211XL U30844 ( .A0(n32578), .A1(n42915), .B0(n13663), .C0(n13664), .Y(
        n34727) );
  OA22XL U30845 ( .A0(net263824), .A1(n32906), .B0(n32914), .B1(n40049), .Y(
        n14695) );
  OA22XL U30846 ( .A0(net263083), .A1(n32842), .B0(n32850), .B1(n40091), .Y(
        n14503) );
  OA22XL U30847 ( .A0(net263083), .A1(n32834), .B0(n32842), .B1(n40090), .Y(
        n14479) );
  OAI211XL U30848 ( .A0(n32538), .A1(n42921), .B0(n13543), .C0(n13544), .Y(
        n34687) );
  OA22XL U30849 ( .A0(net263102), .A1(n32826), .B0(n32834), .B1(n40090), .Y(
        n14455) );
  OAI211XL U30850 ( .A0(n32866), .A1(n42971), .B0(n14527), .C0(n14528), .Y(
        n35015) );
  OAI211XL U30851 ( .A0(n32874), .A1(n42970), .B0(n14551), .C0(n14552), .Y(
        n35023) );
  OAI211XL U30852 ( .A0(n32522), .A1(n42923), .B0(n13495), .C0(n13496), .Y(
        n34671) );
  OAI211XL U30853 ( .A0(n32530), .A1(n42922), .B0(n13519), .C0(n13520), .Y(
        n34679) );
  OAI211XL U30854 ( .A0(n32858), .A1(n42972), .B0(n14503), .C0(n14504), .Y(
        n35007) );
  OA22XL U30855 ( .A0(net262969), .A1(n32698), .B0(n32706), .B1(n40098), .Y(
        n14071) );
  OA22XL U30856 ( .A0(net262969), .A1(n32690), .B0(n32698), .B1(n40097), .Y(
        n14047) );
  OAI211XL U30857 ( .A0(n32650), .A1(n42873), .B0(n13879), .C0(n13880), .Y(
        n34799) );
  OA22XL U30858 ( .A0(net263672), .A1(n33314), .B0(n33322), .B1(n40126), .Y(
        n15919) );
  OA22XL U30859 ( .A0(net261905), .A1(n33706), .B0(n33714), .B1(n40149), .Y(
        n17095) );
  OA22XL U30860 ( .A0(net261905), .A1(n33698), .B0(n33706), .B1(n40148), .Y(
        n17071) );
  OA22XL U30861 ( .A0(net262722), .A1(n33946), .B0(n33954), .B1(n40084), .Y(
        n17815) );
  OA22XL U30862 ( .A0(net262741), .A1(n33938), .B0(n33946), .B1(n40108), .Y(
        n17791) );
  OA22XL U30863 ( .A0(net262019), .A1(n33850), .B0(n33858), .B1(net218850),
        .Y(n17527) );
  OA22XL U30864 ( .A0(net262019), .A1(n33842), .B0(n33850), .B1(n40142), .Y(
        n17503) );
  OAI211XL U30865 ( .A0(n33994), .A1(n42810), .B0(n17911), .C0(n17912), .Y(
        n36143) );
  OAI211XL U30866 ( .A0(n32986), .A1(n42986), .B0(n14887), .C0(n14888), .Y(
        n35135) );
  OA22XL U30867 ( .A0(net263881), .A1(n33114), .B0(n33122), .B1(n40046), .Y(
        n15319) );
  OAI211XL U30868 ( .A0(n33746), .A1(n42845), .B0(n17167), .C0(n17168), .Y(
        n35895) );
  OAI211XL U30869 ( .A0(n33954), .A1(n42847), .B0(n17791), .C0(n17792), .Y(
        n36103) );
  OAI211XL U30870 ( .A0(n33986), .A1(n42811), .B0(n17887), .C0(n17888), .Y(
        n36135) );
  OA22XL U30871 ( .A0(net262304), .A1(n33586), .B0(n33594), .B1(n40128), .Y(
        n16735) );
  OAI211XL U30872 ( .A0(n32634), .A1(n42875), .B0(n13831), .C0(n13832), .Y(
        n34783) );
  OA22XL U30873 ( .A0(net263634), .A1(n33338), .B0(n33346), .B1(n40059), .Y(
        n15991) );
  OAI211XL U30874 ( .A0(n32865), .A1(n42971), .B0(n14524), .C0(n14525), .Y(
        n35014) );
  OAI211XL U30875 ( .A0(n32404), .A1(n42908), .B0(n13141), .C0(n13142), .Y(
        n34553) );
  OA22XL U30876 ( .A0(net262703), .A1(n33970), .B0(n33978), .B1(n40109), .Y(
        n17887) );
  OAI211XL U30877 ( .A0(n33066), .A1(n42942), .B0(n15127), .C0(n15128), .Y(
        n35215) );
  OAI211XL U30878 ( .A0(n33274), .A1(n42945), .B0(n15751), .C0(n15752), .Y(
        n35423) );
  OA22XL U30879 ( .A0(net263900), .A1(n33098), .B0(n33106), .B1(n40045), .Y(
        n15271) );
  OA22XL U30880 ( .A0(net263900), .A1(n33090), .B0(n33098), .B1(n40044), .Y(
        n15247) );
  OA22XL U30881 ( .A0(net263634), .A1(n33346), .B0(n33354), .B1(n40059), .Y(
        n16015) );
  OA22XL U30882 ( .A0(net262000), .A1(n33866), .B0(n33874), .B1(n40143), .Y(
        n17575) );
  OAI211XL U30883 ( .A0(n33698), .A1(n42755), .B0(n17023), .C0(n17024), .Y(
        n35847) );
  OAI211XL U30884 ( .A0(n33418), .A1(n42795), .B0(n16183), .C0(n16184), .Y(
        n35567) );
  OA22XL U30885 ( .A0(net262190), .A1(n33426), .B0(n33434), .B1(n40133), .Y(
        n16255) );
  OA22XL U30886 ( .A0(net262209), .A1(n33418), .B0(n33426), .B1(n40133), .Y(
        n16231) );
  OA22XL U30887 ( .A0(net262361), .A1(n33530), .B0(n33538), .B1(n40125), .Y(
        n16567) );
  OA22XL U30888 ( .A0(net263957), .A1(n33042), .B0(n33050), .B1(n40042), .Y(
        n15103) );
  OAI211XL U30889 ( .A0(n33050), .A1(n42977), .B0(n15079), .C0(n15080), .Y(
        n35199) );
  OAI211XL U30890 ( .A0(n33002), .A1(n42984), .B0(n14935), .C0(n14936), .Y(
        n35151) );
  OAI211XL U30891 ( .A0(n33338), .A1(n42775), .B0(n15943), .C0(n15944), .Y(
        n35487) );
  OAI211XL U30892 ( .A0(n33378), .A1(n42769), .B0(n16063), .C0(n16064), .Y(
        n35527) );
  XOR2X1 U30893 ( .A(n33932), .B(n36829), .Y(n43582) );
  OAI211XL U30894 ( .A0(n33730), .A1(n42750), .B0(n17119), .C0(n17120), .Y(
        n35879) );
  OAI211XL U30895 ( .A0(n33738), .A1(n42846), .B0(n17143), .C0(n17144), .Y(
        n35887) );
  OAI211XL U30896 ( .A0(n33450), .A1(n42791), .B0(n16279), .C0(n16280), .Y(
        n35599) );
  OAI211XL U30897 ( .A0(n33642), .A1(n42763), .B0(n16855), .C0(n16856), .Y(
        n35791) );
  OA22XL U30898 ( .A0(net261924), .A1(n33682), .B0(n33690), .B1(n40147), .Y(
        n17023) );
  OA22XL U30899 ( .A0(net262874), .A1(n34066), .B0(n34074), .B1(n40102), .Y(
        n18175) );
  OA22XL U30900 ( .A0(net262285), .A1(n33594), .B0(n33602), .B1(n40078), .Y(
        n16759) );
  OA22XL U30901 ( .A0(net262285), .A1(n33602), .B0(n33610), .B1(net218866),
        .Y(n16783) );
  OA22XL U30902 ( .A0(net262380), .A1(n33506), .B0(n33514), .B1(n40123), .Y(
        n16495) );
  OA22XL U30903 ( .A0(net262114), .A1(n33498), .B0(n33506), .B1(n40138), .Y(
        n16471) );
  OAI211XL U30904 ( .A0(n33498), .A1(n42784), .B0(n16423), .C0(n16424), .Y(
        n35647) );
  OAI211XL U30905 ( .A0(n32786), .A1(n42885), .B0(n14287), .C0(n14288), .Y(
        n34935) );
  OAI211XL U30906 ( .A0(n32794), .A1(n42884), .B0(n14311), .C0(n14312), .Y(
        n34943) );
  OAI211XL U30907 ( .A0(n32778), .A1(n42886), .B0(n14263), .C0(n14264), .Y(
        n34927) );
  OAI211XL U30908 ( .A0(n32642), .A1(n42874), .B0(n13855), .C0(n13856), .Y(
        n34791) );
  OAI211XL U30909 ( .A0(n32658), .A1(n42872), .B0(n13903), .C0(n13904), .Y(
        n34807) );
  OA22XL U30910 ( .A0(net262133), .A1(n33490), .B0(n33498), .B1(n40137), .Y(
        n16447) );
  OA22XL U30911 ( .A0(net262133), .A1(n33482), .B0(n33490), .B1(n40137), .Y(
        n16423) );
  OAI211XL U30912 ( .A0(n33114), .A1(n42935), .B0(n15271), .C0(n15272), .Y(
        n35263) );
  OAI211XL U30913 ( .A0(n33122), .A1(n42934), .B0(n15295), .C0(n15296), .Y(
        n35271) );
  OA22XL U30914 ( .A0(net263539), .A1(n33186), .B0(n33194), .B1(n40065), .Y(
        n15535) );
  OA22XL U30915 ( .A0(net263539), .A1(n33178), .B0(n33186), .B1(n40065), .Y(
        n15511) );
  OA22XL U30916 ( .A0(net263007), .A1(n33234), .B0(n33242), .B1(n40068), .Y(
        n15679) );
  OAI211XL U30917 ( .A0(n32716), .A1(n42863), .B0(n14077), .C0(n14078), .Y(
        n34865) );
  OAI211XL U30918 ( .A0(n32708), .A1(n42864), .B0(n14053), .C0(n14054), .Y(
        n34857) );
  OAI211XL U30919 ( .A0(n32460), .A1(n42900), .B0(n13309), .C0(n13310), .Y(
        n34609) );
  OAI211XL U30920 ( .A0(n32561), .A1(n42918), .B0(n13612), .C0(n13613), .Y(
        n34710) );
  OAI211XL U30921 ( .A0(n32524), .A1(n42923), .B0(n13501), .C0(n13502), .Y(
        n34673) );
  OAI211XL U30922 ( .A0(n34026), .A1(n42805), .B0(n18007), .C0(n18008), .Y(
        n36175) );
  OA22XL U30923 ( .A0(net262722), .A1(n33954), .B0(n33962), .B1(n40091), .Y(
        n17839) );
  OA22XL U30924 ( .A0(net263710), .A1(n33266), .B0(n33274), .B1(n40055), .Y(
        n15775) );
  OAI211XL U30925 ( .A0(n33866), .A1(n42860), .B0(n17527), .C0(n17528), .Y(
        n36015) );
  OAI211XL U30926 ( .A0(n33594), .A1(n42738), .B0(n16711), .C0(n16712), .Y(
        n35743) );
  OAI211XL U30927 ( .A0(n33858), .A1(n42861), .B0(n17503), .C0(n17504), .Y(
        n36007) );
  OAI211XL U30928 ( .A0(n33610), .A1(n42737), .B0(n16759), .C0(n16760), .Y(
        n35759) );
  OAI211XL U30929 ( .A0(n33602), .A1(n42864), .B0(n16735), .C0(n16736), .Y(
        n35751) );
  OAI211XL U30930 ( .A0(n32994), .A1(n42985), .B0(n14911), .C0(n14912), .Y(
        n35143) );
  OAI211XL U30931 ( .A0(n33058), .A1(n42943), .B0(n15103), .C0(n15104), .Y(
        n35207) );
  OAI211XL U30932 ( .A0(n33106), .A1(n42937), .B0(n15247), .C0(n15248), .Y(
        n35255) );
  OAI211XL U30933 ( .A0(n33306), .A1(n42779), .B0(n15847), .C0(n15848), .Y(
        n35455) );
  OAI211XL U30934 ( .A0(n33138), .A1(n42932), .B0(n15343), .C0(n15344), .Y(
        n35287) );
  OAI211XL U30935 ( .A0(n33146), .A1(n42931), .B0(n15367), .C0(n15368), .Y(
        n35295) );
  OAI211XL U30936 ( .A0(n33178), .A1(n42958), .B0(n15463), .C0(n15464), .Y(
        n35327) );
  OA22XL U30937 ( .A0(net263691), .A1(n33282), .B0(n33290), .B1(n40056), .Y(
        n15823) );
  OA22XL U30938 ( .A0(net263710), .A1(n33274), .B0(n33282), .B1(n40056), .Y(
        n15799) );
  OAI211XL U30939 ( .A0(n33194), .A1(n42956), .B0(n15511), .C0(n15512), .Y(
        n35343) );
  OAI211XL U30940 ( .A0(n33226), .A1(n42951), .B0(n15607), .C0(n15608), .Y(
        n35375) );
  OAI211XL U30941 ( .A0(n33234), .A1(n42950), .B0(n15631), .C0(n15632), .Y(
        n35383) );
  OAI211XL U30942 ( .A0(n33186), .A1(n42957), .B0(n15487), .C0(n15488), .Y(
        n35335) );
  OAI211XL U30943 ( .A0(n33010), .A1(n42982), .B0(n14959), .C0(n14960), .Y(
        n35159) );
  OA22XL U30944 ( .A0(net262912), .A1(n34034), .B0(n34042), .B1(n40101), .Y(
        n18079) );
  OA22XL U30945 ( .A0(net262912), .A1(n34026), .B0(n34034), .B1(n40101), .Y(
        n18055) );
  XNOR2X1 U30946 ( .A(n50524), .B(n36709), .Y(n25205) );
  OAI211XL U30947 ( .A0(n32585), .A1(n42914), .B0(n13684), .C0(n13685), .Y(
        n34734) );
  OAI211XL U30948 ( .A0(n32428), .A1(n42905), .B0(n13213), .C0(n13214), .Y(
        n34577) );
  OAI211XL U30949 ( .A0(n32569), .A1(n42916), .B0(n13636), .C0(n13637), .Y(
        n34718) );
  OAI211XL U30950 ( .A0(n32601), .A1(n42912), .B0(n13732), .C0(n13733), .Y(
        n34750) );
  OAI211XL U30951 ( .A0(n32609), .A1(n42879), .B0(n13756), .C0(n13757), .Y(
        n34758) );
  OAI211XL U30952 ( .A0(n32593), .A1(n42913), .B0(n13708), .C0(n13709), .Y(
        n34742) );
  OAI211XL U30953 ( .A0(n32553), .A1(n42919), .B0(n13588), .C0(n13589), .Y(
        n34702) );
  OAI211XL U30954 ( .A0(n32489), .A1(n42896), .B0(n13396), .C0(n13397), .Y(
        n34638) );
  OAI211XL U30955 ( .A0(n32801), .A1(n42883), .B0(n14332), .C0(n14333), .Y(
        n34950) );
  OAI211XL U30956 ( .A0(n32617), .A1(n42878), .B0(n13780), .C0(n13781), .Y(
        n34766) );
  XNOR2X1 U30957 ( .A(n33778), .B(n42565), .Y(n46175) );
  XOR2X1 U30958 ( .A(n34427), .B(n36881), .Y(n45035) );
  XOR2X1 U30959 ( .A(n34420), .B(n42637), .Y(n45039) );
  XOR2X1 U30960 ( .A(n34420), .B(n36822), .Y(n45282) );
  XOR2X1 U30961 ( .A(n34431), .B(n42515), .Y(n45228) );
  XOR2X1 U30962 ( .A(n34431), .B(n42612), .Y(n45261) );
  OAI211XL U30963 ( .A0(n34097), .A1(n42827), .B0(n18220), .C0(n18221), .Y(
        n36246) );
  OAI211XL U30964 ( .A0(n34098), .A1(n42827), .B0(n18223), .C0(n18224), .Y(
        n36247) );
  OAI211XL U30965 ( .A0(n32972), .A1(n42988), .B0(n14845), .C0(n14846), .Y(
        n35121) );
  OAI211XL U30966 ( .A0(n32964), .A1(n42989), .B0(n14821), .C0(n14822), .Y(
        n35113) );
  OAI211XL U30967 ( .A0(n32548), .A1(n42920), .B0(n13573), .C0(n13574), .Y(
        n34697) );
  OAI211XL U30968 ( .A0(n32540), .A1(n42921), .B0(n13549), .C0(n13550), .Y(
        n34689) );
  XOR2X1 U30969 ( .A(n34422), .B(n42533), .Y(n45279) );
  OAI211XL U30970 ( .A0(n32740), .A1(n42892), .B0(n14149), .C0(n14150), .Y(
        n34889) );
  OAI211XL U30971 ( .A0(n32572), .A1(n42916), .B0(n13645), .C0(n13646), .Y(
        n34721) );
  OAI211XL U30972 ( .A0(n32580), .A1(n42915), .B0(n13669), .C0(n13670), .Y(
        n34729) );
  OAI211XL U30973 ( .A0(n32564), .A1(n42917), .B0(n13621), .C0(n13622), .Y(
        n34713) );
  OAI211XL U30974 ( .A0(n32468), .A1(n42899), .B0(n13333), .C0(n13334), .Y(
        n34617) );
  OAI211XL U30975 ( .A0(n32476), .A1(n42898), .B0(n13357), .C0(n13358), .Y(
        n34625) );
  OAI211XL U30976 ( .A0(n32484), .A1(n42896), .B0(n13381), .C0(n13382), .Y(
        n34633) );
  OAI211XL U30977 ( .A0(n32956), .A1(n42990), .B0(n14797), .C0(n14798), .Y(
        n35105) );
  OAI211XL U30978 ( .A0(n32492), .A1(n42895), .B0(n13405), .C0(n13406), .Y(
        n34641) );
  OAI211XL U30979 ( .A0(n32860), .A1(n42972), .B0(n14509), .C0(n14510), .Y(
        n35009) );
  OAI211XL U30980 ( .A0(n32868), .A1(n42971), .B0(n14533), .C0(n14534), .Y(
        n35017) );
  OAI211XL U30981 ( .A0(n32876), .A1(n42970), .B0(n14557), .C0(n14558), .Y(
        n35025) );
  OAI211XL U30982 ( .A0(n32532), .A1(n42922), .B0(n13525), .C0(n13526), .Y(
        n34681) );
  OAI211XL U30983 ( .A0(n32417), .A1(n42906), .B0(n13180), .C0(n13181), .Y(
        n34566) );
  OAI211XL U30984 ( .A0(n32732), .A1(n42893), .B0(n14125), .C0(n14126), .Y(
        n34881) );
  OAI211XL U30985 ( .A0(n32596), .A1(n42913), .B0(n13717), .C0(n13718), .Y(
        n34745) );
  OAI211XL U30986 ( .A0(n32604), .A1(n42911), .B0(n13741), .C0(n13742), .Y(
        n34753) );
  OAI211XL U30987 ( .A0(n32425), .A1(n42905), .B0(n13204), .C0(n13205), .Y(
        n34574) );
  XOR2X1 U30988 ( .A(n36853), .B(n34424), .Y(n46598) );
  XOR2X1 U30989 ( .A(n34424), .B(net219434), .Y(n45010) );
  XOR2X1 U30990 ( .A(n34424), .B(n36730), .Y(n45277) );
  OAI211XL U30991 ( .A0(n32724), .A1(n42894), .B0(n14101), .C0(n14102), .Y(
        n34873) );
  OAI211XL U30992 ( .A0(n32713), .A1(n42864), .B0(n14068), .C0(n14069), .Y(
        n34862) );
  OAI211XL U30993 ( .A0(n32588), .A1(n42914), .B0(n13693), .C0(n13694), .Y(
        n34737) );
  OAI211XL U30994 ( .A0(n32780), .A1(n42886), .B0(n14269), .C0(n14270), .Y(
        n34929) );
  OAI211XL U30995 ( .A0(n32788), .A1(n42885), .B0(n14293), .C0(n14294), .Y(
        n34937) );
  OAI211XL U30996 ( .A0(n32796), .A1(n42884), .B0(n14317), .C0(n14318), .Y(
        n34945) );
  OAI211XL U30997 ( .A0(n32804), .A1(n42883), .B0(n14341), .C0(n14342), .Y(
        n34953) );
  OAI211XL U30998 ( .A0(n32620), .A1(n42877), .B0(n13789), .C0(n13790), .Y(
        n34769) );
  XOR2X1 U30999 ( .A(n34421), .B(n42549), .Y(n45280) );
  XOR2X1 U31000 ( .A(n34421), .B(n41281), .Y(n45007) );
  NAND2X1 U31001 ( .A(n34421), .B(n36802), .Y(n41644) );
  XOR2X1 U31002 ( .A(n34198), .B(net219330), .Y(n44112) );
  XOR2X1 U31003 ( .A(n34197), .B(n41281), .Y(n44113) );
  XNOR2X1 U31004 ( .A(n34336), .B(n36730), .Y(n45226) );
  XNOR2X1 U31005 ( .A(n36856), .B(n34336), .Y(n46520) );
  XNOR2X1 U31006 ( .A(n36856), .B(n34152), .Y(n46230) );
  XOR2X1 U31007 ( .A(n34204), .B(n42697), .Y(n44145) );
  XNOR2X1 U31008 ( .A(n36851), .B(n34216), .Y(n46399) );
  XNOR2XL U31009 ( .A(n34216), .B(n42504), .Y(n44671) );
  XOR2X1 U31010 ( .A(n34150), .B(n42617), .Y(n43981) );
  XNOR2X1 U31011 ( .A(n36856), .B(n34344), .Y(n46542) );
  XOR2X1 U31012 ( .A(n34289), .B(n42719), .Y(n45362) );
  XOR2X1 U31013 ( .A(n34297), .B(n34435), .Y(n45393) );
  XOR2X1 U31014 ( .A(n34258), .B(n41641), .Y(n44809) );
  XOR2X1 U31015 ( .A(n34257), .B(n34435), .Y(n44810) );
  XOR2X1 U31016 ( .A(n34298), .B(n41642), .Y(n45392) );
  XOR2X1 U31017 ( .A(n36766), .B(n34361), .Y(n47606) );
  XOR2X1 U31018 ( .A(n34318), .B(net219336), .Y(n45476) );
  XOR2X1 U31019 ( .A(n34341), .B(n34447), .Y(n45200) );
  XNOR2X1 U31020 ( .A(n36853), .B(n34280), .Y(n46374) );
  XOR2X1 U31021 ( .A(n34214), .B(n42538), .Y(n44663) );
  XOR2X1 U31022 ( .A(n34337), .B(n42680), .Y(n45204) );
  XNOR2X1 U31023 ( .A(n34360), .B(n42501), .Y(n44993) );
  XNOR2X1 U31024 ( .A(n36851), .B(n34360), .Y(n46498) );
  XOR2X1 U31025 ( .A(n34349), .B(n42630), .Y(n45111) );
  XNOR2X1 U31026 ( .A(n34382), .B(n42538), .Y(n44905) );
  XNOR2X1 U31027 ( .A(n34381), .B(n42550), .Y(n44904) );
  XNOR2X1 U31028 ( .A(n34312), .B(n34458), .Y(n45464) );
  XNOR2X1 U31029 ( .A(n34288), .B(n42505), .Y(n45407) );
  XNOR2X1 U31030 ( .A(n34296), .B(n42505), .Y(net213701) );
  XOR2X1 U31031 ( .A(n34202), .B(n42705), .Y(n44147) );
  OAI211XL U31032 ( .A0(n32889), .A1(n42968), .B0(n14596), .C0(n14597), .Y(
        n35038) );
  OAI211XL U31033 ( .A0(n32897), .A1(n42966), .B0(n14620), .C0(n14621), .Y(
        n35046) );
  OAI211XL U31034 ( .A0(n32881), .A1(n42969), .B0(n14572), .C0(n14573), .Y(
        n35030) );
  XOR2X1 U31035 ( .A(n34290), .B(n42705), .Y(n45361) );
  XOR2X1 U31036 ( .A(n34366), .B(n36868), .Y(n44967) );
  XOR2X1 U31037 ( .A(n34365), .B(n36832), .Y(n44942) );
  XOR2X1 U31038 ( .A(n34320), .B(net219468), .Y(n45474) );
  XNOR2X1 U31039 ( .A(n34304), .B(n42505), .Y(net213732) );
  XNOR2X1 U31040 ( .A(n34389), .B(n42552), .Y(n45102) );
  XOR2X1 U31041 ( .A(n34389), .B(n41281), .Y(n44921) );
  XOR2X1 U31042 ( .A(n34144), .B(net219444), .Y(n43894) );
  XOR2X1 U31043 ( .A(n34306), .B(n42558), .Y(n45461) );
  OAI211XL U31044 ( .A0(n32753), .A1(n42890), .B0(n14188), .C0(n14189), .Y(
        n34902) );
  OAI211XL U31045 ( .A0(n32761), .A1(n42889), .B0(n14212), .C0(n14213), .Y(
        n34910) );
  OAI211XL U31046 ( .A0(n32505), .A1(n42926), .B0(n13444), .C0(n13445), .Y(
        n34654) );
  OAI211XL U31047 ( .A0(n32641), .A1(n42874), .B0(n13852), .C0(n13853), .Y(
        n34790) );
  XOR2X1 U31048 ( .A(n34390), .B(n36868), .Y(n44882) );
  XOR2X1 U31049 ( .A(n36860), .B(n34400), .Y(n46588) );
  XOR2X1 U31050 ( .A(n34406), .B(net219308), .Y(n45092) );
  XOR2X1 U31051 ( .A(n34406), .B(n42613), .Y(n45065) );
  XOR2X1 U31052 ( .A(n34384), .B(n42592), .Y(n44910) );
  XOR2X1 U31053 ( .A(n34378), .B(n42672), .Y(n44916) );
  OAI211XL U31054 ( .A0(n32625), .A1(n42876), .B0(n13804), .C0(n13805), .Y(
        n34774) );
  OAI211XL U31055 ( .A0(n32433), .A1(n42904), .B0(n13228), .C0(n13229), .Y(
        n34582) );
  OAI211XL U31056 ( .A0(n32441), .A1(n42903), .B0(n13252), .C0(n13253), .Y(
        n34590) );
  OAI211XL U31057 ( .A0(n32449), .A1(n42901), .B0(n13276), .C0(n13277), .Y(
        n34598) );
  OAI211XL U31058 ( .A0(n32769), .A1(n42888), .B0(n14236), .C0(n14237), .Y(
        n34918) );
  OAI211XL U31059 ( .A0(n32633), .A1(n42875), .B0(n13828), .C0(n13829), .Y(
        n34782) );
  OAI211XL U31060 ( .A0(n32497), .A1(n42927), .B0(n13420), .C0(n13421), .Y(
        n34646) );
  OAI211XL U31061 ( .A0(n32513), .A1(n42925), .B0(n13468), .C0(n13469), .Y(
        n34662) );
  XOR2X1 U31062 ( .A(n34168), .B(net219450), .Y(n43956) );
  XNOR2X1 U31063 ( .A(n51119), .B(n42552), .Y(n31831) );
  NOR2XL U31064 ( .A(n50147), .B(n50148), .Y(n9704) );
  XNOR2XL U31065 ( .A(n32399), .B(n50147), .Y(n9726) );
  NAND2X1 U31066 ( .A(n34423), .B(n36908), .Y(n41206) );
  XOR2X1 U31067 ( .A(n34376), .B(net219434), .Y(n44973) );
  XNOR2X1 U31068 ( .A(n34376), .B(n42505), .Y(n44937) );
  XOR2X1 U31069 ( .A(n34200), .B(net219468), .Y(n44110) );
  XOR2X1 U31070 ( .A(n34419), .B(n42659), .Y(n45033) );
  XOR2X1 U31071 ( .A(n34419), .B(n36877), .Y(n45281) );
  XOR2X1 U31072 ( .A(n34393), .B(n36875), .Y(n44895) );
  XOR2X1 U31073 ( .A(n34393), .B(n42575), .Y(n45059) );
  XOR2X1 U31074 ( .A(n34248), .B(n42592), .Y(n44764) );
  XOR2X1 U31075 ( .A(n34394), .B(n42705), .Y(n44894) );
  XOR2X1 U31076 ( .A(n34394), .B(n42557), .Y(n45061) );
  XOR2X1 U31077 ( .A(n36847), .B(n34394), .Y(n46593) );
  XOR2X1 U31078 ( .A(n34397), .B(n42629), .Y(n45085) );
  XOR2X1 U31079 ( .A(n34397), .B(n36832), .Y(n45057) );
  XOR2X1 U31080 ( .A(n34358), .B(n36868), .Y(n45139) );
  XOR2X1 U31081 ( .A(n34358), .B(n42533), .Y(n44985) );
  XOR2X1 U31082 ( .A(n34350), .B(net219310), .Y(n45207) );
  XOR2X1 U31083 ( .A(n41293), .B(n34350), .Y(n46545) );
  XOR2X1 U31084 ( .A(n34324), .B(n42638), .Y(n45421) );
  XOR2X1 U31085 ( .A(n34324), .B(n36825), .Y(n45191) );
  XOR2X1 U31086 ( .A(n41302), .B(n34324), .Y(n46527) );
  XOR2X1 U31087 ( .A(n34328), .B(net219468), .Y(n45445) );
  XNOR2X1 U31088 ( .A(n34328), .B(n42505), .Y(n45195) );
  XNOR2X1 U31089 ( .A(n36852), .B(n34328), .Y(n46531) );
  NAND2X1 U31090 ( .A(n34201), .B(n41228), .Y(n41229) );
  NAND2X1 U31091 ( .A(n34368), .B(n42509), .Y(n41350) );
  XOR2X1 U31092 ( .A(n34386), .B(n42705), .Y(n44924) );
  XNOR2X1 U31093 ( .A(n34386), .B(n42560), .Y(n45098) );
  XNOR2X1 U31094 ( .A(n36845), .B(n34386), .Y(n46579) );
  XNOR2X1 U31095 ( .A(n36733), .B(n34386), .Y(n47687) );
  NAND2X1 U31096 ( .A(n34408), .B(net259034), .Y(n41235) );
  XOR2X1 U31097 ( .A(n34398), .B(n36870), .Y(n44890) );
  XOR2X1 U31098 ( .A(n34398), .B(n42538), .Y(n45058) );
  NAND2X1 U31099 ( .A(n34208), .B(n37015), .Y(n41232) );
  XOR2X1 U31100 ( .A(n34364), .B(n42637), .Y(n44969) );
  NAND2X1 U31101 ( .A(n34364), .B(n36923), .Y(n41271) );
  INVX12 U31102 ( .A(n37536), .Y(codeword[5]) );
  INVX12 U31103 ( .A(n37538), .Y(enc_num[11]) );
  INVX12 U31104 ( .A(n37537), .Y(enc_num[10]) );
  INVX12 U31105 ( .A(n37539), .Y(enc_num[9]) );
  INVX12 U31106 ( .A(n37531), .Y(enc_num[8]) );
  INVX12 U31107 ( .A(n37532), .Y(enc_num[7]) );
  INVX12 U31108 ( .A(n37533), .Y(enc_num[6]) );
  INVX12 U31109 ( .A(n37524), .Y(enc_num[1]) );
  INVX12 U31110 ( .A(n37523), .Y(enc_num[2]) );
  INVX12 U31111 ( .A(n37522), .Y(enc_num[3]) );
  INVX12 U31112 ( .A(n37535), .Y(enc_num[4]) );
  INVX12 U31113 ( .A(n37534), .Y(enc_num[5]) );
  INVX12 U31114 ( .A(n37521), .Y(enc_num[0]) );
  CLKINVX1 U31115 ( .A(n37600), .Y(n37589) );
  INVX12 U31116 ( .A(n37589), .Y(n37590) );
  INVX12 U31117 ( .A(n37589), .Y(n37591) );
  INVX20 U31118 ( .A(n37597), .Y(n37592) );
  INVX20 U31119 ( .A(n37597), .Y(n37593) );
  INVX16 U31120 ( .A(reset), .Y(n37594) );
  INVX16 U31121 ( .A(reset), .Y(n37595) );
  INVX16 U31122 ( .A(reset), .Y(n37596) );
  INVX20 U31123 ( .A(n37597), .Y(n37599) );
  INVX20 U31124 ( .A(n37597), .Y(n37600) );
  INVX20 U31125 ( .A(n37597), .Y(n37601) );
  NAND2BX4 U32515 ( .AN(n39293), .B(net214879), .Y(n10543) );
  NAND2BX4 U32516 ( .AN(n39307), .B(net214389), .Y(net209930) );
  NAND3X6 U32517 ( .A(n39308), .B(net213703), .C(net213700), .Y(net209894) );
  NAND2BX4 U32518 ( .AN(n39318), .B(net216020), .Y(n10559) );
  NAND2BX4 U32519 ( .AN(n39323), .B(net215271), .Y(n10608) );
  NAND2BX4 U32520 ( .AN(n39324), .B(net215298), .Y(n10607) );
  NAND2BX4 U32521 ( .AN(n39325), .B(net215289), .Y(n10606) );
  NAND2BX4 U32522 ( .AN(n_cell_301249_net267075), .B(net211962), .Y(n39345) );
  NAND2BX4 U32523 ( .AN(n39371), .B(net211147), .Y(n10044) );
  NAND2BX4 U32524 ( .AN(n39372), .B(net211152), .Y(n10045) );
  NAND2BX4 U32525 ( .AN(n39404), .B(net213402), .Y(n10852) );
  NAND2BX4 U32526 ( .AN(n39405), .B(net212711), .Y(n10855) );
  NAND2BX4 U32527 ( .AN(n39406), .B(net212716), .Y(n10854) );
  NAND2BX4 U32528 ( .AN(n39407), .B(net212726), .Y(n10853) );
  NAND2BX4 U32529 ( .AN(n39410), .B(net213357), .Y(n10863) );
  NAND2BX4 U32530 ( .AN(n39411), .B(net213352), .Y(n10872) );
  CLKINVX6 U32531 ( .A(net209253), .Y(net171433) );
  NAND2BX4 U32532 ( .AN(n39413), .B(net212691), .Y(n11147) );
  NAND4BX4 U32533 ( .AN(n37236), .B(net215432), .C(net215429), .D(net215430),
        .Y(n10395) );
  NAND4BX4 U32534 ( .AN(n37220), .B(net215821), .C(net215818), .D(net215819),
        .Y(net209565) );
  NAND3X6 U32535 ( .A(net215438), .B(net215439), .C(n39458), .Y(n10126) );
  NAND3X6 U32536 ( .A(net215827), .B(net215828), .C(n39459), .Y(n10128) );
  NAND4X4 U32537 ( .A(net215402), .B(net215403), .C(net215404), .D(net215405),
        .Y(n10387) );
  NAND4X4 U32538 ( .A(net215375), .B(net215376), .C(net215377), .D(net215378),
        .Y(n10385) );
  NAND3X6 U32539 ( .A(net215395), .B(net215396), .C(n39465), .Y(n10384) );
  NAND4BX4 U32540 ( .AN(n37218), .B(net215385), .C(net215386), .D(net215387),
        .Y(n10383) );
  NAND4BX4 U32541 ( .AN(n37302), .B(net215304), .C(net215305), .D(net215306),
        .Y(n10423) );
  OR4X8 U32542 ( .A(net171425), .B(net171427), .C(net151673), .D(net151712),
        .Y(n39505) );
  NOR2BX4 U32543 ( .AN(net214154), .B(n37234), .Y(n39463) );
  NAND2X4 U32544 ( .A(n39776), .B(net214392), .Y(n39307) );
  NAND2X4 U32545 ( .A(n39784), .B(net215274), .Y(n39323) );
  NAND3X6 U32546 ( .A(net213364), .B(net213365), .C(net213363), .Y(n39412) );
  NAND2X4 U32547 ( .A(n39951), .B(net213350), .Y(n39424) );
  NAND2X4 U32548 ( .A(n39955), .B(net213360), .Y(n39410) );
  NAND2X4 U32549 ( .A(n39960), .B(net212719), .Y(n39406) );
  NAND2X4 U32550 ( .A(n39961), .B(net212714), .Y(n39405) );
  INVX8 U32551 ( .A(n12024), .Y(net171214) );
  INVX8 U32552 ( .A(n40386), .Y(net171218) );
  INVX6 U32553 ( .A(n11398), .Y(net171551) );
  NOR2X8 U32554 ( .A(n37009), .B(n37231), .Y(n39459) );
  NOR2X8 U32555 ( .A(n37105), .B(n37314), .Y(n39784) );
  NOR2X8 U32556 ( .A(n36951), .B(n37335), .Y(n39955) );
  NOR2X8 U32557 ( .A(n36950), .B(n37334), .Y(n39951) );
  AND2X6 U32558 ( .A(net214391), .B(net214390), .Y(n39776) );
  NAND2BX4 U32559 ( .AN(n_cell_301249_net267379), .B(net216328), .Y(
        n_cell_303546_net275967) );
  AOI21X4 U32560 ( .A0(n40477), .A1(n40478), .B0(n40479), .Y(n40476) );
  AOI21X4 U32561 ( .A0(n11874), .A1(n40509), .B0(n_cell_303546_net277494), .Y(
        n40508) );
  NOR2X6 U32562 ( .A(n40508), .B(n_cell_303546_net277496), .Y(n40510) );
  AOI21X4 U32563 ( .A0(n40512), .A1(n11551), .B0(n_cell_303546_net277497), .Y(
        n40511) );
  AOI21X4 U32564 ( .A0(n40521), .A1(n40522), .B0(n40523), .Y(n40520) );
  AOI21X4 U32565 ( .A0(n40526), .A1(n40527), .B0(n40528), .Y(n40525) );
  NOR2X6 U32566 ( .A(n40525), .B(n40530), .Y(n40529) );
  AOI21X4 U32567 ( .A0(n40532), .A1(n40533), .B0(n40534), .Y(n40531) );
  AOI21X4 U32568 ( .A0(n40551), .A1(n40552), .B0(n40553), .Y(n40550) );
  AOI21X4 U32569 ( .A0(n40555), .A1(n40556), .B0(n40557), .Y(n40554) );
  AOI21X4 U32570 ( .A0(n40559), .A1(n40560), .B0(n40561), .Y(n40558) );
  AOI21X4 U32571 ( .A0(n40563), .A1(net210555), .B0(n40002), .Y(n40562) );
  AOI21X4 U32572 ( .A0(n_cell_303546_net277735), .A1(n10957), .B0(n40658), .Y(
        n40552) );
  OAI21X4 U32573 ( .A0(n10205), .A1(net151584), .B0(n40659), .Y(n40553) );
  AOI21X4 U32574 ( .A0(n_cell_303546_net277759), .A1(n10928), .B0(n40676), .Y(
        n40677) );
  OAI21X4 U32575 ( .A0(n40467), .A1(n40725), .B0(n40728), .Y(n40761) );
  OAI21X4 U32576 ( .A0(n40474), .A1(n40734), .B0(n40737), .Y(n40477) );
  OAI21X4 U32577 ( .A0(n40476), .A1(n40743), .B0(n40745), .Y(n40762) );
  OAI21X4 U32578 ( .A0(n40497), .A1(n40622), .B0(n40624), .Y(n40765) );
  NAND2X4 U32579 ( .A(n40765), .B(n40626), .Y(n40503) );
  OAI21X4 U32580 ( .A0(n_cell_303546_net277957), .A1(n40510), .B0(n10064), .Y(
        n40512) );
  OAI21X4 U32581 ( .A0(n39699), .A1(n40511), .B0(n11550), .Y(n40767) );
  OAI21X4 U32582 ( .A0(net259031), .A1(n40687), .B0(n40690), .Y(n40522) );
  OAI21X4 U32583 ( .A0(n40520), .A1(n40694), .B0(n40697), .Y(n40768) );
  NAND2X4 U32584 ( .A(n40768), .B(n40698), .Y(n40526) );
  OAI21X4 U32585 ( .A0(n40529), .A1(n40705), .B0(n40708), .Y(n40769) );
  NAND2X4 U32586 ( .A(n40709), .B(n40769), .Y(n40532) );
  OAI21X4 U32587 ( .A0(n40548), .A1(n40654), .B0(n40657), .Y(n40551) );
  OAI21X4 U32588 ( .A0(n40550), .A1(n40662), .B0(n40665), .Y(n40771) );
  NAND2X4 U32589 ( .A(n40667), .B(n40771), .Y(n40555) );
  OAI21X4 U32590 ( .A0(n40554), .A1(n40674), .B0(n40677), .Y(n40560) );
  OAI21X4 U32591 ( .A0(n40558), .A1(n40681), .B0(net210556), .Y(n40563) );
  NAND3X8 U32592 ( .A(n12194), .B(n10928), .C(n40675), .Y(n40674) );
  NAND3X6 U32593 ( .A(n40802), .B(n40803), .C(n40804), .Y(net152412) );
  NOR2X6 U32594 ( .A(n10994), .B(n37179), .Y(n40805) );
  NOR2X6 U32595 ( .A(n40805), .B(n40807), .Y(n40806) );
  AOI21X4 U32596 ( .A0(n40809), .A1(n40810), .B0(n40811), .Y(n40808) );
  AOI21X4 U32597 ( .A0(n40813), .A1(n40814), .B0(n40815), .Y(n40812) );
  AOI21X4 U32598 ( .A0(n40817), .A1(n40818), .B0(n40819), .Y(n40816) );
  AOI21X4 U32599 ( .A0(n40821), .A1(n40822), .B0(n40823), .Y(n40820) );
  AOI21X4 U32600 ( .A0(n40825), .A1(n40826), .B0(n40827), .Y(n40824) );
  AOI21X4 U32601 ( .A0(n40843), .A1(n40844), .B0(n40845), .Y(n40842) );
  NOR2X6 U32602 ( .A(n40842), .B(n40847), .Y(n40846) );
  AOI21X4 U32603 ( .A0(n40861), .A1(n40862), .B0(n40863), .Y(n40860) );
  AOI21X4 U32604 ( .A0(n40895), .A1(n40896), .B0(n40897), .Y(n40894) );
  AOI21X4 U32605 ( .A0(n40906), .A1(n40907), .B0(n40908), .Y(n40905) );
  NAND2X4 U32606 ( .A(n41147), .B(n41146), .Y(n41148) );
  NOR2X6 U32607 ( .A(net171414), .B(net171412), .Y(n41168) );
  OAI21X4 U32608 ( .A0(n37120), .A1(n_cell_301249_net269022), .B0(n41170), .Y(
        n41171) );
  AOI21X4 U32609 ( .A0(n41122), .A1(n41190), .B0(n40913), .Y(n40802) );
  OAI21X4 U32610 ( .A0(n40806), .A1(n41148), .B0(n41155), .Y(n40809) );
  OAI21X4 U32611 ( .A0(n40808), .A1(n41163), .B0(n41164), .Y(n40814) );
  OAI21X4 U32612 ( .A0(n40812), .A1(n41167), .B0(n41168), .Y(n40818) );
  OAI21X4 U32613 ( .A0(n40816), .A1(n41171), .B0(n41172), .Y(n40822) );
  OAI21X4 U32614 ( .A0(n40820), .A1(n41175), .B0(n41178), .Y(n40825) );
  OAI21X4 U32615 ( .A0(n40832), .A1(n41081), .B0(n41087), .Y(n40835) );
  OAI21X4 U32616 ( .A0(n40838), .A1(n41102), .B0(n41103), .Y(n40843) );
  OAI21X4 U32617 ( .A0(n40850), .A1(n41115), .B0(n41116), .Y(n40856) );
  OAI21X4 U32618 ( .A0(n40864), .A1(n41037), .B0(n41040), .Y(n40867) );
  OAI21X4 U32619 ( .A0(n40901), .A1(n41012), .B0(n41013), .Y(n40907) );
  OAI21X4 U32620 ( .A0(n40905), .A1(n41016), .B0(n41017), .Y(n40911) );
  NAND2X4 U32621 ( .A(n41187), .B(n41192), .Y(n40803) );
  CLKINVX12 U32622 ( .A(net260488), .Y(net151420) );
  NOR2X8 U32623 ( .A(n_cell_301249_net269831), .B(n39481), .Y(n41172) );
  NAND2X6 U32624 ( .A(n10958), .B(n10957), .Y(n41167) );
  NOR4X8 U32625 ( .A(n41153), .B(n41152), .C(net171401), .D(net171396), .Y(
        n41155) );
  NAND4XL U32626 ( .A(n37468), .B(net209308), .C(net209311), .D(n41764), .Y(
        n47798) );
  NOR2X4 U32627 ( .A(n47347), .B(net209308), .Y(n47357) );
  XOR2XL U32628 ( .A(n41319), .B(n34121), .Y(n43862) );
  NOR2BX1 U32629 ( .AN(net209900), .B(net209899), .Y(n47714) );
  NAND4X4 U32630 ( .A(n45454), .B(n45453), .C(n45452), .D(n45451), .Y(
        net209606) );
  NOR4X2 U32631 ( .A(n45440), .B(n45439), .C(n45438), .D(n45437), .Y(n45454)
         );
  NAND4X2 U32632 ( .A(n45747), .B(n45746), .C(n45745), .D(n45744), .Y(
        net211656) );
  NOR2X4 U32633 ( .A(n47391), .B(net209300), .Y(n47401) );
  XOR2X1 U32634 ( .A(n36765), .B(n34369), .Y(n47617) );
  NAND4X4 U32635 ( .A(n44177), .B(n44176), .C(n44175), .D(n44174), .Y(n12751)
         );
  XOR2X1 U32636 ( .A(n34366), .B(net219310), .Y(n45147) );
  XOR2X1 U32637 ( .A(n36733), .B(n34402), .Y(n47680) );
  NOR4X1 U32638 ( .A(n44947), .B(n44946), .C(n44945), .D(n44944), .Y(n44963)
         );
  XOR2X1 U32639 ( .A(n34402), .B(n42670), .Y(n45069) );
  NOR2X8 U32640 ( .A(n12746), .B(n45693), .Y(net213347) );
  INVX1 U32641 ( .A(net209320), .Y(net210772) );
  XOR2X1 U32642 ( .A(n34396), .B(n41385), .Y(n44892) );
  NOR2X2 U32643 ( .A(n47402), .B(net209298), .Y(n47412) );
  XOR2X1 U32644 ( .A(n41827), .B(n36895), .Y(n44682) );
  INVXL U32645 ( .A(n48435), .Y(n48445) );
  NOR4X1 U32646 ( .A(n45481), .B(n45480), .C(n45479), .D(n45478), .Y(n45482)
         );
  XOR2X1 U32647 ( .A(n34316), .B(n42693), .Y(n45478) );
  XNOR2XL U32648 ( .A(n36857), .B(n34240), .Y(n46454) );
  XOR2X1 U32649 ( .A(n34317), .B(n41282), .Y(n45477) );
  XOR2X1 U32650 ( .A(n42071), .B(n42660), .Y(n45142) );
  NOR2X2 U32651 ( .A(n47468), .B(net209296), .Y(n47478) );
  XOR2X1 U32652 ( .A(n34222), .B(net219314), .Y(n44743) );
  XOR2X1 U32653 ( .A(n42495), .B(n42081), .Y(n47350) );
  AOI21X1 U32654 ( .A0(n47987), .A1(net210209), .B0(net210210), .Y(n47988) );
  NOR2X4 U32655 ( .A(net210567), .B(net209289), .Y(n47785) );
  NOR4X4 U32656 ( .A(n45074), .B(n45073), .C(n45072), .D(n45071), .Y(n45078)
         );
  XOR2X1 U32657 ( .A(n34285), .B(n41283), .Y(n45300) );
  XOR2X1 U32658 ( .A(n42065), .B(n42659), .Y(n45068) );
  NOR2X2 U32659 ( .A(n47612), .B(n48441), .Y(n47622) );
  XOR2X1 U32660 ( .A(n34306), .B(n42707), .Y(n45506) );
  NOR4X2 U32661 ( .A(n45448), .B(n45447), .C(n45446), .D(n45445), .Y(n45452)
         );
  NOR4X2 U32662 ( .A(n45247), .B(n45246), .C(n45245), .D(n45244), .Y(n45252)
         );
  AOI21XL U32663 ( .A0(n48300), .A1(net209603), .B0(net209627), .Y(n48324) );
  NAND3XL U32664 ( .A(net209602), .B(net209603), .C(net209604), .Y(n48314) );
  NAND2XL U32665 ( .A(n48312), .B(n48307), .Y(n47731) );
  XOR2X1 U32666 ( .A(n34361), .B(n36875), .Y(n45152) );
  XOR2X1 U32667 ( .A(n36736), .B(n34314), .Y(n47299) );
  XOR2X1 U32668 ( .A(n36736), .B(n34290), .Y(n47331) );
  XOR2X1 U32669 ( .A(n41333), .B(n34397), .Y(n46589) );
  CLKINVX8 U32670 ( .A(net209919), .Y(net212238) );
  XOR2X1 U32671 ( .A(n34269), .B(n41281), .Y(n44864) );
  NOR2X1 U32672 ( .A(n48437), .B(n48436), .Y(n48438) );
  NOR2X1 U32673 ( .A(n47490), .B(net209287), .Y(n47500) );
  OAI21XL U32674 ( .A0(n48178), .A1(n48177), .B0(net209873), .Y(n48181) );
  NOR2X4 U32675 ( .A(n47457), .B(net209341), .Y(n47467) );
  INVXL U32676 ( .A(n48467), .Y(n48469) );
  NOR2X8 U32677 ( .A(n47286), .B(n48467), .Y(n47290) );
  NAND4X8 U32678 ( .A(n46199), .B(n46198), .C(n46197), .D(n46196), .Y(n48467)
         );
  NAND2X8 U32679 ( .A(n37235), .B(n44962), .Y(n48151) );
  XOR2X1 U32680 ( .A(n34382), .B(n40039), .Y(n44956) );
  INVX1 U32681 ( .A(net219468), .Y(net259034) );
  NAND2X4 U32682 ( .A(net210479), .B(n46473), .Y(n48145) );
  INVX4 U32683 ( .A(net210580), .Y(net209333) );
  XOR2X1 U32684 ( .A(n34301), .B(n41281), .Y(n45389) );
  INVXL U32685 ( .A(n48439), .Y(n48440) );
  NOR2X6 U32686 ( .A(n10395), .B(n44188), .Y(n44192) );
  INVXL U32687 ( .A(n10395), .Y(net209547) );
  NAND2XL U32688 ( .A(n11770), .B(n10395), .Y(n11769) );
  XNOR2X1 U32689 ( .A(n36851), .B(n34384), .Y(n46480) );
  AOI21X1 U32690 ( .A0(n48176), .A1(n48175), .B0(n48174), .Y(n48177) );
  NAND2X1 U32691 ( .A(n34398), .B(n41368), .Y(n41369) );
  AOI21XL U32692 ( .A0(n48442), .A1(n48441), .B0(n48440), .Y(n48444) );
  XOR2X1 U32693 ( .A(n34358), .B(net219310), .Y(n45118) );
  XOR2X1 U32694 ( .A(n41297), .B(n34358), .Y(n46490) );
  NOR2X4 U32695 ( .A(net210616), .B(net210617), .Y(n47764) );
  XOR2X1 U32696 ( .A(n34390), .B(net219330), .Y(n44920) );
  AOI21XL U32697 ( .A0(n48010), .A1(n48009), .B0(n48008), .Y(n48013) );
  NAND2XL U32698 ( .A(n48009), .B(n48005), .Y(n47977) );
  NOR4X2 U32699 ( .A(n44802), .B(n44801), .C(n44800), .D(n44799), .Y(n44813)
         );
  NAND3X1 U32700 ( .A(net210699), .B(n48147), .C(net209919), .Y(n47713) );
  AOI21XL U32701 ( .A0(net209622), .A1(net209623), .B0(net209624), .Y(n48304)
         );
  NOR4X2 U32702 ( .A(n44837), .B(n44836), .C(n44835), .D(n44834), .Y(n44840)
         );
  XNOR2XL U32703 ( .A(n36748), .B(n34388), .Y(n47691) );
  XOR2X1 U32704 ( .A(n36768), .B(n34313), .Y(n47297) );
  XOR2XL U32705 ( .A(n42066), .B(n41321), .Y(n45060) );
  XNOR2X1 U32706 ( .A(n36735), .B(n34378), .Y(n47654) );
  XNOR2XL U32707 ( .A(n36735), .B(n34106), .Y(n47560) );
  OR4X4 U32708 ( .A(n45066), .B(n45065), .C(n45064), .D(n45063), .Y(n41709) );
  XOR2X1 U32709 ( .A(n42080), .B(n41321), .Y(n45401) );
  XOR2X1 U32710 ( .A(n42096), .B(n41321), .Y(n43940) );
  NOR2X6 U32711 ( .A(n45367), .B(net209602), .Y(n45377) );
  XOR2X1 U32712 ( .A(n34294), .B(net219330), .Y(n45357) );
  NOR2X4 U32713 ( .A(n11148), .B(n47291), .Y(net211152) );
  NOR2X4 U32714 ( .A(n43820), .B(net209565), .Y(n43824) );
  XOR2X1 U32715 ( .A(n34341), .B(n41283), .Y(n45179) );
  NOR2X4 U32716 ( .A(n44784), .B(net213687), .Y(n44794) );
  NAND4X4 U32717 ( .A(n44794), .B(n44793), .C(n44792), .D(n44791), .Y(
        net209927) );
  XOR2X1 U32718 ( .A(n36733), .B(n34394), .Y(n47703) );
  NOR2X2 U32719 ( .A(net171547), .B(net171546), .Y(n11431) );
  BUFX20 U32720 ( .A(n42475), .Y(n42471) );
  NOR2X2 U32721 ( .A(n47380), .B(net209301), .Y(n47390) );
  XOR2X1 U32722 ( .A(n34418), .B(n42706), .Y(n45004) );
  XOR2X1 U32723 ( .A(n34262), .B(n40039), .Y(n44805) );
  NOR2X8 U32724 ( .A(n45157), .B(n48312), .Y(n45167) );
  NOR4X4 U32725 ( .A(n44972), .B(n44971), .C(n44970), .D(n44969), .Y(n44983)
         );
  XOR2X1 U32726 ( .A(n34362), .B(n42670), .Y(n44971) );
  XOR2X1 U32727 ( .A(n34333), .B(n41282), .Y(n45428) );
  NAND2X1 U32728 ( .A(n9657), .B(n41218), .Y(n41219) );
  INVX1 U32729 ( .A(n42669), .Y(n41218) );
  NAND2X2 U32730 ( .A(n41219), .B(n41220), .Y(n45242) );
  INVX1 U32731 ( .A(net209605), .Y(net210668) );
  INVX1 U32732 ( .A(n48465), .Y(n48428) );
  INVX2 U32733 ( .A(n48130), .Y(n48131) );
  NOR2XL U32734 ( .A(n47557), .B(n48465), .Y(n47561) );
  NOR2X6 U32735 ( .A(n46205), .B(n48130), .Y(n46209) );
  XOR2X1 U32736 ( .A(n42584), .B(n42061), .Y(n44033) );
  XOR2X1 U32737 ( .A(n34348), .B(n36871), .Y(n45209) );
  XOR2XL U32738 ( .A(n34316), .B(n36861), .Y(n45441) );
  NAND2X1 U32739 ( .A(n41345), .B(net219330), .Y(n41347) );
  AOI31XL U32740 ( .A0(n48450), .A1(n48449), .A2(net209320), .B0(n48448), .Y(
        n48454) );
  NOR2X8 U32741 ( .A(n46544), .B(n48149), .Y(n46554) );
  NAND4X8 U32742 ( .A(n45167), .B(n45166), .C(n45165), .D(n45164), .Y(n48158)
         );
  INVXL U32743 ( .A(n48449), .Y(n48447) );
  NOR4X1 U32744 ( .A(n45223), .B(n45222), .C(n45221), .D(n45220), .Y(n45224)
         );
  NAND2X1 U32745 ( .A(n48151), .B(n48149), .Y(net210698) );
  XOR2X1 U32746 ( .A(n34431), .B(n36900), .Y(n45026) );
  CLKINVX8 U32747 ( .A(n48305), .Y(n44962) );
  AOI21X2 U32748 ( .A0(n48388), .A1(n12490), .B0(net171119), .Y(n48389) );
  OAI2BB1X4 U32749 ( .A0N(n12449), .A1N(n41740), .B0(n11626), .Y(n48411) );
  AO21X4 U32750 ( .A0(n48410), .A1(n12452), .B0(net209455), .Y(n41740) );
  OAI21X4 U32751 ( .A0(n48397), .A1(n48396), .B0(net209476), .Y(n48398) );
  AOI21X1 U32752 ( .A0(n48281), .A1(n11688), .B0(net209663), .Y(n48386) );
  OAI21X1 U32753 ( .A0(n48275), .A1(n48274), .B0(n11709), .Y(n48276) );
  AOI21X1 U32754 ( .A0(n11711), .A1(net209675), .B0(net209676), .Y(n48274) );
  XOR2X1 U32755 ( .A(n34369), .B(n36875), .Y(n44980) );
  XOR2X1 U32756 ( .A(n34370), .B(n42705), .Y(n44979) );
  XOR2X1 U32757 ( .A(n34389), .B(n42628), .Y(n44883) );
  NOR2X4 U32758 ( .A(n46260), .B(n48179), .Y(n46270) );
  NAND4X4 U32759 ( .A(n44101), .B(n44100), .C(n44099), .D(n44098), .Y(n48179)
         );
  NOR2X4 U32760 ( .A(n47634), .B(n48443), .Y(n47644) );
  NAND2X6 U32761 ( .A(n41211), .B(n11638), .Y(n11632) );
  OR2X8 U32762 ( .A(net171474), .B(n48547), .Y(n41240) );
  AOI21X2 U32763 ( .A0(n48542), .A1(n11017), .B0(net209165), .Y(n48543) );
  AO21X4 U32764 ( .A0(n48424), .A1(n12324), .B0(n48423), .Y(n41782) );
  XOR2X1 U32765 ( .A(n34432), .B(net219434), .Y(n45034) );
  OAI2BB1X1 U32766 ( .A0N(net210233), .A1N(net210148), .B0(n10044), .Y(n47970)
         );
  NAND2X2 U32767 ( .A(n41234), .B(net219468), .Y(n41236) );
  NOR2X2 U32768 ( .A(n47446), .B(net209313), .Y(n47456) );
  NAND2X4 U32769 ( .A(n41206), .B(n41207), .Y(n45278) );
  BUFX16 U32770 ( .A(n42475), .Y(n42470) );
  NAND2X2 U32771 ( .A(n11147), .B(n11149), .Y(n48468) );
  NOR2X4 U32772 ( .A(n43829), .B(n48293), .Y(n43833) );
  NOR2X2 U32773 ( .A(net210476), .B(net210665), .Y(n41363) );
  XOR2X1 U32774 ( .A(n9659), .B(n41319), .Y(n45243) );
  XOR2X1 U32775 ( .A(n41810), .B(n42607), .Y(n44911) );
  XOR2X1 U32776 ( .A(n34381), .B(n41281), .Y(n44957) );
  XNOR2XL U32777 ( .A(n50800), .B(net258262), .Y(n26552) );
  XNOR2XL U32778 ( .A(n50814), .B(n40039), .Y(n26281) );
  XNOR2XL U32779 ( .A(n50854), .B(net219336), .Y(n30132) );
  XNOR2XL U32780 ( .A(n50828), .B(net219310), .Y(n26101) );
  XNOR2XL U32781 ( .A(n50844), .B(net258262), .Y(n29832) );
  XNOR2XL U32782 ( .A(n50981), .B(net219310), .Y(n29380) );
  XOR2X1 U32783 ( .A(n34351), .B(n36894), .Y(n45206) );
  XOR2X1 U32784 ( .A(n34349), .B(n41281), .Y(n45208) );
  XNOR2X1 U32785 ( .A(n34376), .B(n42592), .Y(n41654) );
  XNOR2X1 U32786 ( .A(n41811), .B(n42605), .Y(n41653) );
  OAI211XL U32787 ( .A0(n48447), .A1(net209323), .B0(n48446), .C0(net209325),
        .Y(n48448) );
  AOI21X1 U32788 ( .A0(n47970), .A1(n10045), .B0(net151670), .Y(n47971) );
  NAND3XL U32789 ( .A(n13014), .B(n11442), .C(n10045), .Y(n48041) );
  XOR2X1 U32790 ( .A(n34357), .B(n41282), .Y(n45119) );
  XOR2X1 U32791 ( .A(n34350), .B(n42534), .Y(n45158) );
  NOR2X6 U32792 ( .A(n47552), .B(n48426), .Y(n47556) );
  NAND4X4 U32793 ( .A(n43874), .B(n43873), .C(n43872), .D(n43871), .Y(n48335)
         );
  NOR4X2 U32794 ( .A(n43858), .B(n43857), .C(n43856), .D(n43855), .Y(n43874)
         );
  NOR3X4 U32795 ( .A(n45075), .B(n41711), .C(n45076), .Y(n45077) );
  XOR2X1 U32796 ( .A(n41798), .B(n42692), .Y(n45075) );
  XOR2X1 U32797 ( .A(n42064), .B(n36880), .Y(n45076) );
  NOR2X1 U32798 ( .A(n11140), .B(n47025), .Y(net211508) );
  NOR2X4 U32799 ( .A(n47435), .B(net209344), .Y(n47445) );
  XOR2X1 U32800 ( .A(n34265), .B(n41319), .Y(n45327) );
  CLKXOR2X2 U32801 ( .A(n41818), .B(n42523), .Y(n45455) );
  XOR2X1 U32802 ( .A(n41811), .B(n36892), .Y(n44974) );
  NAND4X4 U32803 ( .A(n46482), .B(n46481), .C(n46480), .D(n46479), .Y(n46488)
         );
  AOI21X4 U32804 ( .A0(n47747), .A1(n47746), .B0(net210639), .Y(n47749) );
  XOR2X1 U32805 ( .A(n34365), .B(n41281), .Y(n45148) );
  NOR4X2 U32806 ( .A(n44917), .B(n44916), .C(n44915), .D(n44914), .Y(n44928)
         );
  XNOR2XL U32807 ( .A(n50578), .B(n41380), .Y(n28054) );
  NOR2X8 U32808 ( .A(n46354), .B(net209894), .Y(n46364) );
  NAND2XL U32809 ( .A(net209894), .B(n48159), .Y(n48162) );
  NOR4X2 U32810 ( .A(n44105), .B(n44104), .C(n44103), .D(n44102), .Y(n44121)
         );
  XOR2X1 U32811 ( .A(n41832), .B(n36898), .Y(n44111) );
  XOR2X1 U32812 ( .A(n41812), .B(n36897), .Y(n45146) );
  NOR2X1 U32813 ( .A(n47562), .B(n48427), .Y(n47566) );
  NAND4X4 U32814 ( .A(n46220), .B(n46219), .C(n46218), .D(n46217), .Y(n48427)
         );
  NOR4X2 U32815 ( .A(n45404), .B(n45403), .C(n45402), .D(n45401), .Y(n45405)
         );
  XOR2X1 U32816 ( .A(n34166), .B(net219314), .Y(n43958) );
  XOR2X1 U32817 ( .A(n34361), .B(n41319), .Y(n44972) );
  NAND2XL U32818 ( .A(net209605), .B(net209606), .Y(n48315) );
  XOR2X1 U32819 ( .A(n34273), .B(n34435), .Y(n45335) );
  INVXL U32820 ( .A(n48149), .Y(n48150) );
  XOR2X1 U32821 ( .A(n34273), .B(n42684), .Y(n45296) );
  OAI2BB1X1 U32822 ( .A0N(n48039), .A1N(n48038), .B0(n48037), .Y(n48044) );
  NOR2X2 U32823 ( .A(n47601), .B(n48439), .Y(n47611) );
  XOR2X1 U32824 ( .A(n34397), .B(n41283), .Y(n44891) );
  XNOR2XL U32825 ( .A(n34264), .B(n42505), .Y(n45345) );
  XOR2X1 U32826 ( .A(n34326), .B(n42533), .Y(n45187) );
  XOR2X1 U32827 ( .A(n34254), .B(n42533), .Y(n44874) );
  NAND3X2 U32828 ( .A(n10585), .B(n12089), .C(n12090), .Y(n12088) );
  XOR2X1 U32829 ( .A(n41800), .B(n42627), .Y(n45015) );
  NOR2X6 U32830 ( .A(n46434), .B(net209927), .Y(n46444) );
  CLKINVX3 U32831 ( .A(n42510), .Y(n42502) );
  NOR2X6 U32832 ( .A(n41635), .B(net171421), .Y(n11106) );
  NAND4X4 U32833 ( .A(n44703), .B(n44702), .C(n44701), .D(n44700), .Y(n48172)
         );
  XOR2X1 U32834 ( .A(n34238), .B(net219314), .Y(n44683) );
  XOR2X1 U32835 ( .A(n34301), .B(n42624), .Y(n45495) );
  OAI21XL U32836 ( .A0(net210211), .A1(n47986), .B0(net210213), .Y(n47987) );
  NOR4X1 U32837 ( .A(n44051), .B(n44050), .C(n44049), .D(n44048), .Y(n44057)
         );
  NOR2X2 U32838 ( .A(n47510), .B(net209284), .Y(n47520) );
  XOR2X1 U32839 ( .A(n34182), .B(net219324), .Y(n44050) );
  XOR2X1 U32840 ( .A(n34232), .B(n34450), .Y(n44673) );
  NOR2X6 U32841 ( .A(n46445), .B(net209893), .Y(n46455) );
  NOR4X2 U32842 ( .A(n44082), .B(n44081), .C(n44080), .D(n44079), .Y(n44088)
         );
  XOR2X1 U32843 ( .A(n41822), .B(n42595), .Y(n45290) );
  OAI21X1 U32844 ( .A0(net209347), .A1(n48430), .B0(n11148), .Y(n48432) );
  XOR2X1 U32845 ( .A(n34281), .B(n36903), .Y(n45354) );
  NOR2X4 U32846 ( .A(n47479), .B(net209291), .Y(n47489) );
  XOR2X1 U32847 ( .A(n36721), .B(n34397), .Y(n47699) );
  NOR4X2 U32848 ( .A(n27598), .B(n27599), .C(n27600), .D(n27601), .Y(net215465) );
  NAND4X4 U32849 ( .A(n44168), .B(n44167), .C(n44166), .D(n44165), .Y(n12747)
         );
  NOR4X2 U32850 ( .A(n28083), .B(n28084), .C(n28085), .D(n28086), .Y(n43816)
         );
  NAND4X2 U32851 ( .A(n43817), .B(n43816), .C(n43815), .D(n43814), .Y(
        net210460) );
  NOR2X4 U32852 ( .A(n11147), .B(n46992), .Y(n46996) );
  CLKINVX8 U32853 ( .A(n12976), .Y(net151670) );
  NOR4X2 U32854 ( .A(n44829), .B(n44828), .C(n44827), .D(n44826), .Y(n44841)
         );
  XOR2X1 U32855 ( .A(n41827), .B(n36819), .Y(n44827) );
  INVXL U32856 ( .A(net210222), .Y(net210221) );
  OAI31X2 U32857 ( .A0(n11675), .A1(net171119), .A2(net171129), .B0(net151263),
        .Y(n11674) );
  XOR2X1 U32858 ( .A(n41814), .B(n42597), .Y(n45198) );
  OR4X8 U32859 ( .A(n41705), .B(n41706), .C(n41707), .D(n41652), .Y(n48305) );
  OAI211X2 U32860 ( .A0(n11037), .A1(n11038), .B0(n11039), .C0(n11040), .Y(
        n11036) );
  OAI21X4 U32861 ( .A0(n36936), .A1(n47761), .B0(n47760), .Y(n47763) );
  NOR4X2 U32862 ( .A(n45002), .B(n45001), .C(n45000), .D(n44999), .Y(n45023)
         );
  XNOR2X1 U32863 ( .A(n34369), .B(n42579), .Y(n44932) );
  XOR2X1 U32864 ( .A(n34305), .B(n42717), .Y(n45507) );
  CLKINVX6 U32865 ( .A(n47705), .Y(n48437) );
  XOR2X1 U32866 ( .A(n34417), .B(n36905), .Y(n45027) );
  NAND4X4 U32867 ( .A(n43947), .B(n43946), .C(n43945), .D(n43944), .Y(n48182)
         );
  XOR2X1 U32868 ( .A(n34174), .B(n36870), .Y(n43927) );
  XOR2X1 U32869 ( .A(n41835), .B(n36893), .Y(n43926) );
  XOR2X1 U32870 ( .A(n34290), .B(n42558), .Y(n45518) );
  NOR2X4 U32871 ( .A(n44153), .B(n48319), .Y(n44163) );
  OAI211X2 U32872 ( .A0(n10093), .A1(n50116), .B0(n11672), .C0(n11673), .Y(
        n11670) );
  AOI21X4 U32873 ( .A0(n47743), .A1(n47742), .B0(net210646), .Y(n47745) );
  OAI21X4 U32874 ( .A0(n47732), .A1(n47731), .B0(net210659), .Y(n47734) );
  AOI21X4 U32875 ( .A0(n47730), .A1(n47729), .B0(n47728), .Y(n47732) );
  INVX3 U32876 ( .A(n11674), .Y(n50116) );
  NOR2X2 U32877 ( .A(n47293), .B(n48446), .Y(n47303) );
  NOR4X2 U32878 ( .A(n44684), .B(n44683), .C(n44682), .D(n44681), .Y(n44690)
         );
  XNOR2X1 U32879 ( .A(n34385), .B(n42579), .Y(n45100) );
  NOR2X4 U32880 ( .A(n12344), .B(n47002), .Y(n47006) );
  XOR2X1 U32881 ( .A(n41823), .B(n42597), .Y(n45321) );
  NOR2X4 U32882 ( .A(n47017), .B(net209267), .Y(n47021) );
  NAND2XL U32883 ( .A(net209267), .B(n12344), .Y(n48431) );
  NAND4X4 U32884 ( .A(n44186), .B(n44185), .C(n44184), .D(n44183), .Y(n12089)
         );
  NOR2X2 U32885 ( .A(net151672), .B(net151670), .Y(n11437) );
  XOR2X1 U32886 ( .A(n41825), .B(n42605), .Y(n44796) );
  XNOR2X1 U32887 ( .A(n50335), .B(n42670), .Y(n26819) );
  OAI21X2 U32888 ( .A0(n37253), .A1(net210109), .B0(n12942), .Y(n48073) );
  XNOR2X1 U32889 ( .A(n50539), .B(n41319), .Y(n26820) );
  AOI21X1 U32890 ( .A0(n48076), .A1(n10752), .B0(n39636), .Y(n48077) );
  OAI211X2 U32891 ( .A0(n11047), .A1(n11048), .B0(n11049), .C0(n11050), .Y(
        n11043) );
  NAND2X6 U32892 ( .A(n41651), .B(net151599), .Y(n11119) );
  XNOR2X1 U32893 ( .A(n34338), .B(n41642), .Y(n41727) );
  OAI211X2 U32894 ( .A0(n12091), .A1(n10182), .B0(n10184), .C0(n39304), .Y(
        n12090) );
  OAI211X2 U32895 ( .A0(n11995), .A1(n10522), .B0(n10520), .C0(n10519), .Y(
        n11993) );
  AOI211X2 U32896 ( .A0(n11980), .A1(n11981), .B0(net209760), .C0(net151495),
        .Y(n11974) );
  OAI211X2 U32897 ( .A0(n12046), .A1(n12047), .B0(n40392), .C0(n12049), .Y(
        n12043) );
  XNOR2X1 U32898 ( .A(n34353), .B(n34435), .Y(n41730) );
  XNOR2X1 U32899 ( .A(n34354), .B(n42706), .Y(n41731) );
  OAI211X2 U32900 ( .A0(n11356), .A1(n11357), .B0(n11358), .C0(n11359), .Y(
        n11353) );
  NAND2X2 U32901 ( .A(n48020), .B(n48018), .Y(n47759) );
  AOI31X2 U32902 ( .A0(n11057), .A1(n11058), .A2(n11059), .B0(n39488), .Y(
        n11053) );
  OAI21X4 U32903 ( .A0(net171114), .A1(n48399), .B0(n10339), .Y(n48400) );
  OAI21X4 U32904 ( .A0(net171129), .A1(n48389), .B0(n12488), .Y(n48390) );
  OAI21X1 U32905 ( .A0(net209664), .A1(n48280), .B0(n11694), .Y(n48281) );
  AOI21X4 U32906 ( .A0(n48398), .A1(n12474), .B0(net171319), .Y(n48399) );
  XOR2X1 U32907 ( .A(n34329), .B(n42576), .Y(n45221) );
  AOI211X2 U32908 ( .A0(n11053), .A1(n11054), .B0(net151458), .C0(net151473),
        .Y(n11047) );
  AOI211X2 U32909 ( .A0(n11067), .A1(n11068), .B0(net171456), .C0(net171453),
        .Y(n11061) );
  CLKINVX3 U32910 ( .A(n42623), .Y(n42613) );
  NAND4X4 U32911 ( .A(n43998), .B(n43997), .C(n43996), .D(n43995), .Y(n48289)
         );
  NOR2X2 U32912 ( .A(n47567), .B(n48464), .Y(n47577) );
  NOR2X4 U32913 ( .A(n46294), .B(n48166), .Y(n46304) );
  NAND2X1 U32914 ( .A(n34396), .B(n41388), .Y(n41389) );
  XOR2X1 U32915 ( .A(n41828), .B(n42605), .Y(n44674) );
  XOR2X1 U32916 ( .A(n41835), .B(n42605), .Y(n44041) );
  XOR2X1 U32917 ( .A(n41836), .B(n42605), .Y(n43918) );
  XOR2X1 U32918 ( .A(n41832), .B(n42605), .Y(n44134) );
  NAND3XL U32919 ( .A(n48151), .B(n48145), .C(net209919), .Y(n48154) );
  NOR2X4 U32920 ( .A(n46271), .B(n48185), .Y(n46281) );
  INVXL U32921 ( .A(net209312), .Y(net209342) );
  NAND4BX4 U32922 ( .AN(n46488), .B(n46487), .C(n46486), .D(net209620), .Y(
        n48441) );
  OAI21X4 U32923 ( .A0(net171156), .A1(n48271), .B0(net260431), .Y(n48272) );
  OAI21X4 U32924 ( .A0(net209750), .A1(n48264), .B0(net260277), .Y(n48265) );
  OAI21X4 U32925 ( .A0(n48247), .A1(n48246), .B0(n12799), .Y(n48248) );
  AOI21X4 U32926 ( .A0(n48254), .A1(n10520), .B0(net209772), .Y(n48255) );
  OAI21X4 U32927 ( .A0(net209773), .A1(n48253), .B0(n12672), .Y(n48254) );
  AOI21X2 U32928 ( .A0(n48117), .A1(n12711), .B0(net209969), .Y(n48118) );
  XNOR2X1 U32929 ( .A(n50952), .B(n42618), .Y(n25012) );
  OAI21X4 U32930 ( .A0(net209764), .A1(n48257), .B0(n11991), .Y(n48258) );
  AOI21X2 U32931 ( .A0(n48256), .A1(net209767), .B0(net209768), .Y(n48257) );
  AOI211X2 U32932 ( .A0(n11342), .A1(n11343), .B0(net171532), .C0(n37240), .Y(
        n11339) );
  XOR2X1 U32933 ( .A(n34292), .B(n41385), .Y(n45359) );
  INVX4 U32934 ( .A(n11122), .Y(n41650) );
  BUFX20 U32935 ( .A(n42648), .Y(n42658) );
  NAND3X6 U32936 ( .A(n41650), .B(net211197), .C(net209249), .Y(n41651) );
  AOI21X4 U32937 ( .A0(n48544), .A1(n40395), .B0(net209161), .Y(n48545) );
  OAI21X4 U32938 ( .A0(n39485), .A1(n48543), .B0(n11016), .Y(n48544) );
  OAI21X1 U32939 ( .A0(n48490), .A1(n48489), .B0(n48488), .Y(n48496) );
  OAI21X4 U32940 ( .A0(net209172), .A1(n48537), .B0(n11031), .Y(n48538) );
  AOI21X4 U32941 ( .A0(n48536), .A1(n40390), .B0(net209175), .Y(n48537) );
  AOI21X4 U32942 ( .A0(n48552), .A1(n10990), .B0(net209144), .Y(net209142) );
  NAND4X4 U32943 ( .A(n46209), .B(n46208), .C(n46207), .D(n46206), .Y(n48465)
         );
  XOR2X1 U32944 ( .A(n36838), .B(n34402), .Y(n46555) );
  XOR2X1 U32945 ( .A(n36840), .B(n34378), .Y(n46485) );
  XOR2X1 U32946 ( .A(n36844), .B(n34306), .Y(n46316) );
  XOR2X1 U32947 ( .A(n36845), .B(n34354), .Y(n46495) );
  AOI21X4 U32948 ( .A0(n47764), .A1(n47763), .B0(n47762), .Y(n47765) );
  NOR4X2 U32949 ( .A(n44990), .B(n44989), .C(n44988), .D(n44987), .Y(n44991)
         );
  XOR2X1 U32950 ( .A(n34209), .B(n42579), .Y(n44666) );
  CLKINVX6 U32951 ( .A(n11008), .Y(n50089) );
  OAI2BB1X4 U32952 ( .A0N(n11316), .A1N(n41692), .B0(n11317), .Y(n48109) );
  OAI21X4 U32953 ( .A0(n47960), .A1(n47959), .B0(n11510), .Y(n47962) );
  AOI21X1 U32954 ( .A0(n47962), .A1(n11509), .B0(n47961), .Y(n48092) );
  AOI211X2 U32955 ( .A0(n12050), .A1(n12051), .B0(net171247), .C0(net171245),
        .Y(n12046) );
  OAI211X2 U32956 ( .A0(n11986), .A1(n11987), .B0(n11988), .C0(n11989), .Y(
        n11981) );
  NOR3X2 U32957 ( .A(n11996), .B(net171136), .C(net171139), .Y(n11995) );
  NOR2X1 U32958 ( .A(net209885), .B(net210702), .Y(n47724) );
  AOI211X2 U32959 ( .A0(n11019), .A1(n11020), .B0(n39487), .C0(net171472), .Y(
        n11013) );
  AND3X8 U32960 ( .A(n50089), .B(n11006), .C(n11007), .Y(n11003) );
  OAI21X4 U32961 ( .A0(n47779), .A1(n47778), .B0(net234488), .Y(n47781) );
  OAI211X2 U32962 ( .A0(n11013), .A1(n11014), .B0(n11015), .C0(n11016), .Y(
        n11010) );
  OAI21X4 U32963 ( .A0(n47741), .A1(n47740), .B0(n47739), .Y(n47742) );
  INVX12 U32964 ( .A(net210477), .Y(net209620) );
  OAI211X2 U32965 ( .A0(n50115), .A1(n11667), .B0(n10090), .C0(n10089), .Y(
        n11663) );
  INVX3 U32966 ( .A(n11670), .Y(n50115) );
  OAI21X4 U32967 ( .A0(n47745), .A1(net210641), .B0(n47744), .Y(n47746) );
  AOI211X2 U32968 ( .A0(n11713), .A1(n11714), .B0(net151401), .C0(net209675),
        .Y(n11707) );
  OAI211X2 U32969 ( .A0(n11659), .A1(n11660), .B0(n10336), .C0(n10339), .Y(
        n11654) );
  AOI211X2 U32970 ( .A0(net151265), .A1(n11663), .B0(net171113), .C0(net151253), .Y(n11659) );
  AOI211X2 U32971 ( .A0(n11009), .A1(n11010), .B0(net171471), .C0(net171470),
        .Y(n11008) );
  NAND3X6 U32972 ( .A(n11023), .B(n11024), .C(n11025), .Y(n11020) );
  NAND4X4 U32973 ( .A(n45408), .B(n45407), .C(n45406), .D(n45405), .Y(n48137)
         );
  OAI211X2 U32974 ( .A0(n11322), .A1(n11323), .B0(n11324), .C0(n11325), .Y(
        n11319) );
  OAI211X2 U32975 ( .A0(n11346), .A1(n11347), .B0(n11348), .C0(n11349), .Y(
        n11343) );
  NAND2X2 U32976 ( .A(n48028), .B(n48030), .Y(n47771) );
  AOI21X4 U32977 ( .A0(n47782), .A1(n47781), .B0(n47780), .Y(n47783) );
  XOR2X1 U32978 ( .A(n34176), .B(net219460), .Y(n43925) );
  AOI211X2 U32979 ( .A0(n11390), .A1(n11391), .B0(n39900), .C0(net151847), .Y(
        n11384) );
  NOR4X2 U32980 ( .A(n45231), .B(n45230), .C(n45229), .D(n45228), .Y(n45256)
         );
  AOI211X2 U32981 ( .A0(n11042), .A1(n11043), .B0(net171467), .C0(net151477),
        .Y(n11037) );
  OAI211X2 U32982 ( .A0(n11026), .A1(n11027), .B0(n40399), .C0(n11029), .Y(
        n11025) );
  XOR2X1 U32983 ( .A(n34326), .B(n40039), .Y(n45447) );
  AOI21X4 U32984 ( .A0(n48100), .A1(n48099), .B0(n41735), .Y(n48101) );
  INVX1 U32985 ( .A(n47980), .Y(n47983) );
  OAI21X2 U32986 ( .A0(n48045), .A1(n48044), .B0(n48043), .Y(n48051) );
  AOI211X2 U32987 ( .A0(n11328), .A1(n11329), .B0(net151445), .C0(net151448),
        .Y(n11322) );
  AOI211X2 U32988 ( .A0(n12018), .A1(n12019), .B0(net171201), .C0(net171200),
        .Y(n12012) );
  AOI211X2 U32989 ( .A0(net151456), .A1(n11993), .B0(net209768), .C0(net171117), .Y(n11986) );
  OAI211X2 U32990 ( .A0(n12060), .A1(n12061), .B0(n12062), .C0(n12063), .Y(
        n12057) );
  AOI211X2 U32991 ( .A0(n12066), .A1(n12067), .B0(n49508), .C0(n49509), .Y(
        n12060) );
  OAI211X2 U32992 ( .A0(n12012), .A1(n12013), .B0(n12014), .C0(n12015), .Y(
        n12009) );
  AOI211X2 U32993 ( .A0(n12042), .A1(n12043), .B0(net171307), .C0(net171304),
        .Y(n12040) );
  OAI2BB1X4 U32994 ( .A0N(n11621), .A1N(n41739), .B0(n11620), .Y(n48412) );
  AO21X4 U32995 ( .A0(n48411), .A1(n11625), .B0(n39702), .Y(n41739) );
  AOI21X4 U32996 ( .A0(n48412), .A1(n10425), .B0(net171146), .Y(net209446) );
  OAI21X4 U32997 ( .A0(net171321), .A1(n48409), .B0(n12455), .Y(n48410) );
  AOI21X4 U32998 ( .A0(n48408), .A1(n12457), .B0(net171098), .Y(n48409) );
  OAI21X2 U32999 ( .A0(net171101), .A1(n48404), .B0(n11645), .Y(n48405) );
  OAI21X4 U33000 ( .A0(net171152), .A1(n48273), .B0(n10483), .Y(net209732) );
  AOI21X4 U33001 ( .A0(n48272), .A1(n10485), .B0(net209736), .Y(n48273) );
  AOI21X2 U33002 ( .A0(n48218), .A1(n48217), .B0(n48216), .Y(n48233) );
  NOR2X4 U33003 ( .A(n10126), .B(n44187), .Y(net215433) );
  AOI211X2 U33004 ( .A0(n11689), .A1(n11690), .B0(net151327), .C0(net209664),
        .Y(n11683) );
  OAI211X2 U33005 ( .A0(n11695), .A1(n11696), .B0(n11697), .C0(n11698), .Y(
        n11690) );
  AOI211X2 U33006 ( .A0(n11734), .A1(n11735), .B0(net151356), .C0(net209517),
        .Y(n11729) );
  OAI211X2 U33007 ( .A0(n11729), .A1(n11730), .B0(n11731), .C0(n11732), .Y(
        n11726) );
  AOI211X2 U33008 ( .A0(n11679), .A1(n11680), .B0(net151261), .C0(net151258),
        .Y(n11675) );
  OAI211X2 U33009 ( .A0(n11683), .A1(n11684), .B0(n11685), .C0(n11686), .Y(
        n11680) );
  BUFX20 U33010 ( .A(n42666), .Y(n42659) );
  OAI211X2 U33011 ( .A0(n11647), .A1(n11648), .B0(n11649), .C0(n11650), .Y(
        n11642) );
  AOI211X2 U33012 ( .A0(n11653), .A1(n11654), .B0(net151271), .C0(net151270),
        .Y(n11647) );
  OAI2BB1X4 U33013 ( .A0N(n40400), .A1N(n41772), .B0(n11002), .Y(n48549) );
  OAI21X2 U33014 ( .A0(net171472), .A1(n48541), .B0(n12390), .Y(n48542) );
  AOI21X2 U33015 ( .A0(n48538), .A1(n40399), .B0(net209171), .Y(n48539) );
  OAI21X4 U33016 ( .A0(net171470), .A1(n48545), .B0(n12391), .Y(n48546) );
  AOI21X1 U33017 ( .A0(n48500), .A1(n10853), .B0(net209231), .Y(n48501) );
  OAI21X1 U33018 ( .A0(net209228), .A1(n48501), .B0(n40396), .Y(n48502) );
  NAND4X2 U33019 ( .A(n45653), .B(n45652), .C(n45651), .D(n45650), .Y(
        net209242) );
  AOI21X4 U33020 ( .A0(n41761), .A1(n47788), .B0(net210539), .Y(n47789) );
  AOI211X2 U33021 ( .A0(n11076), .A1(n11077), .B0(net171449), .C0(net171448),
        .Y(n11070) );
  AOI211X2 U33022 ( .A0(net151452), .A1(n11033), .B0(net171469), .C0(net209175), .Y(n11026) );
  NAND2XL U33023 ( .A(n42122), .B(n36917), .Y(n41200) );
  NAND2XL U33024 ( .A(n37246), .B(n42661), .Y(n41201) );
  NAND2X1 U33025 ( .A(n41200), .B(n41201), .Y(n27334) );
  NOR4X2 U33026 ( .A(n27331), .B(n27332), .C(n27333), .D(n27334), .Y(n44226)
         );
  INVXL U33027 ( .A(n48158), .Y(n41202) );
  NAND3XL U33028 ( .A(net209903), .B(net209900), .C(n48156), .Y(n48157) );
  OAI21X4 U33029 ( .A0(n48165), .A1(n48164), .B0(n48163), .Y(n48169) );
  AOI21X4 U33030 ( .A0(n48110), .A1(net210047), .B0(net238947), .Y(n48111) );
  XNOR2XL U33031 ( .A(n50974), .B(n36870), .Y(n26793) );
  XNOR2XL U33032 ( .A(n51188), .B(n41283), .Y(n26794) );
  XNOR2XL U33033 ( .A(n50760), .B(net219434), .Y(n26795) );
  NAND2XL U33034 ( .A(n51182), .B(n42628), .Y(n41208) );
  NAND2X1 U33035 ( .A(n33773), .B(n36803), .Y(n41209) );
  NAND2X1 U33036 ( .A(n41208), .B(n41209), .Y(n26876) );
  OR2X6 U33037 ( .A(n39491), .B(n48518), .Y(n41210) );
  AO21X4 U33038 ( .A0(n48519), .A1(n11073), .B0(net171458), .Y(n41695) );
  OA21X4 U33039 ( .A0(n11635), .A1(n11636), .B0(n11637), .Y(n41211) );
  AOI211X2 U33040 ( .A0(n11641), .A1(n11642), .B0(net151249), .C0(net151248),
        .Y(n11635) );
  OR2X6 U33041 ( .A(n47722), .B(net210682), .Y(n41212) );
  NAND2X6 U33042 ( .A(n41212), .B(net234527), .Y(n47723) );
  AOI21X4 U33043 ( .A0(n47721), .A1(n47720), .B0(n47719), .Y(n47722) );
  CLKAND2X2 U33044 ( .A(n48171), .B(n48173), .Y(net234527) );
  NAND2X8 U33045 ( .A(n10341), .B(n37014), .Y(n41213) );
  NAND2X6 U33046 ( .A(n41213), .B(n11657), .Y(n48401) );
  INVX1 U33047 ( .A(n10341), .Y(net171140) );
  CLKINVX1 U33048 ( .A(n12929), .Y(net151857) );
  OR3X4 U33049 ( .A(n11628), .B(net171098), .C(net171321), .Y(n41215) );
  AOI211X2 U33050 ( .A0(n11631), .A1(n11632), .B0(net151246), .C0(net151243),
        .Y(n11628) );
  NAND2X2 U33051 ( .A(n41216), .B(n11770), .Y(n48349) );
  AOI21X2 U33052 ( .A0(n48349), .A1(n10387), .B0(net209546), .Y(n48350) );
  NAND2X1 U33053 ( .A(n34242), .B(n41222), .Y(n41223) );
  NAND2XL U33054 ( .A(n41221), .B(n42559), .Y(n41224) );
  INVXL U33055 ( .A(n42559), .Y(n41222) );
  CLKINVX1 U33056 ( .A(n42573), .Y(n42559) );
  NOR4X2 U33057 ( .A(n44821), .B(n44820), .C(n44819), .D(n44818), .Y(n44822)
         );
  OA21X4 U33058 ( .A0(n12002), .A1(n12003), .B0(n12004), .Y(n41225) );
  NAND2X6 U33059 ( .A(n41225), .B(n12005), .Y(n11999) );
  AOI211X2 U33060 ( .A0(n12008), .A1(n12009), .B0(n39557), .C0(net171127), .Y(
        n12002) );
  NAND2X2 U33061 ( .A(n12006), .B(n12007), .Y(n12003) );
  NAND4X4 U33062 ( .A(n43254), .B(n43253), .C(n43252), .D(n43251), .Y(n12004)
         );
  NAND3X2 U33063 ( .A(n10996), .B(n10997), .C(n10998), .Y(n10994) );
  CLKINVX1 U33064 ( .A(n10807), .Y(net151503) );
  CLKINVX1 U33065 ( .A(n12959), .Y(net151601) );
  NAND2XL U33066 ( .A(n41227), .B(n42725), .Y(n41230) );
  INVXL U33067 ( .A(n36708), .Y(n41228) );
  NAND2X1 U33068 ( .A(n41232), .B(n41233), .Y(n44141) );
  NOR4X2 U33069 ( .A(n44868), .B(n44867), .C(n44866), .D(n44865), .Y(n44869)
         );
  OR2X6 U33070 ( .A(net210034), .B(n48115), .Y(net259031) );
  AOI21X4 U33071 ( .A0(n48114), .A1(n39345), .B0(net151514), .Y(n48115) );
  NAND2XL U33072 ( .A(n42161), .B(n41237), .Y(n41238) );
  NAND2XL U33073 ( .A(n37247), .B(n42655), .Y(n41239) );
  NAND2X1 U33074 ( .A(n41238), .B(n41239), .Y(n25199) );
  INVXL U33075 ( .A(n42655), .Y(n41237) );
  NAND2X6 U33076 ( .A(n41240), .B(n10810), .Y(n48548) );
  AOI21X4 U33077 ( .A0(n48546), .A1(n11006), .B0(net209158), .Y(n48547) );
  AO21X4 U33078 ( .A0(n48548), .A1(n10274), .B0(net209155), .Y(n41772) );
  NOR2X2 U33079 ( .A(net209629), .B(n48299), .Y(n41241) );
  INVXL U33080 ( .A(net209631), .Y(net259019) );
  OR2X8 U33081 ( .A(n41241), .B(net259019), .Y(n48300) );
  INVXL U33082 ( .A(net209602), .Y(net209629) );
  NAND2XL U33083 ( .A(n50968), .B(n41647), .Y(n41242) );
  NAND2X1 U33084 ( .A(n33774), .B(n42621), .Y(n41243) );
  NAND2X1 U33085 ( .A(n41242), .B(n41243), .Y(n26875) );
  NAND2XL U33086 ( .A(n50310), .B(n42672), .Y(n41245) );
  NAND2X1 U33087 ( .A(n41244), .B(n36924), .Y(n41246) );
  NAND2X1 U33088 ( .A(n41245), .B(n41246), .Y(n24806) );
  INVXL U33089 ( .A(n50310), .Y(n41244) );
  XNOR2XL U33090 ( .A(n33810), .B(n42568), .Y(n43676) );
  NAND2XL U33091 ( .A(n50336), .B(n42674), .Y(n41248) );
  NAND2X1 U33092 ( .A(n41248), .B(n41249), .Y(n26879) );
  INVXL U33093 ( .A(n50336), .Y(n41247) );
  NAND2XL U33094 ( .A(n51367), .B(n42643), .Y(n41252) );
  NAND2X1 U33095 ( .A(n41250), .B(n41251), .Y(n41253) );
  NAND2X1 U33096 ( .A(n41252), .B(n41253), .Y(n28116) );
  INVXL U33097 ( .A(n51367), .Y(n41250) );
  INVXL U33098 ( .A(n42643), .Y(n41251) );
  NAND2X1 U33099 ( .A(n41863), .B(n36919), .Y(n41254) );
  NAND2XL U33100 ( .A(n37248), .B(n42607), .Y(n41255) );
  NAND2X1 U33101 ( .A(n41254), .B(n41255), .Y(n27330) );
  NOR4X2 U33102 ( .A(n27327), .B(n27328), .C(n27329), .D(n27330), .Y(n44227)
         );
  NAND2X1 U33103 ( .A(n50772), .B(net219468), .Y(n41256) );
  NAND2X1 U33104 ( .A(n34184), .B(net258961), .Y(n41260) );
  NAND2X1 U33105 ( .A(n41259), .B(net219450), .Y(n41261) );
  NAND2XL U33106 ( .A(n50757), .B(n36865), .Y(n41262) );
  NAND2X2 U33107 ( .A(n41262), .B(n41263), .Y(n26727) );
  NAND2XL U33108 ( .A(n51156), .B(n42633), .Y(n41264) );
  NAND2X1 U33109 ( .A(n33565), .B(n36804), .Y(n41265) );
  NAND2X1 U33110 ( .A(n41264), .B(n41265), .Y(n24803) );
  NAND2XL U33111 ( .A(n50514), .B(n36728), .Y(n41266) );
  NAND2X1 U33112 ( .A(n33561), .B(n36922), .Y(n41267) );
  NAND2X1 U33113 ( .A(n41266), .B(n41267), .Y(n24807) );
  NOR2X2 U33114 ( .A(n43891), .B(n37206), .Y(n43904) );
  XOR2XL U33115 ( .A(n42099), .B(n42651), .Y(n43891) );
  NAND4X4 U33116 ( .A(n43905), .B(n43904), .C(n43903), .D(n43902), .Y(n48288)
         );
  NAND2XL U33117 ( .A(n37249), .B(n36893), .Y(n41269) );
  NAND2X1 U33118 ( .A(n41268), .B(n41269), .Y(n29112) );
  NAND2XL U33119 ( .A(n50309), .B(n42712), .Y(n41274) );
  NAND2X1 U33120 ( .A(n41274), .B(n41275), .Y(n28122) );
  INVXL U33121 ( .A(n50309), .Y(n41273) );
  NAND2X6 U33122 ( .A(n41276), .B(n47725), .Y(n47726) );
  INVXL U33123 ( .A(net210675), .Y(net258903) );
  NAND2XL U33124 ( .A(n48182), .B(n48185), .Y(net210675) );
  AOI21X4 U33125 ( .A0(n36947), .A1(n47726), .B0(net210673), .Y(n12091) );
  NAND2X2 U33126 ( .A(n42064), .B(n36939), .Y(n41277) );
  OR2X6 U33127 ( .A(net209483), .B(n48391), .Y(n41279) );
  NAND2X6 U33128 ( .A(n41279), .B(n11672), .Y(n48392) );
  CLKINVX1 U33129 ( .A(n12482), .Y(net209483) );
  AOI21X4 U33130 ( .A0(n48390), .A1(n12485), .B0(net209486), .Y(n48391) );
  XOR2X1 U33131 ( .A(n34353), .B(n41379), .Y(n45144) );
  XOR2X1 U33132 ( .A(n34357), .B(n42625), .Y(n45140) );
  XNOR2X1 U33133 ( .A(n50313), .B(n42672), .Y(n24776) );
  XNOR2X1 U33134 ( .A(n50343), .B(n42707), .Y(n29023) );
  XOR2X1 U33135 ( .A(n41867), .B(n36899), .Y(n29323) );
  XOR2X1 U33136 ( .A(n41913), .B(n42600), .Y(n28113) );
  XNOR2X1 U33137 ( .A(n50786), .B(n42592), .Y(n27600) );
  NOR4X2 U33138 ( .A(n26875), .B(n26876), .C(n26877), .D(n26878), .Y(net215227) );
  XNOR2X1 U33139 ( .A(n51155), .B(n41282), .Y(n28119) );
  XOR2X1 U33140 ( .A(n42112), .B(n42663), .Y(n27605) );
  XOR2X1 U33141 ( .A(n34417), .B(n42575), .Y(n45283) );
  AOI211X2 U33142 ( .A0(n11437), .A1(n11438), .B0(net151708), .C0(net151711),
        .Y(n11435) );
  XNOR2X1 U33143 ( .A(n50315), .B(n36907), .Y(n24926) );
  XNOR2X1 U33144 ( .A(n51159), .B(n42631), .Y(n24773) );
  XNOR2X1 U33145 ( .A(n50368), .B(n42711), .Y(n27520) );
  NAND4X2 U33146 ( .A(n47203), .B(n47202), .C(n47201), .D(n47200), .Y(n12316)
         );
  OAI21X2 U33147 ( .A0(net209617), .A1(n48304), .B0(n48303), .Y(n48313) );
  NOR4X2 U33148 ( .A(n24776), .B(n24777), .C(n24778), .D(n24779), .Y(n44554)
         );
  XNOR2X1 U33149 ( .A(n50517), .B(n36905), .Y(n24777) );
  XOR2X1 U33150 ( .A(n41884), .B(n36893), .Y(n26886) );
  XNOR2X1 U33151 ( .A(n50311), .B(n42708), .Y(n24814) );
  XNOR2X1 U33152 ( .A(n50540), .B(n36905), .Y(n26880) );
  OAI211X2 U33153 ( .A0(n11768), .A1(n11769), .B0(n10387), .C0(n10383), .Y(
        n11765) );
  AOI211X2 U33154 ( .A0(n11771), .A1(n11772), .B0(net151340), .C0(net209549),
        .Y(n11768) );
  XNOR2X1 U33155 ( .A(n51369), .B(n42641), .Y(n24808) );
  AOI21X1 U33156 ( .A0(n48417), .A1(n11208), .B0(net171441), .Y(n48418) );
  AOI211X2 U33157 ( .A0(n11418), .A1(n11419), .B0(net151594), .C0(net151593),
        .Y(n11412) );
  INVX1 U33158 ( .A(net209814), .Y(net171245) );
  NAND4X4 U33159 ( .A(n44260), .B(n44259), .C(n44258), .D(n44257), .Y(
        net209814) );
  XNOR2X1 U33160 ( .A(n50728), .B(n36863), .Y(n24804) );
  NOR2X1 U33161 ( .A(n43999), .B(n48289), .Y(n44009) );
  XOR2X1 U33162 ( .A(n34427), .B(n42660), .Y(n45266) );
  OAI211X2 U33163 ( .A0(n11760), .A1(n40393), .B0(n11762), .C0(n11763), .Y(
        n11758) );
  AOI211X2 U33164 ( .A0(n11764), .A1(n11765), .B0(net209543), .C0(net151348),
        .Y(n11760) );
  XNOR2X1 U33165 ( .A(n50971), .B(n42615), .Y(n26725) );
  NAND2X1 U33166 ( .A(net209898), .B(net209894), .Y(n47716) );
  XOR2X1 U33167 ( .A(n42088), .B(n42658), .Y(n44647) );
  XOR2X1 U33168 ( .A(n9669), .B(n36871), .Y(n45268) );
  INVXL U33169 ( .A(net210442), .Y(net214016) );
  AOI21XL U33170 ( .A0(n48181), .A1(net209868), .B0(n48180), .Y(n48183) );
  AOI211X2 U33171 ( .A0(n11400), .A1(n11401), .B0(net151744), .C0(net151746),
        .Y(n11394) );
  NAND4BBX4 U33172 ( .AN(n46510), .BN(n41723), .C(n46509), .D(n48306), .Y(
        n48435) );
  NOR4X4 U33173 ( .A(n44017), .B(n44016), .C(n44015), .D(n44014), .Y(n44028)
         );
  XOR2X1 U33174 ( .A(n34140), .B(n42638), .Y(n44014) );
  XOR2X2 U33175 ( .A(n42070), .B(n42659), .Y(n44970) );
  XNOR2X1 U33176 ( .A(n51373), .B(n36867), .Y(n24958) );
  XOR2X1 U33177 ( .A(n34128), .B(net219450), .Y(n43845) );
  XOR2X1 U33178 ( .A(n42111), .B(n42662), .Y(n27575) );
  CLKBUFX4 U33179 ( .A(n42646), .Y(n42662) );
  XNOR2X1 U33180 ( .A(n50733), .B(n36865), .Y(n24924) );
  XNOR2X1 U33181 ( .A(n49510), .B(n42711), .Y(n27731) );
  XNOR2X1 U33182 ( .A(n50574), .B(n42724), .Y(n27581) );
  CLKINVX4 U33183 ( .A(n42726), .Y(n42724) );
  CLKINVX1 U33184 ( .A(n47716), .Y(n45519) );
  XNOR2X1 U33185 ( .A(n51372), .B(n36867), .Y(n24778) );
  XNOR2X1 U33186 ( .A(n49514), .B(n42618), .Y(n27719) );
  XOR2X1 U33187 ( .A(n41907), .B(n42608), .Y(n24955) );
  XOR2X1 U33188 ( .A(n34228), .B(n42637), .Y(n44677) );
  XOR2X1 U33189 ( .A(n42167), .B(n42663), .Y(n24779) );
  OAI211X2 U33190 ( .A0(n11739), .A1(n11740), .B0(n11741), .C0(n11742), .Y(
        n11738) );
  XOR2X1 U33191 ( .A(n34429), .B(n41283), .Y(n45025) );
  XNOR2X1 U33192 ( .A(n50733), .B(net258207), .Y(n24962) );
  XOR2X1 U33193 ( .A(n41852), .B(n42608), .Y(n27571) );
  XOR2X1 U33194 ( .A(n41907), .B(n36899), .Y(n24783) );
  XNOR2X1 U33195 ( .A(n50947), .B(n42618), .Y(n24922) );
  XOR2X1 U33196 ( .A(n42087), .B(n42658), .Y(n44678) );
  XOR2X1 U33197 ( .A(n34230), .B(n41284), .Y(n44675) );
  OAI21X1 U33198 ( .A0(net171418), .A1(n48503), .B0(n10845), .Y(n48508) );
  XOR2X1 U33199 ( .A(n42069), .B(n42659), .Y(n44951) );
  OAI211X2 U33200 ( .A0(n11412), .A1(n11413), .B0(n11414), .C0(n11415), .Y(
        n11407) );
  XNOR2X1 U33201 ( .A(n50314), .B(n42708), .Y(n24784) );
  XOR2X1 U33202 ( .A(n41839), .B(n42605), .Y(n44011) );
  XNOR2X1 U33203 ( .A(n50731), .B(n36863), .Y(n24774) );
  XNOR2X1 U33204 ( .A(n51214), .B(n41283), .Y(n27517) );
  XOR2X1 U33205 ( .A(n34330), .B(n42707), .Y(n45431) );
  XOR2X2 U33206 ( .A(n41812), .B(n42597), .Y(n44966) );
  AOI21X1 U33207 ( .A0(n48284), .A1(n11850), .B0(n48283), .Y(n48285) );
  NOR2X2 U33208 ( .A(n45398), .B(net210669), .Y(n45408) );
  XOR2X1 U33209 ( .A(n34360), .B(n42592), .Y(n45137) );
  XNOR2X1 U33210 ( .A(n50518), .B(n41287), .Y(n24785) );
  XNOR2X1 U33211 ( .A(n50316), .B(n42707), .Y(n24934) );
  OAI21X2 U33212 ( .A0(n12078), .A1(net209956), .B0(n12145), .Y(n48124) );
  OAI211X2 U33213 ( .A0(n12076), .A1(n12077), .B0(n12078), .C0(n12079), .Y(
        n12075) );
  XNOR2X1 U33214 ( .A(n51162), .B(n41281), .Y(n24931) );
  XOR2X1 U33215 ( .A(n42059), .B(n41319), .Y(n45011) );
  CLKBUFX2 U33216 ( .A(n42692), .Y(n42691) );
  OR4X4 U33217 ( .A(n44953), .B(n44952), .C(n44951), .D(n44950), .Y(n41706) );
  XOR2X1 U33218 ( .A(n34372), .B(n42637), .Y(n44950) );
  XNOR2X1 U33219 ( .A(n34370), .B(n42560), .Y(n44930) );
  XOR2X1 U33220 ( .A(n34425), .B(n41379), .Y(n45271) );
  XNOR2X1 U33221 ( .A(n51185), .B(n42632), .Y(n26726) );
  XNOR2X1 U33222 ( .A(n50732), .B(n36865), .Y(n24954) );
  XNOR2X1 U33223 ( .A(n50543), .B(n41319), .Y(n26730) );
  XOR2X1 U33224 ( .A(n34428), .B(n42638), .Y(n45257) );
  AND2XL U33225 ( .A(n12151), .B(n12152), .Y(n12042) );
  OAI21X2 U33226 ( .A0(n12152), .A1(net209971), .B0(n10544), .Y(n48116) );
  XOR2X1 U33227 ( .A(n34405), .B(n42631), .Y(n45066) );
  XOR2X1 U33228 ( .A(n41908), .B(n42605), .Y(n24775) );
  XNOR2X1 U33229 ( .A(n51216), .B(n41283), .Y(n27577) );
  XNOR2X1 U33230 ( .A(n51416), .B(n36861), .Y(n29228) );
  XOR2X1 U33231 ( .A(n41820), .B(n42610), .Y(n45379) );
  XOR2X1 U33232 ( .A(n34356), .B(n42638), .Y(n45141) );
  XOR2X1 U33233 ( .A(n34304), .B(net219468), .Y(n45386) );
  CLKINVX4 U33234 ( .A(n41289), .Y(n41297) );
  XNOR2X1 U33235 ( .A(n50787), .B(n42592), .Y(n27570) );
  XOR2X1 U33236 ( .A(n34345), .B(n42576), .Y(n45161) );
  XOR2X1 U33237 ( .A(n34406), .B(n42533), .Y(n44998) );
  XOR2X1 U33238 ( .A(n34368), .B(net219434), .Y(n45145) );
  AOI211X2 U33239 ( .A0(n11431), .A1(n11432), .B0(net151720), .C0(net151721),
        .Y(n11429) );
  XNOR2X1 U33240 ( .A(n50946), .B(n42613), .Y(n24952) );
  XNOR2X1 U33241 ( .A(n50314), .B(n42672), .Y(n24956) );
  NOR2X4 U33242 ( .A(n10843), .B(n47174), .Y(n47178) );
  XOR2X1 U33243 ( .A(n34354), .B(n42669), .Y(n45143) );
  XNOR2X1 U33244 ( .A(n51358), .B(n42698), .Y(n28304) );
  XOR2X1 U33245 ( .A(n34362), .B(n42707), .Y(n45151) );
  NAND4X4 U33246 ( .A(n43634), .B(n43633), .C(n43632), .D(n43631), .Y(n12794)
         );
  OAI21X4 U33247 ( .A0(n48193), .A1(n48192), .B0(n48191), .Y(n48199) );
  OAI21X1 U33248 ( .A0(n48184), .A1(n48183), .B0(n48182), .Y(n48192) );
  XNOR2X1 U33249 ( .A(n50518), .B(n36905), .Y(n24957) );
  XOR2X1 U33250 ( .A(n34292), .B(n42638), .Y(n45382) );
  XNOR2X1 U33251 ( .A(n50370), .B(n42711), .Y(n27580) );
  XOR2X1 U33252 ( .A(n34293), .B(n42633), .Y(n45381) );
  XNOR2X1 U33253 ( .A(n51213), .B(n41282), .Y(n27547) );
  XOR2X1 U33254 ( .A(n42068), .B(n42659), .Y(n44915) );
  NOR4X2 U33255 ( .A(n24934), .B(n24935), .C(n24936), .D(n24937), .Y(n44508)
         );
  XNOR2X1 U33256 ( .A(n50520), .B(n36709), .Y(n24935) );
  NOR4X4 U33257 ( .A(n29023), .B(n29024), .C(n29025), .D(n29026), .Y(n43671)
         );
  XNOR2X1 U33258 ( .A(n51402), .B(n42701), .Y(n29025) );
  XOR2X1 U33259 ( .A(n34408), .B(n34450), .Y(n45063) );
  XOR2X1 U33260 ( .A(n34356), .B(n42690), .Y(n45120) );
  XOR2X1 U33261 ( .A(n34352), .B(net219468), .Y(n45205) );
  XOR2X1 U33262 ( .A(n34340), .B(n42638), .Y(n45201) );
  XNOR2X1 U33263 ( .A(n34374), .B(n42538), .Y(n44935) );
  XOR2X1 U33264 ( .A(n34426), .B(n42669), .Y(n45269) );
  NOR4X1 U33265 ( .A(n26758), .B(n26756), .C(n26755), .D(n26757), .Y(n44602)
         );
  XNOR2X1 U33266 ( .A(n50972), .B(n42615), .Y(n26755) );
  XOR2X1 U33267 ( .A(n42098), .B(n42658), .Y(n44015) );
  XOR2X1 U33268 ( .A(n34428), .B(n41385), .Y(n45030) );
  XOR2X1 U33269 ( .A(n34360), .B(net219468), .Y(n45116) );
  XOR2X1 U33270 ( .A(n34352), .B(n42592), .Y(n45108) );
  XOR2X1 U33271 ( .A(n41838), .B(n42604), .Y(n43980) );
  XOR2X1 U33272 ( .A(n34300), .B(n42644), .Y(n45496) );
  XNOR2X1 U33273 ( .A(n34373), .B(n42548), .Y(n44934) );
  XOR2X1 U33274 ( .A(n34368), .B(n34450), .Y(n44965) );
  XNOR2X1 U33275 ( .A(n34390), .B(n42537), .Y(n45103) );
  XOR2X1 U33276 ( .A(n34344), .B(n34450), .Y(n45197) );
  XOR2X1 U33277 ( .A(n34372), .B(n41385), .Y(n44977) );
  XOR2X1 U33278 ( .A(n36854), .B(n34408), .Y(n46562) );
  XNOR2X1 U33279 ( .A(n50714), .B(n36857), .Y(n23185) );
  XNOR2X1 U33280 ( .A(n50717), .B(n36852), .Y(n23135) );
  XOR2X1 U33281 ( .A(n34148), .B(n42637), .Y(n43983) );
  CLKINVX6 U33282 ( .A(n41326), .Y(n41333) );
  XOR2X1 U33283 ( .A(n42097), .B(n42658), .Y(n43984) );
  XOR2X1 U33284 ( .A(n34373), .B(n41282), .Y(n44976) );
  XOR2X1 U33285 ( .A(n34401), .B(n42681), .Y(n45070) );
  NOR4X2 U33286 ( .A(n43986), .B(n43985), .C(n43984), .D(n43983), .Y(n43997)
         );
  BUFX12 U33287 ( .A(n51442), .Y(codeword[7]) );
  INVX12 U33288 ( .A(n41796), .Y(busy) );
  NAND2X1 U33289 ( .A(n9679), .B(n41796), .Y(n19382) );
  NAND3BX1 U33290 ( .AN(n19411), .B(n41796), .C(n19336), .Y(n19374) );
  NOR2X4 U33291 ( .A(state[0]), .B(state[1]), .Y(n41796) );
  INVX3 U33292 ( .A(n37182), .Y(n50140) );
  CLKAND2X12 U33293 ( .A(n9679), .B(drop_done), .Y(finish) );
  BUFX12 U33294 ( .A(n51441), .Y(codeword[8]) );
  INVX12 U33295 ( .A(n40772), .Y(codeword[2]) );
  BUFX12 U33296 ( .A(n51440), .Y(codeword[9]) );
  BUFX12 U33297 ( .A(n51446), .Y(codeword[1]) );
  BUFX12 U33298 ( .A(n51447), .Y(codeword[0]) );
  BUFX12 U33299 ( .A(n51439), .Y(codeword[10]) );
  BUFX12 U33300 ( .A(n51443), .Y(codeword[6]) );
  INVX12 U33301 ( .A(n40038), .Y(codeword[4]) );
  NOR2X4 U33302 ( .A(n50149), .B(state[0]), .Y(n41736) );
  OR2X6 U33303 ( .A(net209509), .B(n48372), .Y(n41343) );
  NAND2X6 U33304 ( .A(n41343), .B(net207653), .Y(n48373) );
  AOI21X2 U33305 ( .A0(n48373), .A1(net207642), .B0(net171305), .Y(n48375) );
  NAND2XL U33306 ( .A(n34422), .B(net258261), .Y(n41346) );
  NOR2X4 U33307 ( .A(n43837), .B(n48337), .Y(n43841) );
  XNOR2XL U33308 ( .A(n34098), .B(n42569), .Y(n43840) );
  AO21X2 U33309 ( .A0(n48135), .A1(n48187), .B0(n48134), .Y(n41778) );
  NAND2XL U33310 ( .A(n41349), .B(n36731), .Y(n41351) );
  NOR4X2 U33311 ( .A(n44943), .B(n44942), .C(n44941), .D(n44940), .Y(n44964)
         );
  AOI21X4 U33312 ( .A0(n48517), .A1(n12388), .B0(net209210), .Y(n48518) );
  OR2X6 U33313 ( .A(n39520), .B(n48529), .Y(n41353) );
  NAND2X6 U33314 ( .A(n41353), .B(n11050), .Y(n48531) );
  AOI21X4 U33315 ( .A0(n48528), .A1(n48527), .B0(net171462), .Y(n48529) );
  AOI21X4 U33316 ( .A0(n48531), .A1(n12270), .B0(n48530), .Y(n48533) );
  NAND2XL U33317 ( .A(n51370), .B(n42696), .Y(n41354) );
  NAND2X1 U33318 ( .A(n33572), .B(n36923), .Y(n41355) );
  NAND2X1 U33319 ( .A(n41354), .B(n41355), .Y(n24816) );
  OA21X4 U33320 ( .A0(n11112), .A1(n11113), .B0(n11114), .Y(n41356) );
  AO21X4 U33321 ( .A0(n11108), .A1(n11109), .B0(net171423), .Y(n41635) );
  NAND2XL U33322 ( .A(net209620), .B(n46482), .Y(net258199) );
  AOI2BB1X4 U33323 ( .A0N(n47759), .A1N(n41751), .B0(n47771), .Y(n47775) );
  NAND2X1 U33324 ( .A(n9670), .B(n36923), .Y(n41359) );
  NAND2XL U33325 ( .A(n41358), .B(n42693), .Y(n41360) );
  NAND2X1 U33326 ( .A(n41359), .B(n41360), .Y(n45248) );
  OR2X8 U33327 ( .A(net209479), .B(n48393), .Y(n41361) );
  NAND2X6 U33328 ( .A(n41361), .B(n10089), .Y(n48395) );
  AOI21X4 U33329 ( .A0(n48392), .A1(n11673), .B0(net209482), .Y(n48393) );
  AOI21X4 U33330 ( .A0(n48395), .A1(n10090), .B0(n48394), .Y(n48396) );
  OR2X8 U33331 ( .A(net209466), .B(n48402), .Y(n41362) );
  NAND2X6 U33332 ( .A(n41362), .B(n11649), .Y(n48403) );
  CLKINVX2 U33333 ( .A(n11652), .Y(net209466) );
  AOI21X4 U33334 ( .A0(n48401), .A1(n11658), .B0(net209469), .Y(n48402) );
  AOI21X4 U33335 ( .A0(n48403), .A1(n11650), .B0(net171143), .Y(n48404) );
  OR2X2 U33336 ( .A(n41363), .B(n41364), .Y(n47729) );
  OR2X8 U33337 ( .A(n47749), .B(net210635), .Y(n41365) );
  OR3X4 U33338 ( .A(n11753), .B(net171185), .C(net171192), .Y(n41366) );
  AOI211X2 U33339 ( .A0(n11757), .A1(n11758), .B0(net151308), .C0(net209661),
        .Y(n11753) );
  NAND2XL U33340 ( .A(n41367), .B(n41647), .Y(n41370) );
  INVXL U33341 ( .A(n42615), .Y(n41368) );
  AOI21X4 U33342 ( .A0(n48550), .A1(n40391), .B0(net151503), .Y(n48551) );
  NOR2X6 U33343 ( .A(n12087), .B(n45690), .Y(net213362) );
  NAND4BBX4 U33344 ( .AN(n46478), .BN(n41722), .C(n46477), .D(net210479), .Y(
        n48439) );
  AOI211X2 U33345 ( .A0(n11086), .A1(n11087), .B0(net171441), .C0(net171440),
        .Y(n11080) );
  OAI21X4 U33346 ( .A0(net171099), .A1(n48407), .B0(n12459), .Y(n48408) );
  AOI21X4 U33347 ( .A0(n48406), .A1(n11638), .B0(net171104), .Y(n48407) );
  AO21X4 U33348 ( .A0(n12074), .A1(n12075), .B0(net171191), .Y(n41375) );
  OAI211X2 U33349 ( .A0(n12070), .A1(n12071), .B0(n12072), .C0(n12073), .Y(
        n12067) );
  OAI211X2 U33350 ( .A0(n12022), .A1(n12023), .B0(n10529), .C0(n12024), .Y(
        n12019) );
  AOI211X2 U33351 ( .A0(n12027), .A1(n12028), .B0(net171199), .C0(net171218),
        .Y(n12022) );
  NAND2XL U33352 ( .A(n37202), .B(n42660), .Y(n41378) );
  INVXL U33353 ( .A(n42660), .Y(n41376) );
  BUFX20 U33354 ( .A(n42666), .Y(n42660) );
  NAND2X1 U33355 ( .A(n42130), .B(n36917), .Y(n41382) );
  NAND2XL U33356 ( .A(n37250), .B(n42653), .Y(n41383) );
  NAND2X1 U33357 ( .A(n41382), .B(n41383), .Y(n29289) );
  AOI211X2 U33358 ( .A0(n11361), .A1(n11362), .B0(n50102), .C0(n50103), .Y(
        n11356) );
  XOR2X1 U33359 ( .A(n34380), .B(n42637), .Y(n44914) );
  OA21X4 U33360 ( .A0(n11136), .A1(n11137), .B0(n11138), .Y(n41386) );
  AOI211X2 U33361 ( .A0(n11141), .A1(n11142), .B0(net171427), .C0(net171425),
        .Y(n11136) );
  AOI211X2 U33362 ( .A0(n11134), .A1(n11133), .B0(net171433), .C0(n39953), .Y(
        n11128) );
  NAND2XL U33363 ( .A(n41387), .B(n42638), .Y(n41390) );
  OAI211X2 U33364 ( .A0(n11106), .A1(n11107), .B0(n10852), .C0(n10855), .Y(
        n11103) );
  CLKBUFX2 U33365 ( .A(n42474), .Y(n42473) );
  CLKBUFX2 U33366 ( .A(n42476), .Y(n42469) );
  CLKBUFX2 U33367 ( .A(n42468), .Y(n42460) );
  CLKBUFX2 U33368 ( .A(n42468), .Y(n42467) );
  CLKBUFX2 U33369 ( .A(n42492), .Y(n42491) );
  CLKBUFX2 U33370 ( .A(n42492), .Y(n42489) );
  CLKBUFX2 U33371 ( .A(n42478), .Y(n42484) );
  INVX3 U33372 ( .A(net256309), .Y(net209924) );
  NAND2XL U33373 ( .A(net209620), .B(n46482), .Y(n48147) );
  OAI21X2 U33374 ( .A0(n12040), .A1(n10542), .B0(n12041), .Y(n12037) );
  OAI211X2 U33375 ( .A0(n12030), .A1(n12031), .B0(n12032), .C0(n12033), .Y(
        n12028) );
  OAI2BB1X4 U33376 ( .A0N(n40405), .A1N(n41699), .B0(n10672), .Y(n48110) );
  AO21X4 U33377 ( .A0(n48109), .A1(n11314), .B0(net171534), .Y(n41699) );
  NAND2XL U33378 ( .A(n48439), .B(n48441), .Y(net210582) );
  NOR2X1 U33379 ( .A(n10872), .B(n47026), .Y(n47030) );
  NOR2X1 U33380 ( .A(n11057), .B(n46709), .Y(n46713) );
  NOR2X2 U33381 ( .A(n12323), .B(n47233), .Y(n47237) );
  NAND2XL U33382 ( .A(n41911), .B(n36915), .Y(n41631) );
  NAND2XL U33383 ( .A(n37203), .B(n36898), .Y(n41632) );
  NAND2X1 U33384 ( .A(n41631), .B(n41632), .Y(n28151) );
  NOR4X4 U33385 ( .A(n28148), .B(n28149), .C(n28150), .D(n28151), .Y(n43797)
         );
  AOI211X2 U33386 ( .A0(n11102), .A1(n11103), .B0(net171418), .C0(net171417),
        .Y(n11100) );
  NAND4BBX4 U33387 ( .AN(n46586), .BN(n46585), .C(net212238), .D(n46584), .Y(
        net209335) );
  NAND4BX4 U33388 ( .AN(n46575), .B(n41665), .C(n46574), .D(net209622), .Y(
        n48436) );
  XOR2XL U33389 ( .A(n42062), .B(n42557), .Y(n45050) );
  AOI21X1 U33390 ( .A0(n10529), .A1(net171214), .B0(net171205), .Y(n48241) );
  NOR2X4 U33391 ( .A(n44722), .B(n48320), .Y(n44732) );
  INVX1 U33392 ( .A(n10526), .Y(net171132) );
  INVX3 U33393 ( .A(net211271), .Y(net171421) );
  CLKINVX4 U33394 ( .A(net209242), .Y(net171423) );
  XOR2XL U33395 ( .A(n34418), .B(n41630), .Y(n45284) );
  NAND4X1 U33396 ( .A(n43413), .B(n43412), .C(n43411), .D(n43410), .Y(n10493)
         );
  AOI21X4 U33397 ( .A0(n48270), .A1(net260251), .B0(net209739), .Y(n48271) );
  INVXL U33398 ( .A(n10544), .Y(net171307) );
  AO21X2 U33399 ( .A0(n48126), .A1(n10559), .B0(net209953), .Y(n41704) );
  XOR2X1 U33400 ( .A(n42124), .B(n36882), .Y(n29177) );
  XNOR2XL U33401 ( .A(n50921), .B(n42617), .Y(n31359) );
  XNOR2XL U33402 ( .A(n50289), .B(n36907), .Y(n31363) );
  XNOR2XL U33403 ( .A(n50707), .B(n42588), .Y(n31361) );
  XNOR2XL U33404 ( .A(n51135), .B(n42633), .Y(n31360) );
  NOR2X2 U33405 ( .A(n12539), .B(n43582), .Y(n43586) );
  NOR2XL U33406 ( .A(n10544), .B(n45748), .Y(n45752) );
  NOR2X1 U33407 ( .A(n12488), .B(n43267), .Y(n43271) );
  CLKBUFX3 U33408 ( .A(n33143), .Y(n41964) );
  CLKBUFX3 U33409 ( .A(n33139), .Y(n42223) );
  NAND2XL U33410 ( .A(n41348), .B(n42612), .Y(n41640) );
  INVX2 U33411 ( .A(n42571), .Y(n42563) );
  NOR4X1 U33412 ( .A(n28272), .B(n28273), .C(n28274), .D(n28275), .Y(n43760)
         );
  AOI211X2 U33413 ( .A0(n12036), .A1(n12037), .B0(net171313), .C0(n39561), .Y(
        n12030) );
  XOR2XL U33414 ( .A(n41803), .B(n36868), .Y(n45016) );
  NOR2X1 U33415 ( .A(n46583), .B(n46582), .Y(n46584) );
  OAI21X4 U33416 ( .A0(net209145), .A1(n48551), .B0(n10992), .Y(n48552) );
  OAI211X2 U33417 ( .A0(n39987), .A1(n11000), .B0(n40400), .C0(n11002), .Y(
        n10998) );
  OAI31X2 U33418 ( .A0(n11003), .A1(net171474), .A2(net171476), .B0(n10273),
        .Y(n11000) );
  NAND3X1 U33419 ( .A(n11389), .B(n10752), .C(n10753), .Y(n48065) );
  CLKINVX1 U33420 ( .A(n11417), .Y(net210239) );
  XOR2X1 U33421 ( .A(n42214), .B(n42652), .Y(n31065) );
  XOR2X1 U33422 ( .A(n41955), .B(n42607), .Y(n31061) );
  NOR2XL U33423 ( .A(n47263), .B(net211197), .Y(n47267) );
  NOR2XL U33424 ( .A(n10553), .B(n45618), .Y(n45622) );
  NOR2X2 U33425 ( .A(n11732), .B(n44247), .Y(n44251) );
  NOR2X1 U33426 ( .A(n12329), .B(n47253), .Y(n47257) );
  NOR2X1 U33427 ( .A(n12278), .B(n46769), .Y(n46773) );
  AO21X4 U33428 ( .A0(n48282), .A1(n11756), .B0(net209659), .Y(n41741) );
  AOI31XL U33429 ( .A0(n48313), .A1(n48312), .A2(n48311), .B0(n48310), .Y(
        n48317) );
  NAND4X4 U33430 ( .A(n44312), .B(n44311), .C(n44310), .D(n44309), .Y(n11741)
         );
  NOR3X1 U33431 ( .A(n44496), .B(n44495), .C(n44494), .Y(n44498) );
  XNOR2X1 U33432 ( .A(n50952), .B(n42539), .Y(n24972) );
  XNOR2XL U33433 ( .A(n49515), .B(net219310), .Y(n27727) );
  OA21X2 U33434 ( .A0(n36948), .A1(n48056), .B0(n12962), .Y(n41701) );
  OA21X2 U33435 ( .A0(net171532), .A1(n48098), .B0(n12909), .Y(n41703) );
  OAI2BB1X2 U33436 ( .A0N(n12715), .A1N(n41779), .B0(n40392), .Y(n48232) );
  XOR2X1 U33437 ( .A(n42554), .B(n41802), .Y(n44031) );
  NOR2X1 U33438 ( .A(n44753), .B(n48326), .Y(n44763) );
  OAI21X1 U33439 ( .A0(net151737), .A1(n48075), .B0(n10751), .Y(n48076) );
  INVXL U33440 ( .A(n12967), .Y(net151721) );
  XOR2XL U33441 ( .A(n41316), .B(n41807), .Y(n46561) );
  INVX3 U33442 ( .A(n11366), .Y(n47957) );
  AOI211X2 U33443 ( .A0(n47969), .A1(n11414), .B0(n47968), .C0(n36944), .Y(
        n48072) );
  OAI21X1 U33444 ( .A0(net210239), .A1(n47966), .B0(n11415), .Y(n47969) );
  CLKINVX3 U33445 ( .A(n12342), .Y(net151712) );
  CLKINVX3 U33446 ( .A(n13014), .Y(net151672) );
  AO21X4 U33447 ( .A0(n48073), .A1(n12940), .B0(net171551), .Y(n41694) );
  OAI2BB1X4 U33448 ( .A0N(n11399), .A1N(n41694), .B0(n11397), .Y(n48074) );
  AOI21X4 U33449 ( .A0(n48093), .A1(n12915), .B0(n36942), .Y(n48094) );
  OAI21X1 U33450 ( .A0(n39631), .A1(n48094), .B0(n11350), .Y(n48095) );
  XNOR2XL U33451 ( .A(n51349), .B(n42702), .Y(n31373) );
  XOR2XL U33452 ( .A(n41932), .B(n42605), .Y(n31362) );
  XNOR2XL U33453 ( .A(n50294), .B(n42711), .Y(n31581) );
  XNOR2XL U33454 ( .A(n50925), .B(n42617), .Y(n31569) );
  XNOR2XL U33455 ( .A(n50293), .B(n42670), .Y(n31573) );
  XNOR2XL U33456 ( .A(n50498), .B(n42717), .Y(n31582) );
  XNOR2XL U33457 ( .A(n51139), .B(n34447), .Y(n31570) );
  XNOR2XL U33458 ( .A(n50497), .B(n41380), .Y(n31574) );
  XNOR2XL U33459 ( .A(n50494), .B(n36728), .Y(n31364) );
  XOR2XL U33460 ( .A(n41931), .B(n36897), .Y(n31370) );
  XOR2XL U33461 ( .A(n42190), .B(n36885), .Y(n31374) );
  NOR4X2 U33462 ( .A(n31307), .B(n31308), .C(n31309), .D(n31310), .Y(n43291)
         );
  INVX1 U33463 ( .A(n12904), .Y(net210067) );
  XOR2XL U33464 ( .A(n34238), .B(n36868), .Y(n44828) );
  NOR2X2 U33465 ( .A(n40396), .B(n47154), .Y(n47158) );
  NOR2X2 U33466 ( .A(n12486), .B(n43294), .Y(n43298) );
  AOI211X2 U33467 ( .A0(n11745), .A1(n11746), .B0(n49503), .C0(n49507), .Y(
        n11739) );
  NAND2XL U33468 ( .A(n41643), .B(n42627), .Y(n41645) );
  CLKINVX2 U33469 ( .A(n42572), .Y(n42561) );
  OAI2BB1X1 U33470 ( .A0N(n11751), .A1N(n41741), .B0(n11752), .Y(n48284) );
  AOI21X1 U33471 ( .A0(n41757), .A1(n48332), .B0(n39479), .Y(n48333) );
  NOR4X1 U33472 ( .A(n27034), .B(n27035), .C(n27036), .D(n27037), .Y(n44244)
         );
  NAND4X4 U33473 ( .A(n43799), .B(n43798), .C(n43797), .D(n43796), .Y(n12586)
         );
  NOR4X2 U33474 ( .A(n28140), .B(n28141), .C(n28142), .D(n28143), .Y(n43799)
         );
  NOR4X2 U33475 ( .A(n26853), .B(n26854), .C(n26855), .D(n26856), .Y(n44310)
         );
  NAND2XL U33476 ( .A(n48320), .B(n48319), .Y(net210641) );
  INVXL U33477 ( .A(n47979), .Y(n47991) );
  NAND4X1 U33478 ( .A(n43058), .B(n43057), .C(n43056), .D(n43055), .Y(n12589)
         );
  NAND4X1 U33479 ( .A(n43081), .B(n43080), .C(n43079), .D(n43078), .Y(n12453)
         );
  XOR2X1 U33480 ( .A(n42100), .B(n41286), .Y(n43860) );
  XOR2X1 U33481 ( .A(n41841), .B(n42600), .Y(n43856) );
  XNOR2X1 U33482 ( .A(n51180), .B(n41282), .Y(n26915) );
  XOR2X1 U33483 ( .A(n41889), .B(n42607), .Y(n26939) );
  XOR2X1 U33484 ( .A(n42148), .B(n42663), .Y(n26943) );
  XNOR2X1 U33485 ( .A(n50768), .B(net219450), .Y(n29412) );
  XNOR2XL U33486 ( .A(n51394), .B(n42696), .Y(n26679) );
  NOR4X2 U33487 ( .A(n45444), .B(n45443), .C(n45442), .D(n45441), .Y(n45453)
         );
  XOR2XL U33488 ( .A(n42076), .B(n36801), .Y(n45412) );
  XNOR2XL U33489 ( .A(n51422), .B(n42697), .Y(n27191) );
  OAI211X2 U33490 ( .A0(n11405), .A1(n11404), .B0(n10706), .C0(n10708), .Y(
        n11401) );
  INVXL U33491 ( .A(n11411), .Y(net151753) );
  XOR2XL U33492 ( .A(n36811), .B(n42065), .Y(n46558) );
  XNOR2XL U33493 ( .A(n50765), .B(net219450), .Y(n29442) );
  NOR4X1 U33494 ( .A(n29440), .B(n29441), .C(n29442), .D(n29443), .Y(n43556)
         );
  OAI2BB1X2 U33495 ( .A0N(n48188), .A1N(n41778), .B0(n10184), .Y(n48136) );
  XNOR2X1 U33496 ( .A(n51353), .B(n42701), .Y(n31583) );
  AOI21X1 U33497 ( .A0(n48017), .A1(n48016), .B0(n48015), .Y(n48026) );
  XNOR2X1 U33498 ( .A(n50926), .B(n40039), .Y(n31577) );
  XNOR2X1 U33499 ( .A(n51140), .B(n41281), .Y(n31578) );
  AOI21X1 U33500 ( .A0(n47994), .A1(n47993), .B0(n47992), .Y(n48004) );
  OAI21XL U33501 ( .A0(n47991), .A1(n47990), .B0(n47989), .Y(n47992) );
  XOR2XL U33502 ( .A(n36811), .B(n42077), .Y(n46313) );
  INVX1 U33503 ( .A(n10608), .Y(net209821) );
  INVX1 U33504 ( .A(n12072), .Y(net209953) );
  OAI21X1 U33505 ( .A0(n39560), .A1(n48243), .B0(n12014), .Y(n48244) );
  AOI21XL U33506 ( .A0(n48001), .A1(n48000), .B0(n47999), .Y(n48002) );
  INVXL U33507 ( .A(n47996), .Y(n48001) );
  NAND4BBXL U33508 ( .AN(n48024), .BN(n48023), .C(n48034), .D(n48022), .Y(
        n48025) );
  NAND2XL U33509 ( .A(n48027), .B(n48038), .Y(n48024) );
  NAND2XL U33510 ( .A(n48021), .B(n48020), .Y(n48022) );
  XOR2XL U33511 ( .A(n42544), .B(n41805), .Y(n44030) );
  OAI2BB1X4 U33512 ( .A0N(n41700), .A1N(n41701), .B0(n48061), .Y(n48071) );
  OAI2BB1XL U33513 ( .A0N(n48027), .A1N(n41785), .B0(n48036), .Y(n48039) );
  AO21XL U33514 ( .A0(n48035), .A1(n48034), .B0(n48033), .Y(n41785) );
  INVX3 U33515 ( .A(n12004), .Y(net171125) );
  XOR2XL U33516 ( .A(n41928), .B(n41318), .Y(n23176) );
  INVXL U33517 ( .A(n47975), .Y(n47976) );
  INVX1 U33518 ( .A(n12252), .Y(net171472) );
  INVX1 U33519 ( .A(n11990), .Y(net209764) );
  INVX1 U33520 ( .A(n12246), .Y(net171470) );
  INVX1 U33521 ( .A(n10505), .Y(net171105) );
  XOR2XL U33522 ( .A(n36785), .B(n34393), .Y(n46594) );
  XOR2XL U33523 ( .A(n41331), .B(n34405), .Y(n46559) );
  XOR2XL U33524 ( .A(n9664), .B(n36897), .Y(n45245) );
  XNOR2XL U33525 ( .A(n41296), .B(n34382), .Y(n41795) );
  XNOR2XL U33526 ( .A(n36913), .B(n34381), .Y(n41794) );
  XOR2XL U33527 ( .A(n41303), .B(n34404), .Y(n46557) );
  XOR2XL U33528 ( .A(n36783), .B(n34401), .Y(n46556) );
  XOR2XL U33529 ( .A(n41295), .B(n34406), .Y(n46560) );
  NOR2X1 U33530 ( .A(n20127), .B(n20126), .Y(net211490) );
  NOR2X1 U33531 ( .A(n21092), .B(n21091), .Y(n46922) );
  XOR2XL U33532 ( .A(n36772), .B(n34401), .Y(n47681) );
  XOR2XL U33533 ( .A(n42470), .B(n34408), .Y(n47675) );
  NOR2X2 U33534 ( .A(n10573), .B(n45691), .Y(net213357) );
  NOR2XL U33535 ( .A(n12794), .B(n46108), .Y(n46112) );
  NOR2XL U33536 ( .A(n11139), .B(n47022), .Y(net211523) );
  NOR2X1 U33537 ( .A(n10566), .B(n46088), .Y(n46092) );
  XOR2XL U33538 ( .A(n41299), .B(n33452), .Y(n45853) );
  NOR2X1 U33539 ( .A(n12017), .B(n45910), .Y(n45914) );
  NOR2XL U33540 ( .A(n12793), .B(n45705), .Y(n45709) );
  NOR2XL U33541 ( .A(n12146), .B(n46153), .Y(n46157) );
  NOR2XL U33542 ( .A(n10606), .B(n45628), .Y(n45632) );
  NOR2XL U33543 ( .A(n10559), .B(n46133), .Y(n46137) );
  XOR2XL U33544 ( .A(n36798), .B(n34406), .Y(n47677) );
  XOR2XL U33545 ( .A(n36749), .B(n34404), .Y(n47678) );
  NOR2XL U33546 ( .A(n12005), .B(n45940), .Y(n45944) );
  NOR2XL U33547 ( .A(n11066), .B(n47068), .Y(n47072) );
  NOR2XL U33548 ( .A(n46966), .B(net211656), .Y(net211651) );
  NOR2XL U33549 ( .A(n40398), .B(n46935), .Y(n46939) );
  NOR2XL U33550 ( .A(n12150), .B(n46170), .Y(net212731) );
  NOR2XL U33551 ( .A(n11072), .B(n47108), .Y(n47112) );
  NOR2XL U33552 ( .A(n11074), .B(n47093), .Y(n47097) );
  NOR2XL U33553 ( .A(n12306), .B(n46972), .Y(net211641) );
  NOR2XL U33554 ( .A(n12318), .B(n47194), .Y(n47198) );
  NOR2XL U33555 ( .A(n12015), .B(n45920), .Y(n45924) );
  NOR2XL U33556 ( .A(n12156), .B(n46764), .Y(n46768) );
  NOR2XL U33557 ( .A(n12333), .B(n47897), .Y(n47901) );
  NOR2XL U33558 ( .A(n11201), .B(n47243), .Y(n47247) );
  NOR2XL U33559 ( .A(n45953), .B(net213021), .Y(net213016) );
  NOR2XL U33560 ( .A(n11035), .B(n46675), .Y(n46679) );
  AND4X1 U33561 ( .A(n46828), .B(n46827), .C(n46826), .D(n46825), .Y(net238868) );
  CLKINVX2 U33562 ( .A(n42572), .Y(n42562) );
  AOI21X1 U33563 ( .A0(n48277), .A1(n11699), .B0(net209669), .Y(n48278) );
  NOR2XL U33564 ( .A(net171237), .B(net171238), .Y(n11764) );
  NAND4X4 U33565 ( .A(n44201), .B(n44200), .C(n44199), .D(n44198), .Y(n11770)
         );
  NOR4X1 U33566 ( .A(n28091), .B(n28092), .C(n28093), .D(n28094), .Y(n43814)
         );
  NOR4X2 U33567 ( .A(n27185), .B(n27186), .C(n27187), .D(n27188), .Y(net215395) );
  OAI21XL U33568 ( .A0(n48331), .A1(n48330), .B0(n48329), .Y(n48332) );
  NOR3X1 U33569 ( .A(n45677), .B(n45676), .C(n45675), .Y(n45679) );
  XNOR2XL U33570 ( .A(n51002), .B(n42542), .Y(n27438) );
  NOR4X2 U33571 ( .A(n27189), .B(n27190), .C(n27191), .D(n27192), .Y(net215396) );
  AOI211X2 U33572 ( .A0(n11096), .A1(n11097), .B0(net171445), .C0(net171443),
        .Y(n11090) );
  INVXL U33573 ( .A(n10504), .Y(net209753) );
  XNOR2XL U33574 ( .A(n49512), .B(n42724), .Y(n27732) );
  NAND2XL U33575 ( .A(n10710), .B(n10709), .Y(n11405) );
  XOR2XL U33576 ( .A(n42158), .B(n36889), .Y(n24997) );
  XOR2XL U33577 ( .A(n41843), .B(n36899), .Y(n28000) );
  XNOR2XL U33578 ( .A(n50783), .B(net219444), .Y(n27247) );
  XNOR2XL U33579 ( .A(n42069), .B(n36873), .Y(n44933) );
  XOR2XL U33580 ( .A(n42106), .B(n36889), .Y(n27403) );
  XOR2XL U33581 ( .A(n41849), .B(n42608), .Y(n27421) );
  XOR2XL U33582 ( .A(n42108), .B(n42662), .Y(n27425) );
  XNOR2XL U33583 ( .A(n51005), .B(n40039), .Y(n27426) );
  XNOR2XL U33584 ( .A(n50791), .B(net219466), .Y(n27428) );
  XNOR2XL U33585 ( .A(n50992), .B(n42615), .Y(n27297) );
  XNOR2XL U33586 ( .A(n50993), .B(net219310), .Y(n27305) );
  XNOR2XL U33587 ( .A(n51004), .B(n42618), .Y(n27418) );
  XNOR2XL U33588 ( .A(n50997), .B(net219314), .Y(n27245) );
  XNOR2XL U33589 ( .A(n50790), .B(n42592), .Y(n27420) );
  XNOR2XL U33590 ( .A(n51431), .B(n42642), .Y(n27424) );
  XNOR2XL U33591 ( .A(n51219), .B(n41282), .Y(n27427) );
  XNOR2XL U33592 ( .A(n51218), .B(n42629), .Y(n27419) );
  XNOR2XL U33593 ( .A(n50372), .B(n42675), .Y(n27422) );
  XNOR2XL U33594 ( .A(n50778), .B(n36863), .Y(n27299) );
  XNOR2XL U33595 ( .A(n51419), .B(n42641), .Y(n27303) );
  XNOR2XL U33596 ( .A(n51206), .B(n42628), .Y(n27298) );
  XNOR2XL U33597 ( .A(n50564), .B(n36834), .Y(n27302) );
  XNOR2XL U33598 ( .A(n51211), .B(n41281), .Y(n27246) );
  XNOR2XL U33599 ( .A(n50576), .B(n36903), .Y(n27423) );
  OAI211X2 U33600 ( .A0(n11394), .A1(n11395), .B0(n11396), .C0(n11397), .Y(
        n11391) );
  XOR2XL U33601 ( .A(n41810), .B(n36899), .Y(n44955) );
  XOR2XL U33602 ( .A(n42072), .B(n41324), .Y(n45160) );
  INVXL U33603 ( .A(n11018), .Y(net209165) );
  OAI2BB1X4 U33604 ( .A0N(n11300), .A1N(n41698), .B0(n11301), .Y(n48114) );
  AO21X4 U33605 ( .A0(n48113), .A1(n12873), .B0(net151420), .Y(n41698) );
  OAI21X1 U33606 ( .A0(n48014), .A1(n48013), .B0(n48012), .Y(n48015) );
  XOR2XL U33607 ( .A(n42126), .B(n41322), .Y(n29156) );
  XOR2XL U33608 ( .A(n41842), .B(n42522), .Y(n43875) );
  OAI2BB1X4 U33609 ( .A0N(n11359), .A1N(net210081), .B0(n12918), .Y(n48093) );
  AOI211X2 U33610 ( .A0(n11124), .A1(n11125), .B0(net171483), .C0(net171482),
        .Y(n11122) );
  INVX1 U33611 ( .A(net210091), .Y(net171532) );
  INVXL U33612 ( .A(net209314), .Y(net209307) );
  XNOR2XL U33613 ( .A(n51397), .B(n42697), .Y(n26859) );
  XNOR2XL U33614 ( .A(n51196), .B(n41282), .Y(n29411) );
  XNOR2XL U33615 ( .A(n51187), .B(n41281), .Y(n26764) );
  XNOR2XL U33616 ( .A(n50544), .B(n41319), .Y(n26760) );
  XNOR2XL U33617 ( .A(n50545), .B(n42717), .Y(n26768) );
  XNOR2XL U33618 ( .A(n51400), .B(n42696), .Y(n26769) );
  XOR2XL U33619 ( .A(n41900), .B(n42522), .Y(n25095) );
  XNOR2XL U33620 ( .A(n50741), .B(net258207), .Y(n25112) );
  XOR2XL U33621 ( .A(n41869), .B(n36756), .Y(n19546) );
  XOR2XL U33622 ( .A(n42159), .B(n36883), .Y(n25027) );
  XOR2XL U33623 ( .A(n42113), .B(n36807), .Y(n23998) );
  XOR2XL U33624 ( .A(n41846), .B(n42525), .Y(n28012) );
  XOR2XL U33625 ( .A(n42131), .B(n36815), .Y(n22420) );
  XOR2XL U33626 ( .A(n41884), .B(n42522), .Y(n26688) );
  XOR2XL U33627 ( .A(n42107), .B(n42663), .Y(n27395) );
  XOR2XL U33628 ( .A(n41848), .B(n42609), .Y(n27391) );
  XOR2XL U33629 ( .A(n42109), .B(n42663), .Y(n27455) );
  XOR2XL U33630 ( .A(n42101), .B(n41322), .Y(n43878) );
  XOR2XL U33631 ( .A(n41870), .B(n41310), .Y(n22409) );
  XOR2XL U33632 ( .A(n41885), .B(n42607), .Y(n26878) );
  XOR2XL U33633 ( .A(n42144), .B(n42661), .Y(n26882) );
  XOR2XL U33634 ( .A(n41850), .B(n42609), .Y(n27451) );
  XOR2XL U33635 ( .A(n36887), .B(n42099), .Y(n43868) );
  XNOR2XL U33636 ( .A(n51409), .B(n36871), .Y(n29416) );
  XOR2XL U33637 ( .A(n42122), .B(n36886), .Y(n29237) );
  XOR2XL U33638 ( .A(n41863), .B(n36900), .Y(n29233) );
  XOR2XL U33639 ( .A(n42108), .B(n36889), .Y(n27463) );
  XOR2XL U33640 ( .A(n41854), .B(n42525), .Y(n27591) );
  XOR2XL U33641 ( .A(n41850), .B(n42525), .Y(n27411) );
  XNOR2XL U33642 ( .A(n50928), .B(n42620), .Y(n28440) );
  XNOR2XL U33643 ( .A(n50936), .B(n42620), .Y(n28500) );
  XNOR2XL U33644 ( .A(n50974), .B(n42620), .Y(n29011) );
  XNOR2XL U33645 ( .A(n50291), .B(n42711), .Y(n31611) );
  XNOR2XL U33646 ( .A(n51395), .B(n36867), .Y(n26881) );
  XNOR2XL U33647 ( .A(n50792), .B(net219466), .Y(n27398) );
  XNOR2XL U33648 ( .A(n51217), .B(n42554), .Y(n27409) );
  XNOR2XL U33649 ( .A(n51398), .B(n36867), .Y(n26731) );
  XNOR2XL U33650 ( .A(n51224), .B(n42551), .Y(n27710) );
  XNOR2XL U33651 ( .A(n50360), .B(n42674), .Y(n27301) );
  XNOR2XL U33652 ( .A(n50922), .B(n42617), .Y(n31599) );
  XNOR2XL U33653 ( .A(n50290), .B(n42670), .Y(n31603) );
  XNOR2XL U33654 ( .A(n50791), .B(n42592), .Y(n27390) );
  XNOR2XL U33655 ( .A(n51432), .B(n42642), .Y(n27394) );
  XNOR2XL U33656 ( .A(n51221), .B(n42626), .Y(n28080) );
  XNOR2XL U33657 ( .A(n51220), .B(n41282), .Y(n27397) );
  XNOR2XL U33658 ( .A(n51219), .B(n42633), .Y(n27389) );
  XNOR2XL U33659 ( .A(n50796), .B(n36737), .Y(n27711) );
  XNOR2XL U33660 ( .A(n50495), .B(n42722), .Y(n31612) );
  XNOR2XL U33661 ( .A(n51198), .B(n42554), .Y(n29303) );
  XNOR2XL U33662 ( .A(n51202), .B(n36832), .Y(n29213) );
  XNOR2XL U33663 ( .A(n51136), .B(n42631), .Y(n31600) );
  XNOR2XL U33664 ( .A(n37251), .B(n41380), .Y(n31604) );
  XOR2XL U33665 ( .A(n42129), .B(n36817), .Y(n22410) );
  XNOR2XL U33666 ( .A(n50756), .B(n42508), .Y(n26717) );
  XNOR2XL U33667 ( .A(n50708), .B(n42590), .Y(n31601) );
  XNOR2XL U33668 ( .A(n51209), .B(n36832), .Y(n27228) );
  XNOR2XL U33669 ( .A(n51349), .B(n42644), .Y(n31605) );
  XOR2XL U33670 ( .A(n42086), .B(n36877), .Y(n44787) );
  XNOR2XL U33671 ( .A(n50984), .B(n42535), .Y(n29302) );
  XNOR2XL U33672 ( .A(n50988), .B(n42535), .Y(n29212) );
  XNOR2XL U33673 ( .A(n50323), .B(n42707), .Y(n25114) );
  XNOR2XL U33674 ( .A(n50970), .B(n42540), .Y(n26715) );
  XNOR2XL U33675 ( .A(n50995), .B(n42541), .Y(n27227) );
  XNOR2XL U33676 ( .A(n50563), .B(n42581), .Y(n27292) );
  XNOR2XL U33677 ( .A(n50567), .B(n42581), .Y(n27232) );
  XNOR2XL U33678 ( .A(n50773), .B(n42501), .Y(n29184) );
  XNOR2XL U33679 ( .A(n50560), .B(n42577), .Y(n29217) );
  XNOR2XL U33680 ( .A(n50527), .B(n36709), .Y(n25115) );
  XNOR2XL U33681 ( .A(n50954), .B(n42613), .Y(n25102) );
  XNOR2XL U33682 ( .A(n50322), .B(n36907), .Y(n25106) );
  XNOR2XL U33683 ( .A(n50542), .B(n42576), .Y(n26720) );
  XNOR2XL U33684 ( .A(n50955), .B(net219310), .Y(n25110) );
  XNOR2XL U33685 ( .A(n50740), .B(n36865), .Y(n25104) );
  XOR2XL U33686 ( .A(n42109), .B(n41323), .Y(n27412) );
  XNOR2XL U33687 ( .A(n51168), .B(n42625), .Y(n25103) );
  XNOR2XL U33688 ( .A(n50526), .B(n36905), .Y(n25107) );
  XNOR2XL U33689 ( .A(n51169), .B(n41282), .Y(n25111) );
  XNOR2XL U33690 ( .A(n41890), .B(n36757), .Y(n41714) );
  XOR2XL U33691 ( .A(n41865), .B(n42529), .Y(n29215) );
  XOR2XL U33692 ( .A(n41837), .B(n36895), .Y(n43988) );
  XOR2XL U33693 ( .A(n36899), .B(n41840), .Y(n43864) );
  XNOR2XL U33694 ( .A(n50758), .B(net219434), .Y(n26735) );
  XOR2XL U33695 ( .A(n42124), .B(n36877), .Y(n29216) );
  INVXL U33696 ( .A(n10855), .Y(net209231) );
  XNOR2XL U33697 ( .A(n51219), .B(n42553), .Y(n28040) );
  NAND3XL U33698 ( .A(net209814), .B(n12715), .C(n12150), .Y(n48212) );
  NAND2XL U33699 ( .A(n11411), .B(n10709), .Y(n48063) );
  INVX4 U33700 ( .A(net211656), .Y(net171445) );
  AO21X4 U33701 ( .A0(n48520), .A1(net209202), .B0(net209203), .Y(n41780) );
  OAI2BB1X1 U33702 ( .A0N(n11065), .A1N(n41780), .B0(n48521), .Y(n48523) );
  XNOR2XL U33703 ( .A(n51121), .B(n41283), .Y(n31849) );
  XNOR2XL U33704 ( .A(n50693), .B(net219434), .Y(n31850) );
  XNOR2XL U33705 ( .A(n50907), .B(net219310), .Y(n31848) );
  XNOR2XL U33706 ( .A(n51117), .B(n41281), .Y(n31819) );
  XNOR2XL U33707 ( .A(n50689), .B(net219434), .Y(n31820) );
  XNOR2XL U33708 ( .A(n50903), .B(net219314), .Y(n31818) );
  XNOR2XL U33709 ( .A(n50481), .B(n36709), .Y(n31853) );
  XNOR2XL U33710 ( .A(n51134), .B(n42552), .Y(n31350) );
  XNOR2XL U33711 ( .A(n50706), .B(n42505), .Y(n31351) );
  XNOR2XL U33712 ( .A(n50920), .B(n42537), .Y(n31349) );
  XNOR2XL U33713 ( .A(n50494), .B(n42578), .Y(n31594) );
  XNOR2XL U33714 ( .A(n50493), .B(n42580), .Y(n31354) );
  XOR2XL U33715 ( .A(n42150), .B(n42489), .Y(n19790) );
  XOR2XL U33716 ( .A(n41843), .B(n41318), .Y(n23777) );
  XOR2XL U33717 ( .A(n41891), .B(n36759), .Y(n19789) );
  XOR2XL U33718 ( .A(n42102), .B(n36808), .Y(n23778) );
  INVXL U33719 ( .A(n12318), .Y(net151612) );
  XOR2XL U33720 ( .A(n41854), .B(n41314), .Y(n23997) );
  XOR2XL U33721 ( .A(n41962), .B(n36898), .Y(n32092) );
  XOR2XL U33722 ( .A(n42221), .B(n36886), .Y(n32096) );
  XNOR2XL U33723 ( .A(n51332), .B(n41302), .Y(n22806) );
  XOR2XL U33724 ( .A(n42222), .B(n42657), .Y(n32088) );
  XNOR2XL U33725 ( .A(n50275), .B(n41641), .Y(n31852) );
  XNOR2XL U33726 ( .A(n51333), .B(n42642), .Y(n31846) );
  XOR2XL U33727 ( .A(n41963), .B(n42605), .Y(n32084) );
  INVXL U33728 ( .A(n11969), .Y(net209750) );
  XOR2X1 U33729 ( .A(n34425), .B(n42723), .Y(n45040) );
  XOR2XL U33730 ( .A(n34388), .B(n42699), .Y(n44922) );
  XOR2XL U33731 ( .A(n34012), .B(n36827), .Y(n44193) );
  XNOR2XL U33732 ( .A(n34372), .B(n36831), .Y(n44931) );
  XOR2XL U33733 ( .A(n34262), .B(n36868), .Y(n44855) );
  NOR2X1 U33734 ( .A(n20137), .B(n20136), .Y(net211480) );
  XOR2XL U33735 ( .A(n34350), .B(n41647), .Y(n45110) );
  XOR2XL U33736 ( .A(n34345), .B(n41380), .Y(n45115) );
  XOR2XL U33737 ( .A(n34337), .B(n42576), .Y(n45130) );
  XOR2XL U33738 ( .A(n34348), .B(n42638), .Y(n45112) );
  XOR2XL U33739 ( .A(n34342), .B(n42534), .Y(n45127) );
  XOR2XL U33740 ( .A(n34341), .B(n36832), .Y(n45128) );
  NOR2X2 U33741 ( .A(n19538), .B(n19537), .Y(n47265) );
  NOR4X2 U33742 ( .A(n19536), .B(n19535), .C(n19534), .D(n19533), .Y(n47264)
         );
  XOR2XL U33743 ( .A(n41304), .B(n34380), .Y(n46484) );
  NOR2X2 U33744 ( .A(n11084), .B(n46920), .Y(n46924) );
  XOR2XL U33745 ( .A(n34401), .B(n42575), .Y(n45002) );
  NOR2XL U33746 ( .A(n10846), .B(n46955), .Y(n46959) );
  NOR4X2 U33747 ( .A(n20125), .B(n20124), .C(n20123), .D(n20122), .Y(net211491) );
  NOR2X2 U33748 ( .A(n11209), .B(n46930), .Y(n46934) );
  XOR2XL U33749 ( .A(n34105), .B(n36783), .Y(n46200) );
  XOR2XL U33750 ( .A(n33988), .B(n36829), .Y(n44207) );
  XOR2XL U33751 ( .A(n34394), .B(n42670), .Y(n45088) );
  XOR2XL U33752 ( .A(n34392), .B(n42592), .Y(n44880) );
  XOR2XL U33753 ( .A(n33337), .B(n36780), .Y(n45940) );
  XOR2XL U33754 ( .A(n34154), .B(n42705), .Y(n43993) );
  XOR2XL U33755 ( .A(n42096), .B(n36882), .Y(n43992) );
  NOR2X1 U33756 ( .A(n23198), .B(n23197), .Y(n45850) );
  NOR2X1 U33757 ( .A(n22958), .B(n22957), .Y(n45917) );
  XOR2XL U33758 ( .A(n34160), .B(net219466), .Y(n43987) );
  XOR2XL U33759 ( .A(n41332), .B(n34421), .Y(n46599) );
  XOR2XL U33760 ( .A(n34149), .B(n42625), .Y(n43982) );
  XOR2XL U33761 ( .A(n34145), .B(n41379), .Y(n43986) );
  XOR2XL U33762 ( .A(n34157), .B(n41282), .Y(n43990) );
  XOR2XL U33763 ( .A(n34309), .B(n42549), .Y(n45457) );
  XOR2XL U33764 ( .A(n34156), .B(n41385), .Y(n43991) );
  XOR2XL U33765 ( .A(n34158), .B(net219330), .Y(n43989) );
  XOR2XL U33766 ( .A(n34124), .B(n42638), .Y(n43859) );
  XOR2XL U33767 ( .A(n34128), .B(n36863), .Y(n43855) );
  XOR2XL U33768 ( .A(n34152), .B(n34450), .Y(n43979) );
  NOR2X1 U33769 ( .A(n23605), .B(n23604), .Y(n45719) );
  NOR2X1 U33770 ( .A(n22451), .B(n22450), .Y(n46100) );
  NOR2X1 U33771 ( .A(n23728), .B(n23727), .Y(n45697) );
  XOR2XL U33772 ( .A(n34349), .B(n36832), .Y(n45159) );
  XOR2XL U33773 ( .A(n34237), .B(n42547), .Y(n44786) );
  XOR2XL U33774 ( .A(n34348), .B(n36827), .Y(n45162) );
  XOR2XL U33775 ( .A(n34140), .B(n36829), .Y(n44004) );
  XOR2XL U33776 ( .A(n36767), .B(n33409), .Y(n46709) );
  XOR2XL U33777 ( .A(n36766), .B(n33401), .Y(n46714) );
  XOR2XL U33778 ( .A(n33409), .B(n36784), .Y(n45915) );
  NOR2XL U33779 ( .A(n12388), .B(n47098), .Y(n47102) );
  NOR2X1 U33780 ( .A(n23148), .B(n23147), .Y(n45861) );
  NOR2XL U33781 ( .A(n11210), .B(n47083), .Y(n47087) );
  XOR2XL U33782 ( .A(n34340), .B(n36821), .Y(n45131) );
  XNOR2XL U33783 ( .A(n33466), .B(n42569), .Y(net215904) );
  NAND4X2 U33784 ( .A(n43768), .B(n43767), .C(n43766), .D(n43765), .Y(n12024)
         );
  XNOR2XL U33785 ( .A(n33482), .B(n42558), .Y(n43767) );
  NOR2XL U33786 ( .A(n11200), .B(n47902), .Y(n47906) );
  XOR2XL U33787 ( .A(n34246), .B(n36868), .Y(n44766) );
  XOR2XL U33788 ( .A(n34214), .B(n36868), .Y(n44735) );
  NOR2X1 U33789 ( .A(n22898), .B(n22897), .Y(n45947) );
  NOR2X1 U33790 ( .A(n22857), .B(n22855), .Y(n45987) );
  INVXL U33791 ( .A(n47761), .Y(n47708) );
  CLKBUFX3 U33792 ( .A(net218260), .Y(net218144) );
  CLKBUFX3 U33793 ( .A(net218252), .Y(net218160) );
  CLKBUFX3 U33794 ( .A(net218222), .Y(net218218) );
  CLKBUFX3 U33795 ( .A(net218282), .Y(net218266) );
  CLKBUFX3 U33796 ( .A(net217256), .Y(net217248) );
  CLKBUFX3 U33797 ( .A(net217256), .Y(net217246) );
  CLKBUFX3 U33798 ( .A(net217254), .Y(net217252) );
  CLKBUFX3 U33799 ( .A(net217270), .Y(net217220) );
  CLKBUFX3 U33800 ( .A(net218282), .Y(net218262) );
  CLKBUFX3 U33801 ( .A(net218282), .Y(net218264) );
  CLKBUFX3 U33802 ( .A(n43024), .Y(n43023) );
  CLKBUFX3 U33803 ( .A(net218262), .Y(net218286) );
  CLKBUFX3 U33804 ( .A(n43034), .Y(n43031) );
  CLKBUFX3 U33805 ( .A(net217286), .Y(net217282) );
  CLKBUFX3 U33806 ( .A(net218966), .Y(net218956) );
  CLKBUFX3 U33807 ( .A(net221980), .Y(net221894) );
  CLKINVX2 U33808 ( .A(n42571), .Y(n42565) );
  CLKBUFX3 U33809 ( .A(n42497), .Y(n42495) );
  CLKINVX1 U33810 ( .A(net236115), .Y(n9782) );
  CLKINVX1 U33811 ( .A(n10437), .Y(net210705) );
  INVXL U33812 ( .A(n11645), .Y(net151248) );
  INVXL U33813 ( .A(n10381), .Y(net151348) );
  OAI211X2 U33814 ( .A0(n11775), .A1(n11776), .B0(n11777), .C0(n11778), .Y(
        n11772) );
  OAI21XL U33815 ( .A0(net171309), .A1(net209503), .B0(n11718), .Y(n48379) );
  AOI21X1 U33816 ( .A0(n48279), .A1(n12501), .B0(net171211), .Y(n48280) );
  NAND3XL U33817 ( .A(n11743), .B(n12530), .C(n11850), .Y(n48355) );
  OR2XL U33818 ( .A(n44571), .B(n44570), .Y(net207642) );
  INVXL U33819 ( .A(n11710), .Y(n48275) );
  NOR2BX1 U33820 ( .AN(n9851), .B(n42735), .Y(n9770) );
  NAND2X1 U33821 ( .A(net172112), .B(n9747), .Y(n10197) );
  INVXL U33822 ( .A(net210426), .Y(net210424) );
  OA21X4 U33823 ( .A0(n47770), .A1(net210596), .B0(net210597), .Y(n41751) );
  NOR2X1 U33824 ( .A(n48184), .B(net209885), .Y(n48167) );
  NOR4X4 U33825 ( .A(n28212), .B(n28213), .C(n28214), .D(n28215), .Y(n43778)
         );
  NOR4X4 U33826 ( .A(n28302), .B(n28303), .C(n28304), .D(n28305), .Y(n43751)
         );
  NAND4X2 U33827 ( .A(n43581), .B(n43580), .C(n43579), .D(n43578), .Y(n12539)
         );
  NAND4X2 U33828 ( .A(n43672), .B(n43671), .C(n43670), .D(n43669), .Y(n12530)
         );
  NOR3XL U33829 ( .A(net209620), .B(n48306), .C(n48302), .Y(n48303) );
  INVXL U33830 ( .A(n48307), .Y(n48302) );
  NOR4X2 U33831 ( .A(n29376), .B(n29377), .C(n29378), .D(n29379), .Y(n43571)
         );
  OR4X2 U33832 ( .A(n29192), .B(n29193), .C(n29194), .D(n29195), .Y(n41669) );
  NOR4X2 U33833 ( .A(n28049), .B(n28050), .C(n28051), .D(n28052), .Y(net215827) );
  NOR4X2 U33834 ( .A(n28053), .B(n28054), .C(n28055), .D(n28056), .Y(net215828) );
  OR2X4 U33835 ( .A(n29136), .B(n29145), .Y(n41755) );
  NAND4X2 U33836 ( .A(n44555), .B(n44554), .C(n44553), .D(n44552), .Y(n11712)
         );
  NAND4X2 U33837 ( .A(n44172), .B(n44171), .C(n44170), .D(n44169), .Y(n12582)
         );
  OR2X1 U33838 ( .A(n29167), .B(n29175), .Y(n41756) );
  CLKBUFX2 U33839 ( .A(n42726), .Y(n42727) );
  NOR4X4 U33840 ( .A(n28122), .B(n28123), .C(n28124), .D(n28125), .Y(n43805)
         );
  NOR4X2 U33841 ( .A(n28392), .B(n28393), .C(n28394), .D(n28395), .Y(n43732)
         );
  NAND4X2 U33842 ( .A(n43329), .B(n43328), .C(n43327), .D(n43326), .Y(n10090)
         );
  OR4X2 U33843 ( .A(n31118), .B(n31119), .C(n31120), .D(n31121), .Y(n41679) );
  NAND4X1 U33844 ( .A(n43067), .B(n43066), .C(n43065), .D(n43064), .Y(n12459)
         );
  NAND4X1 U33845 ( .A(n43048), .B(n43047), .C(n43046), .D(n43045), .Y(n12457)
         );
  NAND4X1 U33846 ( .A(n43130), .B(n43129), .C(n43128), .D(n43127), .Y(n12461)
         );
  NAND4X1 U33847 ( .A(n44589), .B(n44588), .C(n44587), .D(n44586), .Y(
        net214669) );
  INVX1 U33848 ( .A(n10686), .Y(net151479) );
  NAND4X1 U33849 ( .A(n43404), .B(n43403), .C(n43402), .D(n43401), .Y(n12449)
         );
  INVX1 U33850 ( .A(n10819), .Y(net151452) );
  NOR3XL U33851 ( .A(net151462), .B(n10686), .C(n10020), .Y(n21446) );
  OR2XL U33852 ( .A(n36935), .B(n41199), .Y(n9719) );
  OR2X1 U33853 ( .A(net218610), .B(n10198), .Y(n9872) );
  CLKBUFX3 U33854 ( .A(net151225), .Y(net221990) );
  OAI211X2 U33855 ( .A0(n11429), .A1(n11430), .B0(n10724), .C0(n10727), .Y(
        n11426) );
  XOR2X1 U33856 ( .A(n41813), .B(n36901), .Y(n45117) );
  XOR2X1 U33857 ( .A(n42057), .B(n42592), .Y(n45018) );
  OAI211X2 U33858 ( .A0(n11435), .A1(n11436), .B0(n10730), .C0(n10732), .Y(
        n11432) );
  INVXL U33859 ( .A(n11422), .Y(net151593) );
  XOR2X1 U33860 ( .A(n41798), .B(n42637), .Y(n45014) );
  OR4X4 U33861 ( .A(n45469), .B(n45468), .C(n45467), .D(n45466), .Y(n41683) );
  XNOR2XL U33862 ( .A(n36755), .B(n41810), .Y(n47660) );
  NOR2X2 U33863 ( .A(n46249), .B(net209868), .Y(n46259) );
  NOR2X2 U33864 ( .A(n43968), .B(n48334), .Y(n43978) );
  NOR2X2 U33865 ( .A(n44693), .B(net210670), .Y(n44703) );
  NOR2X2 U33866 ( .A(n43906), .B(n48288), .Y(n43916) );
  NAND4X4 U33867 ( .A(n44661), .B(n44660), .C(n44659), .D(n44658), .Y(n48325)
         );
  XOR2XL U33868 ( .A(n41808), .B(n36897), .Y(n44889) );
  XNOR2X1 U33869 ( .A(n49513), .B(n36865), .Y(n27721) );
  NAND4X2 U33870 ( .A(n43936), .B(n43935), .C(n43934), .D(n43933), .Y(
        net209572) );
  CLKINVX3 U33871 ( .A(n12007), .Y(net209781) );
  XOR2XL U33872 ( .A(n41831), .B(n36891), .Y(n44142) );
  XOR2XL U33873 ( .A(n36757), .B(n41822), .Y(n47347) );
  XOR2XL U33874 ( .A(n42091), .B(n42658), .Y(n44138) );
  XOR2XL U33875 ( .A(n42063), .B(n42672), .Y(n43892) );
  XOR2XL U33876 ( .A(n41804), .B(net219336), .Y(n43896) );
  XOR2XL U33877 ( .A(n42058), .B(n34450), .Y(n43886) );
  XOR2X1 U33878 ( .A(n41817), .B(n42523), .Y(n45409) );
  XOR2X1 U33879 ( .A(n42125), .B(n42652), .Y(n29169) );
  XNOR2X1 U33880 ( .A(n50996), .B(n42615), .Y(n27237) );
  XNOR2X1 U33881 ( .A(n50944), .B(n42617), .Y(n24742) );
  XNOR2X1 U33882 ( .A(n50364), .B(n42674), .Y(n27241) );
  XNOR2X1 U33883 ( .A(n50312), .B(n42672), .Y(n24746) );
  XNOR2X1 U33884 ( .A(n50945), .B(net219310), .Y(n24750) );
  XNOR2X1 U33885 ( .A(n51423), .B(n42641), .Y(n27243) );
  XNOR2X1 U33886 ( .A(n50782), .B(n36863), .Y(n27239) );
  XNOR2X1 U33887 ( .A(n51371), .B(n36867), .Y(n24748) );
  XNOR2X1 U33888 ( .A(n50730), .B(n36863), .Y(n24744) );
  XNOR2X1 U33889 ( .A(n51188), .B(n34447), .Y(n29012) );
  XNOR2X1 U33890 ( .A(n51210), .B(n42630), .Y(n27238) );
  XNOR2X1 U33891 ( .A(n51158), .B(n42631), .Y(n24743) );
  XNOR2X1 U33892 ( .A(n50568), .B(n36834), .Y(n27242) );
  XNOR2X1 U33893 ( .A(n50516), .B(n36728), .Y(n24747) );
  XNOR2XL U33894 ( .A(n50542), .B(n42717), .Y(n26858) );
  XOR2XL U33895 ( .A(n42157), .B(n36888), .Y(n25117) );
  NAND2X1 U33896 ( .A(n41768), .B(n41769), .Y(n45687) );
  XNOR2XL U33897 ( .A(n41852), .B(n42525), .Y(n41769) );
  XNOR2X1 U33898 ( .A(n50772), .B(n42501), .Y(n29154) );
  INVXL U33899 ( .A(n11029), .Y(net209171) );
  INVXL U33900 ( .A(n12264), .Y(net209176) );
  OAI21X1 U33901 ( .A0(net209176), .A1(n48535), .B0(n12260), .Y(n48536) );
  INVXL U33902 ( .A(n12741), .Y(net209840) );
  OAI21XL U33903 ( .A0(n39561), .A1(n48120), .B0(n12796), .Y(n48121) );
  NAND4XL U33904 ( .A(n48456), .B(net209296), .C(n48455), .D(net209298), .Y(
        n48457) );
  NAND3X4 U33905 ( .A(n44302), .B(n44301), .C(n44300), .Y(n12063) );
  XOR2XL U33906 ( .A(n42157), .B(n42656), .Y(n25139) );
  AO21X2 U33907 ( .A0(n48121), .A1(n12034), .B0(net209964), .Y(n41689) );
  AOI21XL U33908 ( .A0(n48432), .A1(n11147), .B0(n48431), .Y(n48480) );
  CLKINVX1 U33909 ( .A(n12151), .Y(net209971) );
  AOI21X1 U33910 ( .A0(n48074), .A1(n11396), .B0(net171540), .Y(n48075) );
  INVXL U33911 ( .A(n48138), .Y(n48139) );
  INVXL U33912 ( .A(n48172), .Y(n48176) );
  NOR2BX1 U33913 ( .AN(n11410), .B(n13016), .Y(n48064) );
  INVX3 U33914 ( .A(n47967), .Y(n48062) );
  OAI2BB1X2 U33915 ( .A0N(n10709), .A1N(net210238), .B0(n10708), .Y(n47967) );
  XOR2X1 U33916 ( .A(n42100), .B(n36877), .Y(n43909) );
  XOR2XL U33917 ( .A(n41801), .B(n41283), .Y(n43897) );
  XOR2XL U33918 ( .A(n41899), .B(n36900), .Y(n24993) );
  XOR2XL U33919 ( .A(n42159), .B(n42655), .Y(n24989) );
  XOR2XL U33920 ( .A(n41900), .B(n42608), .Y(n24985) );
  XOR2XL U33921 ( .A(n42092), .B(n36873), .Y(n44156) );
  XOR2XL U33922 ( .A(n36809), .B(n42076), .Y(n46346) );
  XOR2X1 U33923 ( .A(n41849), .B(n36895), .Y(n27459) );
  OR2X1 U33924 ( .A(n29153), .B(n29176), .Y(n43603) );
  OAI2BB1XL U33925 ( .A0N(net209903), .A1N(n41777), .B0(net209898), .Y(n48164)
         );
  AO21XL U33926 ( .A0(net209899), .A1(net209900), .B0(net209901), .Y(n41777)
         );
  OAI2BB1XL U33927 ( .A0N(n48160), .A1N(n41775), .B0(net209930), .Y(n48141) );
  AO21XL U33928 ( .A0(n48140), .A1(n48159), .B0(n48139), .Y(n41775) );
  NAND2XL U33929 ( .A(net209312), .B(net209313), .Y(n48451) );
  XOR2X1 U33930 ( .A(n41871), .B(n41309), .Y(n22429) );
  INVXL U33931 ( .A(net209284), .Y(net209283) );
  XNOR2X1 U33932 ( .A(n51350), .B(n42701), .Y(n31613) );
  XNOR2X1 U33933 ( .A(n51135), .B(n42550), .Y(n31590) );
  XNOR2X1 U33934 ( .A(n50760), .B(n42592), .Y(n29013) );
  XNOR2X1 U33935 ( .A(n50707), .B(n42499), .Y(n31591) );
  XOR2X1 U33936 ( .A(n42190), .B(n42667), .Y(n31606) );
  XOR2X1 U33937 ( .A(n41931), .B(n42608), .Y(n31602) );
  XNOR2X1 U33938 ( .A(n51401), .B(n42644), .Y(n29017) );
  XNOR2X1 U33939 ( .A(n50921), .B(n42538), .Y(n31589) );
  XOR2X1 U33940 ( .A(n41932), .B(n42519), .Y(n31592) );
  XOR2X1 U33941 ( .A(n41930), .B(n36892), .Y(n31610) );
  XOR2X1 U33942 ( .A(n42189), .B(n36888), .Y(n31614) );
  XOR2X1 U33943 ( .A(n42130), .B(n36813), .Y(n22430) );
  XOR2X1 U33944 ( .A(n42191), .B(n36877), .Y(n31593) );
  NOR4X1 U33945 ( .A(n29049), .B(n29050), .C(n29051), .D(n29052), .Y(n43662)
         );
  XNOR2XL U33946 ( .A(n50728), .B(net219468), .Y(n28150) );
  INVXL U33947 ( .A(n10879), .Y(net209259) );
  OAI2BB1XL U33948 ( .A0N(n11140), .A1N(net209259), .B0(n11139), .Y(n48481) );
  INVX1 U33949 ( .A(n12064), .Y(n48128) );
  INVX1 U33950 ( .A(n12025), .Y(net209958) );
  NAND2XL U33951 ( .A(n48000), .B(n47995), .Y(n48003) );
  XOR2XL U33952 ( .A(n41892), .B(n41314), .Y(n24099) );
  XOR2XL U33953 ( .A(n41868), .B(n41313), .Y(n22439) );
  XOR2XL U33954 ( .A(n41908), .B(n41313), .Y(n23603) );
  XOR2XL U33955 ( .A(n36734), .B(n42063), .Y(n47547) );
  OAI2BB1X1 U33956 ( .A0N(n12322), .A1N(n41782), .B0(n12323), .Y(n48425) );
  OAI2BB1XL U33957 ( .A0N(n11058), .A1N(n41784), .B0(n12280), .Y(n48525) );
  AO21XL U33958 ( .A0(n48523), .A1(n48522), .B0(net209197), .Y(n41784) );
  XNOR2X1 U33959 ( .A(n50906), .B(n42620), .Y(n31840) );
  XNOR2X1 U33960 ( .A(n50274), .B(n42672), .Y(n31844) );
  XNOR2X1 U33961 ( .A(n50692), .B(n42589), .Y(n31842) );
  XNOR2X1 U33962 ( .A(n51120), .B(n42626), .Y(n31841) );
  XNOR2X1 U33963 ( .A(n50480), .B(n36903), .Y(n31845) );
  NOR4BX1 U33964 ( .AN(n41714), .B(n19808), .C(n19807), .D(n19806), .Y(n47155)
         );
  CLKINVX3 U33965 ( .A(net213021), .Y(net171124) );
  INVXL U33966 ( .A(n11051), .Y(net171461) );
  INVXL U33967 ( .A(n12311), .Y(net171417) );
  INVXL U33968 ( .A(n11116), .Y(net209355) );
  XOR2XL U33969 ( .A(n41909), .B(n36761), .Y(n21100) );
  XOR2XL U33970 ( .A(n41893), .B(n36761), .Y(n19739) );
  XOR2XL U33971 ( .A(n42168), .B(n42484), .Y(n21101) );
  XOR2XL U33972 ( .A(n41889), .B(n36754), .Y(n19799) );
  XOR2XL U33973 ( .A(n41915), .B(n41318), .Y(n23206) );
  XOR2XL U33974 ( .A(n41929), .B(n36756), .Y(n21604) );
  XOR2XL U33975 ( .A(n42152), .B(n42489), .Y(n19740) );
  XOR2XL U33976 ( .A(n42174), .B(n36807), .Y(n23207) );
  XOR2XL U33977 ( .A(n42188), .B(n42489), .Y(n21605) );
  XNOR2X1 U33978 ( .A(n51318), .B(n42697), .Y(n32095) );
  XOR2XL U33979 ( .A(n41933), .B(n36756), .Y(n21504) );
  XOR2XL U33980 ( .A(n42192), .B(n42486), .Y(n21505) );
  NOR3X1 U33981 ( .A(n46485), .B(n46484), .C(n46483), .Y(n46486) );
  XOR2XL U33982 ( .A(n36782), .B(n34369), .Y(n41722) );
  XOR2XL U33983 ( .A(n36784), .B(n34361), .Y(n41723) );
  XOR2X1 U33984 ( .A(n34419), .B(n36879), .Y(n45005) );
  XOR2X1 U33985 ( .A(n34317), .B(n42549), .Y(n45415) );
  XOR2X1 U33986 ( .A(n34318), .B(n42534), .Y(n45414) );
  XNOR2XL U33987 ( .A(n9660), .B(n36875), .Y(n41725) );
  XOR2X1 U33988 ( .A(n42077), .B(n36879), .Y(n45505) );
  NOR2X1 U33989 ( .A(n23789), .B(n23788), .Y(n46207) );
  NOR4X1 U33990 ( .A(n23787), .B(n23786), .C(n23785), .D(n23784), .Y(n46206)
         );
  XOR2XL U33991 ( .A(n34377), .B(n42717), .Y(n44961) );
  XOR2XL U33992 ( .A(n34385), .B(n34435), .Y(n44925) );
  NOR4X1 U33993 ( .A(n47397), .B(n47396), .C(n47395), .D(n47394), .Y(n47398)
         );
  XNOR2XL U33994 ( .A(n34192), .B(n42504), .Y(n44162) );
  NOR4X2 U33995 ( .A(n45518), .B(n45517), .C(n45516), .D(n45515), .Y(net213703) );
  XOR2XL U33996 ( .A(n36789), .B(n34398), .Y(n47700) );
  NOR4X2 U33997 ( .A(n45373), .B(n45372), .C(n45371), .D(n45370), .Y(n45374)
         );
  NOR2X2 U33998 ( .A(n45369), .B(n45368), .Y(n45375) );
  XNOR2XL U33999 ( .A(n42473), .B(n34288), .Y(n47345) );
  XOR2XL U34000 ( .A(n34430), .B(n42534), .Y(n45231) );
  XOR2X1 U34001 ( .A(n42620), .B(n34126), .Y(n43857) );
  XOR2XL U34002 ( .A(n34197), .B(n42625), .Y(n44136) );
  XOR2XL U34003 ( .A(n34194), .B(n36907), .Y(n44139) );
  XOR2XL U34004 ( .A(n34198), .B(n41284), .Y(n44135) );
  XOR2X1 U34005 ( .A(n34423), .B(n36898), .Y(n45009) );
  XOR2XL U34006 ( .A(n34330), .B(n41630), .Y(n45223) );
  OR3X2 U34007 ( .A(n45067), .B(n45070), .C(n45069), .Y(n41734) );
  NOR2X1 U34008 ( .A(n45728), .B(n45727), .Y(n45732) );
  NAND4X4 U34009 ( .A(n43554), .B(n43553), .C(n43552), .D(n43551), .Y(n12147)
         );
  NAND4X4 U34010 ( .A(n43824), .B(n43823), .C(n43822), .D(n43821), .Y(n48188)
         );
  NAND4X4 U34011 ( .A(n43704), .B(n43703), .C(n43702), .D(n43701), .Y(n12797)
         );
  NOR2X2 U34012 ( .A(n25157), .B(n25156), .Y(n44437) );
  NAND4X4 U34013 ( .A(n44197), .B(n44196), .C(n44195), .D(n44194), .Y(n12749)
         );
  NOR2X2 U34014 ( .A(n26690), .B(n26689), .Y(n46174) );
  NOR4X1 U34015 ( .A(n20247), .B(n20246), .C(n20245), .D(n20244), .Y(net211516) );
  NOR4X1 U34016 ( .A(n47516), .B(n47515), .C(n47514), .D(n47513), .Y(n47517)
         );
  NOR2X1 U34017 ( .A(n20413), .B(n20412), .Y(n47564) );
  NOR4X1 U34018 ( .A(n20411), .B(n20410), .C(n20409), .D(n20408), .Y(n47563)
         );
  NAND4X4 U34019 ( .A(n43643), .B(n43642), .C(n43641), .D(n43640), .Y(n12736)
         );
  NOR4X1 U34020 ( .A(n47485), .B(n47484), .C(n47483), .D(n47482), .Y(n47486)
         );
  NOR2X1 U34021 ( .A(n20291), .B(n20290), .Y(n47288) );
  NOR2X1 U34022 ( .A(n20147), .B(n20146), .Y(n47033) );
  XOR2XL U34023 ( .A(n36765), .B(n34033), .Y(n47017) );
  NOR2X4 U34024 ( .A(n11756), .B(n43573), .Y(n43577) );
  NOR2X4 U34025 ( .A(n10422), .B(n44267), .Y(net215289) );
  NOR2X4 U34026 ( .A(n11751), .B(n43559), .Y(n43563) );
  XOR2X1 U34027 ( .A(n33604), .B(n36825), .Y(n44521) );
  NOR2X4 U34028 ( .A(n10384), .B(n44212), .Y(n44216) );
  XOR2XL U34029 ( .A(n36780), .B(n34313), .Y(n46347) );
  XOR2XL U34030 ( .A(n34205), .B(n41282), .Y(n44144) );
  XOR2XL U34031 ( .A(n34124), .B(n42698), .Y(n43846) );
  XOR2XL U34032 ( .A(n34206), .B(net219310), .Y(n44143) );
  XOR2XL U34033 ( .A(n34196), .B(n42637), .Y(n44137) );
  XOR2XL U34034 ( .A(n34200), .B(n34450), .Y(n44133) );
  XOR2XL U34035 ( .A(n34188), .B(n36831), .Y(n44158) );
  XOR2XL U34036 ( .A(n36741), .B(n34308), .Y(n47308) );
  XOR2XL U34037 ( .A(n34189), .B(n42547), .Y(n44155) );
  NOR2X1 U34038 ( .A(n46945), .B(net209225), .Y(n46949) );
  NOR2X1 U34039 ( .A(n47209), .B(net211271), .Y(n47213) );
  XNOR2XL U34040 ( .A(n36837), .B(n33538), .Y(n45831) );
  NOR2X1 U34041 ( .A(n19841), .B(n19840), .Y(n47141) );
  NOR4X1 U34042 ( .A(n19839), .B(n19838), .C(n19837), .D(n19836), .Y(n47140)
         );
  NOR2X1 U34043 ( .A(n22371), .B(n22370), .Y(n46130) );
  NAND4X4 U34044 ( .A(n46132), .B(n46131), .C(n46130), .D(n46129), .Y(n12322)
         );
  NOR4X1 U34045 ( .A(n21090), .B(n21089), .C(n21088), .D(n21087), .Y(n46921)
         );
  NOR2X1 U34046 ( .A(n19952), .B(n19951), .Y(n47080) );
  NOR4X1 U34047 ( .A(n19950), .B(n19949), .C(n19948), .D(n19947), .Y(n47079)
         );
  NOR2X1 U34048 ( .A(n23453), .B(n23452), .Y(n45785) );
  NOR4X1 U34049 ( .A(n23451), .B(n23450), .C(n23449), .D(n23448), .Y(n45784)
         );
  NOR2X1 U34050 ( .A(n19761), .B(n19760), .Y(n47171) );
  NOR4X1 U34051 ( .A(n19759), .B(n19758), .C(n19757), .D(n19756), .Y(n47170)
         );
  NOR2X1 U34052 ( .A(n19851), .B(n19850), .Y(n47136) );
  NAND4X2 U34053 ( .A(n45919), .B(n45918), .C(n45917), .D(n45916), .Y(n11058)
         );
  NOR2X1 U34054 ( .A(n21596), .B(n21595), .Y(n46711) );
  NOR4X1 U34055 ( .A(n21594), .B(n21593), .C(n21592), .D(n21591), .Y(n46710)
         );
  NOR2X1 U34056 ( .A(n19872), .B(n19871), .Y(n47120) );
  NOR4X1 U34057 ( .A(n19870), .B(n19869), .C(n19868), .D(n19867), .Y(n47119)
         );
  NOR2X1 U34058 ( .A(n20117), .B(n20115), .Y(net211485) );
  NOR2X1 U34059 ( .A(n19781), .B(n19780), .Y(n47884) );
  NOR4X1 U34060 ( .A(n19779), .B(n19778), .C(n19777), .D(n19776), .Y(n47883)
         );
  NAND4X2 U34061 ( .A(n45699), .B(n45698), .C(n45697), .D(n45696), .Y(n11131)
         );
  XNOR2XL U34062 ( .A(n36735), .B(n33706), .Y(n47182) );
  NOR2X1 U34063 ( .A(n22471), .B(n22470), .Y(n46090) );
  XOR2XL U34064 ( .A(n36750), .B(n33572), .Y(n46920) );
  NOR2XL U34065 ( .A(n11132), .B(n47041), .Y(net211488) );
  XOR2XL U34066 ( .A(n36773), .B(n33825), .Y(n47149) );
  XOR2XL U34067 ( .A(n36765), .B(n33585), .Y(n47853) );
  NOR2X1 U34068 ( .A(n47053), .B(n48521), .Y(n47057) );
  XNOR2XL U34069 ( .A(n33306), .B(n42569), .Y(n43333) );
  NOR4X1 U34070 ( .A(n31172), .B(n31171), .C(n31170), .D(n31169), .Y(n43331)
         );
  NOR2X1 U34071 ( .A(n21526), .B(n21525), .Y(n46746) );
  NOR4X1 U34072 ( .A(n21524), .B(n21523), .C(n21522), .D(n21521), .Y(n46745)
         );
  NOR2X1 U34073 ( .A(n21576), .B(n21575), .Y(n46721) );
  NOR4X1 U34074 ( .A(n21574), .B(n21573), .C(n21572), .D(n21571), .Y(n46720)
         );
  NOR4X1 U34075 ( .A(n22896), .B(n22895), .C(n22894), .D(n22893), .Y(n45946)
         );
  NOR2X1 U34076 ( .A(n21496), .B(n21495), .Y(n46771) );
  NOR4X1 U34077 ( .A(n21494), .B(n21493), .C(n21492), .D(n21491), .Y(n46770)
         );
  NOR2X1 U34078 ( .A(n43168), .B(net209476), .Y(n43172) );
  NOR2X1 U34079 ( .A(n10089), .B(n43312), .Y(n43316) );
  NOR2X1 U34080 ( .A(n10090), .B(n43330), .Y(n43334) );
  NOR2X1 U34081 ( .A(n11018), .B(n46809), .Y(n46813) );
  NOR2X1 U34082 ( .A(n12251), .B(n46799), .Y(n46803) );
  NOR2X1 U34083 ( .A(n11034), .B(n46895), .Y(n46899) );
  NOR4X1 U34084 ( .A(n22854), .B(n22853), .C(n22852), .D(n22851), .Y(n45986)
         );
  NOR2X1 U34085 ( .A(n10820), .B(n46688), .Y(net211987) );
  NOR2X1 U34086 ( .A(n11007), .B(n46819), .Y(n46823) );
  NOR2X1 U34087 ( .A(n10273), .B(n46689), .Y(net211982) );
  NOR2X1 U34088 ( .A(n12246), .B(n46834), .Y(n46838) );
  NOR2X1 U34089 ( .A(n22755), .B(n22754), .Y(n46012) );
  NAND4X1 U34090 ( .A(n46014), .B(n46013), .C(n46012), .D(n46011), .Y(n11218)
         );
  NOR2X1 U34091 ( .A(n22735), .B(n22734), .Y(n46022) );
  CLKBUFX3 U34092 ( .A(n33127), .Y(n41966) );
  CLKBUFX3 U34093 ( .A(n33119), .Y(n41967) );
  CLKBUFX3 U34094 ( .A(n33111), .Y(n41968) );
  CLKBUFX3 U34095 ( .A(n33103), .Y(n41969) );
  CLKBUFX3 U34096 ( .A(n33095), .Y(n41970) );
  CLKBUFX3 U34097 ( .A(n33087), .Y(n41971) );
  CLKBUFX3 U34098 ( .A(n33071), .Y(n41973) );
  CLKBUFX3 U34099 ( .A(n33063), .Y(n41974) );
  CLKBUFX3 U34100 ( .A(n33123), .Y(n42225) );
  CLKBUFX3 U34101 ( .A(n33115), .Y(n42226) );
  CLKBUFX3 U34102 ( .A(n33107), .Y(n42227) );
  CLKBUFX3 U34103 ( .A(n33099), .Y(n42228) );
  CLKBUFX3 U34104 ( .A(n33091), .Y(n42229) );
  CLKBUFX3 U34105 ( .A(n33083), .Y(n42230) );
  CLKBUFX3 U34106 ( .A(n33067), .Y(n42232) );
  CLKBUFX3 U34107 ( .A(n33059), .Y(n42233) );
  AOI2BB2XL U34108 ( .B0(n9748), .B1(n9715), .A0N(n9737), .A1N(n37241), .Y(
        n9738) );
  CLKBUFX3 U34109 ( .A(n33015), .Y(n41980) );
  CLKBUFX3 U34110 ( .A(n33007), .Y(n41981) );
  CLKBUFX3 U34111 ( .A(n32999), .Y(n41982) );
  CLKBUFX3 U34112 ( .A(n32991), .Y(n41983) );
  CLKBUFX3 U34113 ( .A(n33011), .Y(n42239) );
  CLKBUFX3 U34114 ( .A(n33003), .Y(n42240) );
  CLKBUFX3 U34115 ( .A(n32995), .Y(n42241) );
  CLKBUFX3 U34116 ( .A(n32987), .Y(n42242) );
  AOI2BB2XL U34117 ( .B0(n9873), .B1(n9773), .A0N(n36885), .A1N(net218220),
        .Y(n9807) );
  CLKBUFX3 U34118 ( .A(n33047), .Y(n41976) );
  CLKBUFX3 U34119 ( .A(n33039), .Y(n41977) );
  CLKBUFX3 U34120 ( .A(n33031), .Y(n41978) );
  CLKBUFX3 U34121 ( .A(n33023), .Y(n41979) );
  CLKBUFX3 U34122 ( .A(n33043), .Y(n42235) );
  CLKBUFX3 U34123 ( .A(n33035), .Y(n42236) );
  CLKBUFX3 U34124 ( .A(n33027), .Y(n42237) );
  CLKBUFX3 U34125 ( .A(n33019), .Y(n42238) );
  CLKBUFX3 U34126 ( .A(n33079), .Y(n41972) );
  CLKBUFX3 U34127 ( .A(n33055), .Y(n41975) );
  CLKBUFX3 U34128 ( .A(n33075), .Y(n42231) );
  CLKBUFX3 U34129 ( .A(n33051), .Y(n42234) );
  NAND2X1 U34130 ( .A(n34374), .B(n41656), .Y(n41657) );
  NAND2XL U34131 ( .A(n41655), .B(n36868), .Y(n41658) );
  CLKBUFX3 U34132 ( .A(net218252), .Y(net218158) );
  INVX1 U34133 ( .A(n43010), .Y(n42991) );
  CLKBUFX3 U34134 ( .A(net217248), .Y(net217120) );
  CLKBUFX3 U34135 ( .A(net217250), .Y(net217116) );
  CLKBUFX3 U34136 ( .A(net217250), .Y(net217114) );
  CLKBUFX3 U34137 ( .A(net217248), .Y(net217118) );
  CLKBUFX3 U34138 ( .A(net217252), .Y(net217112) );
  CLKBUFX2 U34139 ( .A(net218222), .Y(net218220) );
  BUFX2 U34140 ( .A(net218276), .Y(net218230) );
  BUFX2 U34141 ( .A(net217254), .Y(net217250) );
  BUFX2 U34142 ( .A(net218284), .Y(net218268) );
  BUFX2 U34143 ( .A(net217266), .Y(net217226) );
  BUFX2 U34144 ( .A(net217258), .Y(net217242) );
  BUFX2 U34145 ( .A(net217270), .Y(net217218) );
  CLKBUFX2 U34146 ( .A(net217276), .Y(net217206) );
  BUFX2 U34147 ( .A(net218948), .Y(net218888) );
  CLKBUFX2 U34148 ( .A(net218934), .Y(net218930) );
  CLKBUFX2 U34149 ( .A(net218934), .Y(net218928) );
  CLKBUFX2 U34150 ( .A(net218948), .Y(net218886) );
  CLKBUFX2 U34151 ( .A(net218948), .Y(net218890) );
  CLKBUFX2 U34152 ( .A(n43034), .Y(n43030) );
  CLKBUFX2 U34153 ( .A(n43034), .Y(n43029) );
  BUFX2 U34154 ( .A(net217288), .Y(net217278) );
  CLKBUFX2 U34155 ( .A(net217286), .Y(net217284) );
  BUFX2 U34156 ( .A(n9874), .Y(net218292) );
  BUFX2 U34157 ( .A(net218602), .Y(net218582) );
  CLKBUFX2 U34158 ( .A(net218602), .Y(net218586) );
  CLKBUFX2 U34159 ( .A(net218602), .Y(net218584) );
  BUFX2 U34160 ( .A(net218964), .Y(net218960) );
  CLKBUFX2 U34161 ( .A(net218966), .Y(net218958) );
  CLKBUFX2 U34162 ( .A(net218964), .Y(net218962) );
  CLKINVX2 U34163 ( .A(n42571), .Y(n42564) );
  CLKBUFX2 U34164 ( .A(n42530), .Y(n42521) );
  NOR3XL U34165 ( .A(net171255), .B(net171248), .C(net209517), .Y(n48361) );
  CLKINVX3 U34166 ( .A(n41222), .Y(n42566) );
  CLKBUFX2 U34167 ( .A(n42529), .Y(n42520) );
  CLKBUFX2 U34168 ( .A(n42472), .Y(n42462) );
  CLKBUFX2 U34169 ( .A(n42478), .Y(n42487) );
  CLKBUFX2 U34170 ( .A(n42472), .Y(n42461) );
  CLKBUFX2 U34171 ( .A(n42519), .Y(n42517) );
  NOR2XL U34172 ( .A(net171314), .B(net171231), .Y(n11771) );
  CLKBUFX2 U34173 ( .A(n42478), .Y(n42485) );
  NAND2BXL U34174 ( .AN(net210705), .B(net260384), .Y(n9852) );
  CLKINVX2 U34175 ( .A(n41222), .Y(n42567) );
  OA22XL U34176 ( .A0(net263330), .A1(n36748), .B0(n41299), .B1(net218918),
        .Y(n13063) );
  NOR4XL U34177 ( .A(n9812), .B(n9813), .C(n50120), .D(net217212), .Y(n9811)
         );
  NOR2XL U34178 ( .A(net171309), .B(net171300), .Y(n11713) );
  INVXL U34179 ( .A(net207653), .Y(net151394) );
  AND2XL U34180 ( .A(n10437), .B(n36928), .Y(net236115) );
  NOR2XL U34181 ( .A(net171140), .B(net171328), .Y(n11653) );
  NOR3BXL U34182 ( .AN(n10355), .B(n10357), .C(net171300), .Y(n10103) );
  AO21X2 U34183 ( .A0(n48386), .A1(n48385), .B0(n48384), .Y(n41659) );
  OA21XL U34184 ( .A0(n11686), .A1(n49506), .B0(n48387), .Y(n41660) );
  OAI2BB1XL U34185 ( .A0N(n10128), .A1N(n41661), .B0(n10126), .Y(n48297) );
  AO21XL U34186 ( .A0(n48296), .A1(net209565), .B0(net209642), .Y(n41661) );
  AOI21X2 U34187 ( .A0(n48287), .A1(n11743), .B0(n48286), .Y(n48366) );
  OAI2BB1X2 U34188 ( .A0N(n41662), .A1N(n41663), .B0(n48359), .Y(n48365) );
  AO21X2 U34189 ( .A0(n48347), .A1(n48346), .B0(n48345), .Y(n41662) );
  AO21X2 U34190 ( .A0(n48405), .A1(n11646), .B0(net209463), .Y(n41738) );
  OAI2BB1X2 U34191 ( .A0N(n11640), .A1N(n41738), .B0(n11637), .Y(n48406) );
  CLKBUFX2 U34192 ( .A(n42648), .Y(n42668) );
  OAI21X1 U34193 ( .A0(net171198), .A1(n48278), .B0(n11698), .Y(n48279) );
  INVX3 U34194 ( .A(n11763), .Y(net209537) );
  NAND2XL U34195 ( .A(net209565), .B(n48337), .Y(n48339) );
  NAND2XL U34196 ( .A(n11777), .B(n10128), .Y(n48338) );
  NAND2XL U34197 ( .A(n10377), .B(n10378), .Y(n48357) );
  NAND2XL U34198 ( .A(n11756), .B(n11751), .Y(n48356) );
  INVXL U34199 ( .A(n10368), .Y(net209529) );
  CLKBUFX2 U34200 ( .A(n42647), .Y(n42667) );
  NAND3XL U34201 ( .A(n11693), .B(n11688), .C(n12501), .Y(n48376) );
  NAND3XL U34202 ( .A(n12506), .B(n11710), .C(n11711), .Y(n48378) );
  NOR2XL U34203 ( .A(net171249), .B(net171255), .Y(n11734) );
  NOR2XL U34204 ( .A(net171101), .B(net171143), .Y(n11641) );
  NOR2XL U34205 ( .A(net171099), .B(net171104), .Y(n11631) );
  NAND2XL U34206 ( .A(n10128), .B(n10126), .Y(n11776) );
  NOR2BXL U34207 ( .AN(n48293), .B(n48295), .Y(n47752) );
  NAND2XL U34208 ( .A(n11711), .B(n11712), .Y(n11708) );
  NAND2XL U34209 ( .A(net209565), .B(net210460), .Y(n47750) );
  NOR2BXL U34210 ( .AN(n12538), .B(net171189), .Y(n11757) );
  NAND2XL U34211 ( .A(n11743), .B(n11744), .Y(n11740) );
  CLKINVX1 U34212 ( .A(net221990), .Y(net221982) );
  OAI211XL U34213 ( .A0(n9784), .A1(n9763), .B0(n49499), .C0(n9770), .Y(n9783)
         );
  NOR2BXL U34214 ( .AN(n48387), .B(n49506), .Y(n11679) );
  NOR4XL U34215 ( .A(n10061), .B(n10062), .C(n10063), .D(net217118), .Y(n10060) );
  NAND2X1 U34216 ( .A(net266255), .B(n41199), .Y(n10058) );
  INVX1 U34217 ( .A(n9759), .Y(n50086) );
  NOR2XL U34218 ( .A(n49505), .B(n49500), .Y(n11701) );
  NOR2XL U34219 ( .A(net171211), .B(net171196), .Y(n11689) );
  NAND2XL U34220 ( .A(n11733), .B(n10424), .Y(n11730) );
  CLKINVX1 U34221 ( .A(net221990), .Y(net221984) );
  CLKINVX1 U34222 ( .A(net221992), .Y(net221986) );
  NAND2XL U34223 ( .A(n12452), .B(n12455), .Y(n10079) );
  NAND4XL U34224 ( .A(n11709), .B(n12506), .C(n12586), .D(n11710), .Y(n10106)
         );
  NAND3X1 U34225 ( .A(n45526), .B(n45525), .C(n45524), .Y(n12592) );
  NAND2XL U34226 ( .A(net210523), .B(net234762), .Y(n47824) );
  CLKINVX1 U34227 ( .A(n9743), .Y(n50082) );
  NAND3BXL U34228 ( .AN(n10088), .B(n10089), .C(n10090), .Y(n10084) );
  NAND4XL U34229 ( .A(n10339), .B(n10341), .C(n10340), .D(n24678), .Y(n9828)
         );
  NOR2BXL U34230 ( .AN(net210473), .B(net210390), .Y(n41742) );
  NAND4X1 U34231 ( .A(n10306), .B(n10302), .C(n24712), .D(net259626), .Y(n9824) );
  NAND4XL U34232 ( .A(n10425), .B(net259641), .C(net259645), .D(n24680), .Y(
        n10075) );
  NAND4XL U34233 ( .A(n10367), .B(n10368), .C(n10369), .D(n24665), .Y(n10108)
         );
  NOR2XL U34234 ( .A(net171255), .B(n10421), .Y(n24665) );
  NAND4X1 U34235 ( .A(n11697), .B(n11688), .C(net151325), .D(n24722), .Y(n9792) );
  AND4XL U34236 ( .A(n10376), .B(n10377), .C(n10378), .D(n24670), .Y(n10110)
         );
  NOR2XL U34237 ( .A(net209661), .B(n10420), .Y(n24670) );
  NAND4X1 U34238 ( .A(net259661), .B(net259665), .C(n10433), .D(n24711), .Y(
        n9816) );
  AND4XL U34239 ( .A(n10362), .B(n11733), .C(n24667), .D(n10424), .Y(n10109)
         );
  NOR2XL U34240 ( .A(net151356), .B(net209517), .Y(n24667) );
  NAND4XL U34241 ( .A(n10393), .B(n10394), .C(n10395), .D(n24718), .Y(n9939)
         );
  AND3XL U34242 ( .A(net210462), .B(n10126), .C(n45531), .Y(n41743) );
  CLKINVX1 U34243 ( .A(n9748), .Y(n50114) );
  AND4X4 U34244 ( .A(n46572), .B(n46571), .C(n46570), .D(n46569), .Y(n41665)
         );
  OR4X4 U34245 ( .A(n26695), .B(n26696), .C(n26697), .D(n26698), .Y(n41666) );
  NAND4BX2 U34246 ( .AN(n41667), .B(n43836), .C(n43835), .D(n43834), .Y(n48337) );
  OR4X2 U34247 ( .A(n27689), .B(n27690), .C(n27691), .D(n27692), .Y(n41667) );
  NAND4X2 U34248 ( .A(n44520), .B(n44519), .C(n44518), .D(n44517), .Y(n11718)
         );
  NAND4X2 U34249 ( .A(n43828), .B(n43827), .C(n43826), .D(n43825), .Y(n48293)
         );
  NOR4X2 U34250 ( .A(n28144), .B(n28145), .C(n28146), .D(n28147), .Y(n43798)
         );
  NOR4X2 U34251 ( .A(n28152), .B(n28153), .C(n28154), .D(n28155), .Y(n43796)
         );
  INVXL U34252 ( .A(n48301), .Y(n48318) );
  OAI2BB1X2 U34253 ( .A0N(n41673), .A1N(n41674), .B0(n48341), .Y(n48346) );
  NAND4X2 U34254 ( .A(n44227), .B(n44226), .C(n44225), .D(n44224), .Y(n12542)
         );
  NAND4X4 U34255 ( .A(n43754), .B(n43753), .C(n43752), .D(n43751), .Y(n11688)
         );
  NAND4BX4 U34256 ( .AN(n41675), .B(n43647), .C(n43646), .D(n43645), .Y(n11850) );
  OR4X2 U34257 ( .A(n29101), .B(n29102), .C(n29103), .D(n29104), .Y(n41675) );
  NAND4X2 U34258 ( .A(n44493), .B(n44492), .C(n44491), .D(n44490), .Y(n11723)
         );
  NAND4X2 U34259 ( .A(n44459), .B(n44458), .C(n44457), .D(n44456), .Y(n44571)
         );
  NOR2X4 U34260 ( .A(n25112), .B(n25113), .Y(n44459) );
  NAND4X2 U34261 ( .A(n44447), .B(n44446), .C(n44445), .D(n44444), .Y(n47947)
         );
  NAND4X2 U34262 ( .A(n44443), .B(n44442), .C(n44441), .D(n44440), .Y(n47948)
         );
  NAND4XL U34263 ( .A(n41757), .B(net209589), .C(n48325), .D(n48321), .Y(
        n48322) );
  NOR2XL U34264 ( .A(net209250), .B(net171433), .Y(n48475) );
  INVXL U34265 ( .A(n48309), .Y(n48310) );
  CLKBUFX2 U34266 ( .A(n42511), .Y(n42528) );
  NAND4X2 U34267 ( .A(n43195), .B(n43194), .C(n43193), .D(n43192), .Y(n12490)
         );
  NAND4X2 U34268 ( .A(n43293), .B(n43292), .C(n43291), .D(n43290), .Y(n12486)
         );
  NOR4X2 U34269 ( .A(n31299), .B(n31300), .C(n31301), .D(n31302), .Y(n43293)
         );
  NOR4X2 U34270 ( .A(n31311), .B(n31312), .C(n31313), .D(n31314), .Y(n43290)
         );
  NAND4X2 U34271 ( .A(n44237), .B(n44236), .C(n44235), .D(n44234), .Y(n48370)
         );
  NAND4X2 U34272 ( .A(n43735), .B(n43734), .C(n43733), .D(n43732), .Y(n48383)
         );
  NOR4X2 U34273 ( .A(n31539), .B(n31540), .C(n31541), .D(n31542), .Y(n43222)
         );
  NOR4X2 U34274 ( .A(n31551), .B(n31552), .C(n31553), .D(n31554), .Y(n43219)
         );
  NAND4X2 U34275 ( .A(n43213), .B(n43212), .C(n43211), .D(n43210), .Y(n48387)
         );
  NAND4X4 U34276 ( .A(n43699), .B(n43698), .C(n43697), .D(n43696), .Y(n11697)
         );
  NAND4X4 U34277 ( .A(n43781), .B(n43780), .C(n43779), .D(n43778), .Y(n11699)
         );
  NAND4X4 U34278 ( .A(n43808), .B(n43807), .C(n43806), .D(n43805), .Y(n11706)
         );
  NOR4X2 U34279 ( .A(n29384), .B(n29385), .C(n29386), .D(n29387), .Y(n43569)
         );
  NOR4XL U34280 ( .A(n26767), .B(n26768), .C(n26770), .D(n26769), .Y(n44599)
         );
  NAND4X2 U34281 ( .A(n44470), .B(n44469), .C(n44468), .D(n44467), .Y(n44598)
         );
  NOR4XL U34282 ( .A(n26759), .B(n26760), .C(n26762), .D(n26761), .Y(n44601)
         );
  NOR4XL U34283 ( .A(n29173), .B(n29170), .C(n29171), .D(n29172), .Y(n44591)
         );
  NOR2XL U34284 ( .A(net171313), .B(n48227), .Y(n48228) );
  NAND3XL U34285 ( .A(n48336), .B(n48335), .C(n48334), .Y(n48340) );
  INVX1 U34286 ( .A(n29174), .Y(n43600) );
  CLKBUFX2 U34287 ( .A(n42513), .Y(n42512) );
  CLKBUFX2 U34288 ( .A(n42457), .Y(n42456) );
  NAND4X2 U34289 ( .A(n43240), .B(n43239), .C(n43238), .D(n43237), .Y(n11669)
         );
  OAI21X4 U34290 ( .A0(n47787), .A1(n47786), .B0(n47785), .Y(n47788) );
  NAND4X2 U34291 ( .A(n43249), .B(n43248), .C(n43247), .D(n43246), .Y(n12482)
         );
  CLKBUFX2 U34292 ( .A(n42480), .Y(n42478) );
  OAI211XL U34293 ( .A0(n9896), .A1(n9876), .B0(n49518), .C0(n9875), .Y(n9895)
         );
  NOR2XL U34294 ( .A(net171210), .B(net171205), .Y(n12018) );
  NAND2XL U34295 ( .A(n40188), .B(n37195), .Y(n49481) );
  NAND2XL U34296 ( .A(n40272), .B(n37554), .Y(n48564) );
  NOR4X1 U34297 ( .A(n10240), .B(n10242), .C(n10235), .D(net171458), .Y(n9798)
         );
  OR4XL U34298 ( .A(n10829), .B(net171453), .C(net171456), .D(net151662), .Y(
        n10235) );
  CLKINVX2 U34299 ( .A(n19180), .Y(n50142) );
  CLKBUFX2 U34300 ( .A(net151225), .Y(net221992) );
  NAND4BBXL U34301 ( .AN(n9840), .BN(n9838), .C(n49521), .D(n30441), .Y(n9763)
         );
  NOR3BXL U34302 ( .AN(n10837), .B(net171447), .C(n10839), .Y(n10244) );
  NOR3BX1 U34303 ( .AN(n10251), .B(n10254), .C(n10253), .Y(n9799) );
  NOR3BXL U34304 ( .AN(n9961), .B(n9963), .C(n9964), .Y(n9845) );
  NAND3BXL U34305 ( .AN(n47823), .B(n36936), .C(n47708), .Y(n47843) );
  NOR4XL U34306 ( .A(net171108), .B(net171327), .C(n10147), .D(n10148), .Y(
        n10144) );
  INVXL U34307 ( .A(net210476), .Y(net213675) );
  NOR2XL U34308 ( .A(net210479), .B(net210475), .Y(n45528) );
  NAND3BXL U34309 ( .AN(net210469), .B(n37126), .C(net209603), .Y(n47815) );
  NOR2XL U34310 ( .A(net209582), .B(net209592), .Y(n45527) );
  NAND4BX1 U34311 ( .AN(n10166), .B(n10196), .C(n28095), .D(net168843), .Y(
        n9787) );
  NOR2XL U34312 ( .A(net171214), .B(net171218), .Y(n28095) );
  NAND3BX1 U34313 ( .AN(n10177), .B(n10174), .C(net168842), .Y(n9788) );
  NOR3X1 U34314 ( .A(n9679), .B(n50145), .C(n19523), .Y(n19449) );
  NOR2X1 U34315 ( .A(n9737), .B(n50146), .Y(n19412) );
  CLKINVX1 U34316 ( .A(n37525), .Y(n42734) );
  INVXL U34317 ( .A(n11989), .Y(net209763) );
  INVXL U34318 ( .A(n11968), .Y(net209749) );
  INVXL U34319 ( .A(net260247), .Y(net209739) );
  OAI21X1 U34320 ( .A0(net209784), .A1(n48245), .B0(n12686), .Y(n48246) );
  OAI21X2 U34321 ( .A0(net209769), .A1(n48255), .B0(n12668), .Y(n48256) );
  INVXL U34322 ( .A(n12671), .Y(net209769) );
  INVXL U34323 ( .A(n10519), .Y(net209772) );
  INVXL U34324 ( .A(n12675), .Y(net209773) );
  AOI21XL U34325 ( .A0(n48136), .A1(n39304), .B0(net171234), .Y(n48200) );
  NAND4XL U34326 ( .A(n48167), .B(n48171), .C(net209884), .D(n48175), .Y(
        n48168) );
  AOI21XL U34327 ( .A0(n48141), .A1(net209893), .B0(net209926), .Y(n48170) );
  NAND2BX2 U34328 ( .AN(n48215), .B(n48214), .Y(n48216) );
  AOI21X2 U34329 ( .A0(n48129), .A1(n12795), .B0(n48128), .Y(n48218) );
  OAI21X2 U34330 ( .A0(n48211), .A1(n48210), .B0(n48209), .Y(n48217) );
  NOR2X4 U34331 ( .A(n43620), .B(n43619), .Y(n43621) );
  XNOR2XL U34332 ( .A(n51001), .B(n42542), .Y(n27468) );
  XNOR2XL U34333 ( .A(n42508), .B(n42058), .Y(n44038) );
  AND3X2 U34334 ( .A(n43594), .B(n43593), .C(n43592), .Y(n41682) );
  NAND4BX2 U34335 ( .AN(n41684), .B(n44028), .C(n44027), .D(n44026), .Y(n48336) );
  OR2X4 U34336 ( .A(n43603), .B(n43602), .Y(n41687) );
  NOR2X4 U34337 ( .A(n44288), .B(n44287), .Y(n44302) );
  NOR2X4 U34338 ( .A(n44299), .B(n44298), .Y(n44300) );
  INVXL U34339 ( .A(n10991), .Y(net209145) );
  INVXL U34340 ( .A(n11092), .Y(net209367) );
  AOI21XL U34341 ( .A0(n12274), .A1(net151458), .B0(net171461), .Y(n48528) );
  OAI21X2 U34342 ( .A0(n48526), .A1(n48525), .B0(n48524), .Y(n48527) );
  XNOR2XL U34343 ( .A(n50774), .B(net258207), .Y(n29172) );
  NAND4X4 U34344 ( .A(n44152), .B(n44151), .C(n44150), .D(n44149), .Y(n48319)
         );
  XNOR2XL U34345 ( .A(n51415), .B(n42693), .Y(n29176) );
  XNOR2XL U34346 ( .A(n36721), .B(n41802), .Y(n47550) );
  XNOR2XL U34347 ( .A(n50560), .B(n34435), .Y(n29175) );
  XNOR2XL U34348 ( .A(n50759), .B(net219434), .Y(n26765) );
  XNOR2XL U34349 ( .A(n50773), .B(net258207), .Y(n29142) );
  XNOR2XL U34350 ( .A(n50758), .B(n36865), .Y(n26757) );
  XNOR2XL U34351 ( .A(n51186), .B(n42631), .Y(n26756) );
  XOR2XL U34352 ( .A(n42068), .B(n36882), .Y(n44959) );
  AOI21XL U34353 ( .A0(n48460), .A1(net209287), .B0(net209288), .Y(n48463) );
  OAI2BB1XL U34354 ( .A0N(n12287), .A1N(n41695), .B0(n10827), .Y(n48520) );
  NOR4X2 U34355 ( .A(n43870), .B(n43869), .C(n43868), .D(n43867), .Y(n43871)
         );
  XNOR2XL U34356 ( .A(n50572), .B(n42724), .Y(n27521) );
  XNOR2XL U34357 ( .A(n51427), .B(n42697), .Y(n27522) );
  XOR2XL U34358 ( .A(n42087), .B(n36885), .Y(n44655) );
  XOR2XL U34359 ( .A(n42075), .B(n36873), .Y(n45189) );
  XOR2XL U34360 ( .A(n41316), .B(n41815), .Y(n46511) );
  XOR2XL U34361 ( .A(n42101), .B(n42663), .Y(n27726) );
  NAND4BBX2 U34362 ( .AN(n43849), .BN(n41696), .C(n43848), .D(n43847), .Y(
        n45530) );
  OR4X2 U34363 ( .A(n27726), .B(n27725), .C(n27724), .D(n27723), .Y(n41696) );
  XOR2XL U34364 ( .A(n42100), .B(n36880), .Y(n27734) );
  XOR2XL U34365 ( .A(n41852), .B(n36899), .Y(n27609) );
  XOR2XL U34366 ( .A(n41851), .B(n36898), .Y(n27579) );
  XOR2XL U34367 ( .A(n41848), .B(n36895), .Y(n27429) );
  XOR2XL U34368 ( .A(n41853), .B(n36894), .Y(n27519) );
  XOR2XL U34369 ( .A(n41851), .B(n42609), .Y(n27481) );
  XOR2XL U34370 ( .A(n42110), .B(n42663), .Y(n27485) );
  XOR2XL U34371 ( .A(n41843), .B(n42609), .Y(n27692) );
  XOR2XL U34372 ( .A(n42102), .B(n42663), .Y(n27696) );
  XOR2XL U34373 ( .A(n41853), .B(n42609), .Y(n27601) );
  XOR2XL U34374 ( .A(n42103), .B(n42663), .Y(n27996) );
  XOR2XL U34375 ( .A(n41844), .B(n42609), .Y(n27992) );
  XOR2XL U34376 ( .A(n42113), .B(n42663), .Y(n27515) );
  XOR2XL U34377 ( .A(n42110), .B(n36888), .Y(n27583) );
  XOR2XL U34378 ( .A(n42107), .B(n36882), .Y(n27433) );
  XOR2XL U34379 ( .A(n42112), .B(n36888), .Y(n27523) );
  XOR2XL U34380 ( .A(n41856), .B(n42526), .Y(n27531) );
  XNOR2XL U34381 ( .A(n51403), .B(n42698), .Y(n29055) );
  XNOR2XL U34382 ( .A(n51367), .B(n42698), .Y(n28184) );
  XNOR2XL U34383 ( .A(n51417), .B(n42693), .Y(n29236) );
  XNOR2XL U34384 ( .A(n51410), .B(n42693), .Y(n29296) );
  XOR2XL U34385 ( .A(n41824), .B(n36899), .Y(n44804) );
  XOR2XL U34386 ( .A(n42084), .B(n42659), .Y(n44800) );
  XOR2XL U34387 ( .A(n41815), .B(n36893), .Y(n45426) );
  XOR2XL U34388 ( .A(n42075), .B(n42660), .Y(n45422) );
  XOR2XL U34389 ( .A(n41814), .B(n36897), .Y(n45177) );
  XOR2XL U34390 ( .A(n41815), .B(n42595), .Y(n45169) );
  XOR2XL U34391 ( .A(n42074), .B(n42660), .Y(n45173) );
  XOR2XL U34392 ( .A(n41826), .B(n36891), .Y(n44835) );
  XOR2XL U34393 ( .A(n42086), .B(n42659), .Y(n44831) );
  XOR2XL U34394 ( .A(n41816), .B(n36892), .Y(n45446) );
  XOR2XL U34395 ( .A(n41820), .B(n36892), .Y(n45356) );
  XOR2XL U34396 ( .A(n42076), .B(n42660), .Y(n45442) );
  XOR2XL U34397 ( .A(n42080), .B(n42660), .Y(n45352) );
  XOR2XL U34398 ( .A(n42081), .B(n42660), .Y(n45294) );
  XOR2XL U34399 ( .A(n41819), .B(n36895), .Y(n45387) );
  XOR2XL U34400 ( .A(n41817), .B(n36899), .Y(n45475) );
  XOR2XL U34401 ( .A(n42079), .B(n42660), .Y(n45383) );
  XOR2XL U34402 ( .A(n42077), .B(n42660), .Y(n45471) );
  XOR2XL U34403 ( .A(n41823), .B(n36898), .Y(n44862) );
  XOR2XL U34404 ( .A(n41822), .B(n36900), .Y(n45329) );
  XOR2XL U34405 ( .A(n42083), .B(n42659), .Y(n44858) );
  XOR2XL U34406 ( .A(n42082), .B(n42660), .Y(n45325) );
  XOR2XL U34407 ( .A(n41838), .B(n36901), .Y(n44019) );
  XOR2XL U34408 ( .A(n41834), .B(n36894), .Y(n44049) );
  XOR2XL U34409 ( .A(n42094), .B(n42658), .Y(n44045) );
  XOR2XL U34410 ( .A(n41833), .B(n42604), .Y(n44103) );
  XOR2XL U34411 ( .A(n42092), .B(n42658), .Y(n44107) );
  XOR2XL U34412 ( .A(n42095), .B(n42658), .Y(n43922) );
  XOR2XL U34413 ( .A(n42088), .B(n36888), .Y(n44746) );
  XOR2XL U34414 ( .A(n41829), .B(n36891), .Y(n44742) );
  XOR2XL U34415 ( .A(n42089), .B(n42659), .Y(n44738) );
  XOR2XL U34416 ( .A(n41836), .B(n36898), .Y(n43957) );
  XOR2XL U34417 ( .A(n41837), .B(n42605), .Y(n43949) );
  XOR2XL U34418 ( .A(n42096), .B(n42658), .Y(n43953) );
  XOR2XL U34419 ( .A(n41830), .B(n42607), .Y(n44734) );
  XOR2XL U34420 ( .A(n41839), .B(n36894), .Y(n43895) );
  XOR2XL U34421 ( .A(n42093), .B(n42658), .Y(n44076) );
  XOR2XL U34422 ( .A(n41834), .B(n42605), .Y(n44072) );
  XOR2XL U34423 ( .A(n41825), .B(n36893), .Y(n44773) );
  XOR2XL U34424 ( .A(n41830), .B(n36897), .Y(n44713) );
  XOR2XL U34425 ( .A(n41831), .B(n42605), .Y(n44705) );
  XOR2XL U34426 ( .A(n42090), .B(n42658), .Y(n44709) );
  XOR2XL U34427 ( .A(n42085), .B(n42659), .Y(n44769) );
  XOR2XL U34428 ( .A(n41826), .B(n42605), .Y(n44765) );
  XOR2XL U34429 ( .A(n41802), .B(n42630), .Y(n43889) );
  XOR2XL U34430 ( .A(n42113), .B(n36881), .Y(n27553) );
  XOR2XL U34431 ( .A(n42117), .B(n36885), .Y(n27192) );
  XOR2XL U34432 ( .A(n41858), .B(n36897), .Y(n27188) );
  XOR2XL U34433 ( .A(n41900), .B(n36893), .Y(n25023) );
  XOR2XL U34434 ( .A(n41901), .B(n42608), .Y(n25015) );
  XOR2XL U34435 ( .A(n42160), .B(n42663), .Y(n25019) );
  XOR2XL U34436 ( .A(n42115), .B(n36886), .Y(n27252) );
  XOR2XL U34437 ( .A(n42145), .B(n36886), .Y(n26680) );
  XOR2XL U34438 ( .A(n41856), .B(n36901), .Y(n27248) );
  XOR2XL U34439 ( .A(n42116), .B(n36879), .Y(n27162) );
  XOR2XL U34440 ( .A(n42104), .B(n42662), .Y(n28026) );
  XOR2XL U34441 ( .A(n41845), .B(n42608), .Y(n28022) );
  XOR2XL U34442 ( .A(n42116), .B(n42662), .Y(n27244) );
  XOR2XL U34443 ( .A(n41857), .B(n42608), .Y(n27240) );
  XOR2XL U34444 ( .A(n41857), .B(n36891), .Y(n27158) );
  XOR2XL U34445 ( .A(n42117), .B(n42662), .Y(n27154) );
  XOR2XL U34446 ( .A(n41858), .B(n42608), .Y(n27150) );
  XOR2XL U34447 ( .A(n42160), .B(n36885), .Y(n25207) );
  XOR2XL U34448 ( .A(n41901), .B(n36892), .Y(n25203) );
  XOR2XL U34449 ( .A(n41888), .B(n36898), .Y(n26947) );
  XOR2XL U34450 ( .A(n42137), .B(n42652), .Y(n29048) );
  XOR2XL U34451 ( .A(n42119), .B(n36881), .Y(n27312) );
  XOR2XL U34452 ( .A(n41877), .B(n36898), .Y(n29052) );
  XOR2XL U34453 ( .A(n41904), .B(n36900), .Y(n24903) );
  XOR2XL U34454 ( .A(n42163), .B(n36880), .Y(n24907) );
  XOR2XL U34455 ( .A(n42102), .B(n36883), .Y(n28004) );
  XOR2XL U34456 ( .A(n42151), .B(n36885), .Y(n27131) );
  XOR2XL U34457 ( .A(n42136), .B(n36887), .Y(n29056) );
  XOR2XL U34458 ( .A(n41860), .B(n36891), .Y(n27308) );
  XOR2XL U34459 ( .A(n41905), .B(n42608), .Y(n24895) );
  XOR2XL U34460 ( .A(n42164), .B(n42665), .Y(n24899) );
  XOR2XL U34461 ( .A(n41902), .B(n42607), .Y(n25195) );
  XOR2XL U34462 ( .A(n41892), .B(n36893), .Y(n27127) );
  XOR2XL U34463 ( .A(n42120), .B(n42662), .Y(n27304) );
  XOR2XL U34464 ( .A(n41861), .B(n42608), .Y(n27300) );
  XOR2XL U34465 ( .A(n42162), .B(n36883), .Y(n24877) );
  XOR2XL U34466 ( .A(n42152), .B(n36888), .Y(n27041) );
  XOR2XL U34467 ( .A(n42148), .B(n36889), .Y(n26981) );
  XOR2XL U34468 ( .A(n41903), .B(n36891), .Y(n24873) );
  XOR2XL U34469 ( .A(n41893), .B(n42607), .Y(n27119) );
  XOR2XL U34470 ( .A(n42152), .B(n42661), .Y(n27123) );
  XOR2XL U34471 ( .A(n42143), .B(n36886), .Y(n26890) );
  XOR2XL U34472 ( .A(n41893), .B(n36900), .Y(n27037) );
  XOR2XL U34473 ( .A(n42114), .B(n36883), .Y(n27282) );
  XOR2XL U34474 ( .A(n42149), .B(n36888), .Y(n27011) );
  XOR2XL U34475 ( .A(n42146), .B(n36889), .Y(n26921) );
  XOR2XL U34476 ( .A(n42118), .B(n36881), .Y(n27222) );
  XOR2XL U34477 ( .A(n41889), .B(n36895), .Y(n26977) );
  XOR2XL U34478 ( .A(n41894), .B(n42608), .Y(n27029) );
  XOR2XL U34479 ( .A(n42153), .B(n42662), .Y(n27033) );
  XOR2XL U34480 ( .A(n42163), .B(n42661), .Y(n24869) );
  XOR2XL U34481 ( .A(n42149), .B(n42661), .Y(n26973) );
  XOR2XL U34482 ( .A(n41890), .B(n36891), .Y(n27007) );
  XOR2XL U34483 ( .A(n41855), .B(n36895), .Y(n27278) );
  XOR2XL U34484 ( .A(n41870), .B(n36899), .Y(n29293) );
  XOR2XL U34485 ( .A(n41890), .B(n42607), .Y(n26969) );
  XOR2XL U34486 ( .A(n41904), .B(n42608), .Y(n24865) );
  XOR2XL U34487 ( .A(n41871), .B(n42602), .Y(n29285) );
  XOR2XL U34488 ( .A(n41859), .B(n36899), .Y(n27218) );
  XOR2XL U34489 ( .A(n41887), .B(n36893), .Y(n26917) );
  XOR2XL U34490 ( .A(n42121), .B(n36881), .Y(n27342) );
  XOR2XL U34491 ( .A(n42129), .B(n36888), .Y(n29297) );
  XOR2XL U34492 ( .A(n41874), .B(n36900), .Y(n29443) );
  XOR2XL U34493 ( .A(n42134), .B(n42653), .Y(n29439) );
  XOR2XL U34494 ( .A(n41875), .B(n42602), .Y(n29435) );
  XOR2XL U34495 ( .A(n42150), .B(n42661), .Y(n27003) );
  XOR2XL U34496 ( .A(n41891), .B(n42607), .Y(n26999) );
  XOR2XL U34497 ( .A(n42165), .B(n36887), .Y(n24967) );
  XOR2XL U34498 ( .A(n41906), .B(n36898), .Y(n24963) );
  XOR2XL U34499 ( .A(n41862), .B(n36892), .Y(n27338) );
  XOR2XL U34500 ( .A(n42119), .B(n42662), .Y(n27214) );
  XOR2XL U34501 ( .A(n41860), .B(n42608), .Y(n27210) );
  XOR2XL U34502 ( .A(n42115), .B(n42662), .Y(n27274) );
  XOR2XL U34503 ( .A(n42133), .B(n36880), .Y(n29447) );
  XOR2XL U34504 ( .A(n42147), .B(n42661), .Y(n26913) );
  XOR2XL U34505 ( .A(n41856), .B(n42608), .Y(n27270) );
  XOR2XL U34506 ( .A(n41888), .B(n42607), .Y(n26909) );
  XOR2XL U34507 ( .A(n42166), .B(n42665), .Y(n24959) );
  XOR2XL U34508 ( .A(n41922), .B(n36897), .Y(n28301) );
  XOR2XL U34509 ( .A(n42181), .B(n36888), .Y(n28305) );
  XOR2XL U34510 ( .A(n41913), .B(n36899), .Y(n28181) );
  XOR2XL U34511 ( .A(n41845), .B(n36891), .Y(n28090) );
  XOR2XL U34512 ( .A(n42172), .B(n36886), .Y(n28185) );
  XOR2XL U34513 ( .A(n42182), .B(n41286), .Y(n28297) );
  XOR2XL U34514 ( .A(n41914), .B(n42600), .Y(n28173) );
  XOR2XL U34515 ( .A(n42173), .B(n41286), .Y(n28177) );
  XOR2XL U34516 ( .A(n41846), .B(n42600), .Y(n28082) );
  XOR2XL U34517 ( .A(n42105), .B(n41286), .Y(n28086) );
  XOR2XL U34518 ( .A(n41805), .B(n42615), .Y(n43888) );
  XOR2XL U34519 ( .A(n42158), .B(n36873), .Y(n25126) );
  XNOR2XL U34520 ( .A(n51002), .B(n42618), .Y(n27478) );
  XNOR2XL U34521 ( .A(n51010), .B(n42618), .Y(n27689) );
  XNOR2XL U34522 ( .A(n50366), .B(n42675), .Y(n27542) );
  XNOR2XL U34523 ( .A(n50999), .B(net219310), .Y(n27546) );
  XNOR2XL U34524 ( .A(n51000), .B(n42618), .Y(n27598) );
  XNOR2XL U34525 ( .A(n50370), .B(n42675), .Y(n27482) );
  XNOR2XL U34526 ( .A(n51003), .B(net219314), .Y(n27486) );
  XNOR2XL U34527 ( .A(n50378), .B(n42675), .Y(n27693) );
  XNOR2XL U34528 ( .A(n49514), .B(net219314), .Y(n27697) );
  XNOR2XL U34529 ( .A(n50368), .B(n42675), .Y(n27602) );
  XNOR2XL U34530 ( .A(n51001), .B(n40039), .Y(n27606) );
  XNOR2XL U34531 ( .A(n50950), .B(n42613), .Y(n25162) );
  XNOR2XL U34532 ( .A(n50320), .B(n42672), .Y(n25016) );
  XNOR2XL U34533 ( .A(n50953), .B(net219330), .Y(n25020) );
  XNOR2XL U34534 ( .A(n50995), .B(n42615), .Y(n27147) );
  XNOR2XL U34535 ( .A(n50318), .B(n42674), .Y(n25166) );
  XNOR2XL U34536 ( .A(n50951), .B(net219310), .Y(n25170) );
  XNOR2XL U34537 ( .A(n51001), .B(n42618), .Y(n27568) );
  XNOR2XL U34538 ( .A(n50964), .B(n42615), .Y(n26936) );
  XNOR2XL U34539 ( .A(n50363), .B(n42674), .Y(n27151) );
  XNOR2XL U34540 ( .A(n50951), .B(n42613), .Y(n25192) );
  XNOR2XL U34541 ( .A(n50948), .B(n36868), .Y(n24892) );
  XNOR2XL U34542 ( .A(n50996), .B(n40039), .Y(n27155) );
  XNOR2XL U34543 ( .A(n50960), .B(n42615), .Y(n27116) );
  XOR2XL U34544 ( .A(n42063), .B(n42558), .Y(n44035) );
  XNOR2XL U34545 ( .A(n50561), .B(n42717), .Y(n29205) );
  XNOR2XL U34546 ( .A(n50557), .B(n36709), .Y(n29355) );
  XNOR2XL U34547 ( .A(n50558), .B(n42717), .Y(n29325) );
  XNOR2XL U34548 ( .A(n50562), .B(n42723), .Y(n29235) );
  XNOR2XL U34549 ( .A(n50549), .B(n42717), .Y(n29114) );
  XNOR2XL U34550 ( .A(n50789), .B(net219466), .Y(n27488) );
  XNOR2XL U34551 ( .A(n50739), .B(net219434), .Y(n25022) );
  XNOR2XL U34552 ( .A(n49513), .B(net219466), .Y(n27699) );
  XNOR2XL U34553 ( .A(n50787), .B(net219466), .Y(n27608) );
  XNOR2XL U34554 ( .A(n50788), .B(n42592), .Y(n27480) );
  XNOR2XL U34555 ( .A(n50737), .B(net219434), .Y(n25172) );
  XNOR2XL U34556 ( .A(n50796), .B(n42592), .Y(n27691) );
  XNOR2XL U34557 ( .A(n50738), .B(n36863), .Y(n25014) );
  XNOR2XL U34558 ( .A(n51429), .B(n42642), .Y(n27484) );
  XNOR2XL U34559 ( .A(n50782), .B(net219468), .Y(n27157) );
  XNOR2XL U34560 ( .A(n51437), .B(n42642), .Y(n27695) );
  XNOR2XL U34561 ( .A(n50738), .B(net219434), .Y(n25202) );
  XNOR2XL U34562 ( .A(n50751), .B(net219434), .Y(n26946) );
  XNOR2XL U34563 ( .A(n51379), .B(n36861), .Y(n25018) );
  XNOR2XL U34564 ( .A(n51427), .B(n42642), .Y(n27604) );
  XNOR2XL U34565 ( .A(n50788), .B(net219466), .Y(n27578) );
  XNOR2XL U34566 ( .A(n50735), .B(net219434), .Y(n24902) );
  XNOR2XL U34567 ( .A(n50736), .B(n36865), .Y(n25164) );
  XNOR2XL U34568 ( .A(n50792), .B(n42592), .Y(n28051) );
  XNOR2XL U34569 ( .A(n50747), .B(net219434), .Y(n27126) );
  XNOR2XL U34570 ( .A(n50779), .B(net219466), .Y(n27307) );
  XNOR2XL U34571 ( .A(n50736), .B(net219434), .Y(n24872) );
  XNOR2XL U34572 ( .A(n50796), .B(net219468), .Y(n27999) );
  XNOR2XL U34573 ( .A(n50781), .B(n36863), .Y(n27149) );
  XNOR2XL U34574 ( .A(n50746), .B(net219434), .Y(n27036) );
  XNOR2XL U34575 ( .A(n51377), .B(n36861), .Y(n25168) );
  XNOR2XL U34576 ( .A(n50750), .B(net219434), .Y(n26976) );
  XNOR2XL U34577 ( .A(n50755), .B(net219434), .Y(n26885) );
  XNOR2XL U34578 ( .A(n50786), .B(net219466), .Y(n27518) );
  XNOR2XL U34579 ( .A(n50784), .B(net219442), .Y(n27277) );
  XNOR2XL U34580 ( .A(n50749), .B(net219442), .Y(n27006) );
  XNOR2XL U34581 ( .A(n50752), .B(net219442), .Y(n26916) );
  XNOR2XL U34582 ( .A(n50780), .B(net219468), .Y(n27217) );
  XNOR2XL U34583 ( .A(n51415), .B(n42642), .Y(n29198) );
  XNOR2XL U34584 ( .A(n51411), .B(n42643), .Y(n29348) );
  XNOR2XL U34585 ( .A(n51216), .B(n42633), .Y(n27479) );
  XNOR2XL U34586 ( .A(n51224), .B(n42627), .Y(n27690) );
  XNOR2XL U34587 ( .A(n51214), .B(n42631), .Y(n27599) );
  XNOR2XL U34588 ( .A(n51166), .B(n34447), .Y(n25013) );
  XNOR2XL U34589 ( .A(n50574), .B(n36903), .Y(n27483) );
  XNOR2XL U34590 ( .A(n51217), .B(n41281), .Y(n27487) );
  XNOR2XL U34591 ( .A(n50582), .B(n36903), .Y(n27694) );
  XNOR2XL U34592 ( .A(n49516), .B(n41282), .Y(n27698) );
  XNOR2XL U34593 ( .A(n50572), .B(n36903), .Y(n27603) );
  XNOR2XL U34594 ( .A(n51215), .B(n41283), .Y(n27607) );
  XNOR2XL U34595 ( .A(n51164), .B(n42629), .Y(n25163) );
  XNOR2XL U34596 ( .A(n50524), .B(n41319), .Y(n25017) );
  XNOR2XL U34597 ( .A(n51167), .B(n41283), .Y(n25021) );
  XNOR2XL U34598 ( .A(n50581), .B(n42724), .Y(n28032) );
  XNOR2XL U34599 ( .A(n51220), .B(n42632), .Y(n28050) );
  XNOR2XL U34600 ( .A(n51209), .B(n42628), .Y(n27148) );
  XNOR2XL U34601 ( .A(n50522), .B(n36905), .Y(n25167) );
  XNOR2XL U34602 ( .A(n51165), .B(n41281), .Y(n25171) );
  XNOR2XL U34603 ( .A(n51215), .B(n42629), .Y(n27569) );
  XNOR2XL U34604 ( .A(n51178), .B(n42633), .Y(n26937) );
  XNOR2XL U34605 ( .A(n50567), .B(n36834), .Y(n27152) );
  XNOR2XL U34606 ( .A(n51165), .B(n42633), .Y(n25193) );
  XNOR2XL U34607 ( .A(n51183), .B(n42624), .Y(n26846) );
  XNOR2XL U34608 ( .A(n51162), .B(n34447), .Y(n24893) );
  XNOR2XL U34609 ( .A(n51210), .B(n41283), .Y(n27156) );
  XNOR2XL U34610 ( .A(n51174), .B(n42629), .Y(n27117) );
  XNOR2XL U34611 ( .A(n51223), .B(n42632), .Y(n27990) );
  XNOR2XL U34612 ( .A(n51202), .B(n42627), .Y(n29193) );
  XNOR2XL U34613 ( .A(n51198), .B(n42633), .Y(n29343) );
  XNOR2XL U34614 ( .A(n50976), .B(n40039), .Y(n29049) );
  XNOR2XL U34615 ( .A(n50762), .B(net219468), .Y(n29051) );
  XNOR2XL U34616 ( .A(n50364), .B(n42710), .Y(n27159) );
  XNOR2XL U34617 ( .A(n50568), .B(n42723), .Y(n27160) );
  XNOR2XL U34618 ( .A(n51423), .B(n42697), .Y(n27161) );
  XNOR2XL U34619 ( .A(n50332), .B(n42710), .Y(n26978) );
  XNOR2XL U34620 ( .A(n50536), .B(n42723), .Y(n26979) );
  XNOR2XL U34621 ( .A(n51391), .B(n42697), .Y(n26980) );
  XOR2XL U34622 ( .A(n42074), .B(n36873), .Y(n45220) );
  XOR2XL U34623 ( .A(n42071), .B(n36873), .Y(n44987) );
  XOR2XL U34624 ( .A(n41899), .B(n42531), .Y(n25125) );
  XOR2XL U34625 ( .A(n42085), .B(n41321), .Y(n44818) );
  XOR2XL U34626 ( .A(n42095), .B(n36877), .Y(n44063) );
  XOR2XL U34627 ( .A(n42093), .B(n41321), .Y(n44125) );
  XOR2XL U34628 ( .A(n42088), .B(n36877), .Y(n44696) );
  XOR2XL U34629 ( .A(n42087), .B(n36801), .Y(n44845) );
  XOR2XL U34630 ( .A(n42077), .B(n36877), .Y(n45458) );
  XOR2XL U34631 ( .A(n42097), .B(n36873), .Y(n43971) );
  XOR2XL U34632 ( .A(n42089), .B(n36877), .Y(n44665) );
  XOR2XL U34633 ( .A(n42094), .B(n36873), .Y(n44094) );
  XOR2XL U34634 ( .A(n42082), .B(n36877), .Y(n45312) );
  XOR2XL U34635 ( .A(n42115), .B(n36801), .Y(n27532) );
  XNOR2XL U34636 ( .A(n51383), .B(n42700), .Y(n25146) );
  XOR2XL U34637 ( .A(n42156), .B(n36881), .Y(n25147) );
  XOR2XL U34638 ( .A(n41897), .B(n36897), .Y(n25143) );
  XOR2XL U34639 ( .A(n41898), .B(n42612), .Y(n25135) );
  XOR2XL U34640 ( .A(n41841), .B(n36892), .Y(n27730) );
  XNOR2XL U34641 ( .A(n51429), .B(n42697), .Y(n27582) );
  XNOR2XL U34642 ( .A(n50320), .B(n42707), .Y(n25204) );
  XNOR2XL U34643 ( .A(n51379), .B(n42691), .Y(n25206) );
  XNOR2XL U34644 ( .A(n50378), .B(n42712), .Y(n28001) );
  XNOR2XL U34645 ( .A(n50582), .B(n36709), .Y(n28002) );
  XNOR2XL U34646 ( .A(n51437), .B(n42697), .Y(n28003) );
  XNOR2XL U34647 ( .A(n50366), .B(n42710), .Y(n27279) );
  XNOR2XL U34648 ( .A(n50570), .B(n42723), .Y(n27280) );
  XNOR2XL U34649 ( .A(n51425), .B(n42697), .Y(n27281) );
  XNOR2XL U34650 ( .A(n50334), .B(n41642), .Y(n26918) );
  XNOR2XL U34651 ( .A(n50538), .B(n36875), .Y(n26919) );
  XNOR2XL U34652 ( .A(n51393), .B(n42697), .Y(n26920) );
  XNOR2XL U34653 ( .A(n50742), .B(net219434), .Y(n25142) );
  XNOR2XL U34654 ( .A(n50955), .B(n36868), .Y(n25132) );
  XNOR2XL U34655 ( .A(n50323), .B(n36907), .Y(n25136) );
  XNOR2XL U34656 ( .A(n50324), .B(n42707), .Y(n25144) );
  XNOR2XL U34657 ( .A(n50741), .B(n36865), .Y(n25134) );
  XNOR2XL U34658 ( .A(n50956), .B(net219310), .Y(n25140) );
  XNOR2XL U34659 ( .A(n50528), .B(n42717), .Y(n25145) );
  XNOR2XL U34660 ( .A(n51169), .B(n42627), .Y(n25133) );
  XNOR2XL U34661 ( .A(n50527), .B(n36903), .Y(n25137) );
  XNOR2XL U34662 ( .A(n51170), .B(n41281), .Y(n25141) );
  XOR2XL U34663 ( .A(n41321), .B(n42099), .Y(n44032) );
  XOR2XL U34664 ( .A(n36809), .B(n42068), .Y(n46483) );
  XOR2XL U34665 ( .A(n36810), .B(n42069), .Y(n46474) );
  XNOR2XL U34666 ( .A(n36813), .B(n42067), .Y(n46581) );
  XNOR2XL U34667 ( .A(n41309), .B(n41809), .Y(n46577) );
  OAI211XL U34668 ( .A0(n48466), .A1(net209277), .B0(n48465), .C0(n48464), .Y(
        n48470) );
  NOR2X4 U34669 ( .A(n44842), .B(net209583), .Y(n44852) );
  XOR2XL U34670 ( .A(n41828), .B(n42522), .Y(n44842) );
  XOR2XL U34671 ( .A(n41830), .B(n42522), .Y(n44662) );
  XOR2XL U34672 ( .A(n41823), .B(n42523), .Y(n45309) );
  NOR2X4 U34673 ( .A(n44815), .B(net210650), .Y(n44825) );
  XOR2XL U34674 ( .A(n41832), .B(n42522), .Y(n44722) );
  XOR2XL U34675 ( .A(n41318), .B(n41841), .Y(n46210) );
  XOR2XL U34676 ( .A(n41311), .B(n41824), .Y(n46376) );
  XOR2XL U34677 ( .A(n41314), .B(n41820), .Y(n46332) );
  XOR2XL U34678 ( .A(n41309), .B(n41823), .Y(n46383) );
  XOR2XL U34679 ( .A(n41310), .B(n41819), .Y(n46321) );
  XOR2XL U34680 ( .A(n36754), .B(n34351), .Y(n47634) );
  XOR2XL U34681 ( .A(n36760), .B(n41815), .Y(n47590) );
  XOR2XL U34682 ( .A(n41836), .B(n42522), .Y(n44060) );
  XOR2XL U34683 ( .A(n36761), .B(n41839), .Y(n47532) );
  NAND2XL U34684 ( .A(n12389), .B(net209185), .Y(n48530) );
  XOR2XL U34685 ( .A(n36759), .B(n41829), .Y(n47380) );
  AOI21XL U34686 ( .A0(n47973), .A1(n11442), .B0(n47972), .Y(n48052) );
  NAND2XL U34687 ( .A(n10734), .B(n10732), .Y(n47972) );
  NAND2XL U34688 ( .A(n12922), .B(n10689), .Y(n47961) );
  INVXL U34689 ( .A(n11365), .Y(n47960) );
  XOR2XL U34690 ( .A(n36761), .B(n41835), .Y(n47490) );
  XOR2XL U34691 ( .A(n41829), .B(n42522), .Y(n44693) );
  XOR2XL U34692 ( .A(n41822), .B(n42523), .Y(n45367) );
  XOR2XL U34693 ( .A(n41835), .B(n42522), .Y(n44091) );
  XOR2XL U34694 ( .A(n41831), .B(n42522), .Y(n44753) );
  XOR2XL U34695 ( .A(n41838), .B(n42522), .Y(n43968) );
  XOR2XL U34696 ( .A(n41318), .B(n41839), .Y(n46271) );
  XOR2XL U34697 ( .A(n41833), .B(n42522), .Y(n44153) );
  XOR2XL U34698 ( .A(n36754), .B(n41837), .Y(n47521) );
  XOR2XL U34699 ( .A(n41318), .B(n41836), .Y(n46260) );
  OAI21X1 U34700 ( .A0(net171538), .A1(net210259), .B0(n12931), .Y(n47953) );
  XOR2XL U34701 ( .A(n36756), .B(n41830), .Y(n47391) );
  XOR2XL U34702 ( .A(n36753), .B(n41838), .Y(n47510) );
  XOR2XL U34703 ( .A(n36753), .B(n41825), .Y(n47424) );
  OAI21X1 U34704 ( .A0(net171443), .A1(n48414), .B0(n11095), .Y(n48415) );
  OAI21X2 U34705 ( .A0(n48533), .A1(n48532), .B0(n11040), .Y(n48534) );
  AOI21XL U34706 ( .A0(n48053), .A1(n12967), .B0(net151728), .Y(n48054) );
  XOR2XL U34707 ( .A(n36754), .B(n41823), .Y(n47369) );
  XOR2XL U34708 ( .A(n36756), .B(n41833), .Y(n47468) );
  XOR2XL U34709 ( .A(n36761), .B(n41831), .Y(n47402) );
  XOR2XL U34710 ( .A(n36757), .B(n41828), .Y(n47457) );
  XOR2XL U34711 ( .A(n41309), .B(n41835), .Y(n46249) );
  XOR2XL U34712 ( .A(n36760), .B(n41832), .Y(n47413) );
  XOR2XL U34713 ( .A(n41311), .B(n41828), .Y(n46434) );
  XOR2XL U34714 ( .A(n36753), .B(n41821), .Y(n47336) );
  XOR2XL U34715 ( .A(n36754), .B(n41834), .Y(n47479) );
  XOR2XL U34716 ( .A(n36756), .B(n41824), .Y(n47358) );
  XOR2XL U34717 ( .A(n36761), .B(n41819), .Y(n47314) );
  OAI21X2 U34718 ( .A0(n48454), .A1(n48453), .B0(n48452), .Y(n48458) );
  OAI21X1 U34719 ( .A0(net210251), .A1(n47956), .B0(n40394), .Y(n47958) );
  NOR2X2 U34720 ( .A(n29126), .B(n29143), .Y(n43610) );
  OAI2BB1X4 U34721 ( .A0N(n41702), .A1N(n41703), .B0(n12906), .Y(n48100) );
  XOR2XL U34722 ( .A(n36754), .B(n41812), .Y(n47601) );
  XOR2XL U34723 ( .A(n36755), .B(n41817), .Y(n47293) );
  XOR2XL U34724 ( .A(n36753), .B(n41827), .Y(n47446) );
  NOR2X2 U34725 ( .A(n25116), .B(n25117), .Y(n44457) );
  XOR2XL U34726 ( .A(n41819), .B(n42523), .Y(n45485) );
  XNOR2XL U34727 ( .A(n51382), .B(n36861), .Y(n25138) );
  CLKINVX3 U34728 ( .A(n29140), .Y(n43615) );
  NOR2X2 U34729 ( .A(n29124), .B(n29146), .Y(n43616) );
  NOR2X2 U34730 ( .A(n25092), .B(n25093), .Y(n44463) );
  AO21X2 U34731 ( .A0(n48202), .A1(n12749), .B0(net209844), .Y(n41783) );
  NAND2XL U34732 ( .A(n11399), .B(n11396), .Y(n48066) );
  AO21X4 U34733 ( .A0(n48224), .A1(net209814), .B0(n48223), .Y(n41779) );
  NAND3XL U34734 ( .A(n39304), .B(n48188), .C(n48187), .Y(n48189) );
  OAI2BB1X2 U34735 ( .A0N(n48201), .A1N(n12751), .B0(n12747), .Y(n48202) );
  NAND2XL U34736 ( .A(n48160), .B(net209893), .Y(n48161) );
  NAND2BXL U34737 ( .AN(net209301), .B(net209300), .Y(n48455) );
  NAND2X2 U34738 ( .A(n48116), .B(n10543), .Y(n48117) );
  OR4X2 U34739 ( .A(n44957), .B(n44956), .C(n44955), .D(n44954), .Y(n41707) );
  NAND2XL U34740 ( .A(net210148), .B(n48040), .Y(n48042) );
  NAND2XL U34741 ( .A(net209341), .B(net209300), .Y(n48433) );
  OAI21X2 U34742 ( .A0(net171240), .A1(n48204), .B0(n12793), .Y(n48205) );
  XOR2XL U34743 ( .A(n41820), .B(n42523), .Y(n45512) );
  CLKINVX3 U34744 ( .A(n10846), .Y(net209372) );
  XNOR2XL U34745 ( .A(n51200), .B(n42550), .Y(n29153) );
  XNOR2X1 U34746 ( .A(n42059), .B(n36875), .Y(n41713) );
  OA21X4 U34747 ( .A0(n12154), .A1(net171218), .B0(n12797), .Y(n41776) );
  XNOR2XL U34748 ( .A(n50973), .B(net219310), .Y(n26763) );
  XNOR2XL U34749 ( .A(n50355), .B(n42704), .Y(n29144) );
  XNOR2XL U34750 ( .A(n51201), .B(n42628), .Y(n29163) );
  XNOR2XL U34751 ( .A(n51399), .B(n36867), .Y(n26761) );
  XNOR2XL U34752 ( .A(n51413), .B(n42638), .Y(n29138) );
  XNOR2XL U34753 ( .A(n51202), .B(n41282), .Y(n29171) );
  XNOR2XL U34754 ( .A(n50986), .B(n41284), .Y(n29132) );
  XNOR2XL U34755 ( .A(n51414), .B(n36867), .Y(n29168) );
  XNOR2XL U34756 ( .A(n50336), .B(n42709), .Y(n26827) );
  XNOR2XL U34757 ( .A(n50540), .B(n34435), .Y(n26828) );
  XNOR2XL U34758 ( .A(n51395), .B(n42696), .Y(n26829) );
  XNOR2XL U34759 ( .A(n50515), .B(n41287), .Y(n24815) );
  XNOR2XL U34760 ( .A(n50360), .B(n42711), .Y(n27369) );
  XNOR2XL U34761 ( .A(n50564), .B(n42724), .Y(n27370) );
  XNOR2XL U34762 ( .A(n51419), .B(n42701), .Y(n27371) );
  XNOR2XL U34763 ( .A(n50330), .B(n42710), .Y(n27098) );
  XNOR2XL U34764 ( .A(n50534), .B(n42723), .Y(n27099) );
  XNOR2XL U34765 ( .A(n51389), .B(n42697), .Y(n27100) );
  XNOR2XL U34766 ( .A(n51191), .B(n41283), .Y(n29110) );
  XNOR2XL U34767 ( .A(n50763), .B(net219468), .Y(n29111) );
  XNOR2XL U34768 ( .A(n51153), .B(n41281), .Y(n28209) );
  XNOR2XL U34769 ( .A(n50725), .B(net219468), .Y(n28210) );
  XNOR2XL U34770 ( .A(n50941), .B(net219310), .Y(n28118) );
  XNOR2XL U34771 ( .A(n50727), .B(net219468), .Y(n28120) );
  XNOR2XL U34772 ( .A(n50982), .B(net219310), .Y(n29410) );
  XNOR2XL U34773 ( .A(n50937), .B(net219310), .Y(n28508) );
  XNOR2XL U34774 ( .A(n51151), .B(n41281), .Y(n28509) );
  XNOR2XL U34775 ( .A(n50723), .B(net219468), .Y(n28510) );
  XNOR2XL U34776 ( .A(n50935), .B(net219336), .Y(n28538) );
  XNOR2XL U34777 ( .A(n51149), .B(n41281), .Y(n28539) );
  XNOR2XL U34778 ( .A(n50721), .B(net219468), .Y(n28540) );
  XOR2XL U34779 ( .A(n41861), .B(n36894), .Y(n27368) );
  XOR2XL U34780 ( .A(n42120), .B(n36885), .Y(n27372) );
  XOR2XL U34781 ( .A(n41844), .B(n42526), .Y(n27682) );
  XOR2XL U34782 ( .A(n41853), .B(n42526), .Y(n27561) );
  XOR2XL U34783 ( .A(n41855), .B(n42526), .Y(n27501) );
  XOR2XL U34784 ( .A(n41845), .B(n42526), .Y(n27982) );
  XOR2XL U34785 ( .A(n41864), .B(n42526), .Y(n27320) );
  XOR2XL U34786 ( .A(n41849), .B(n42526), .Y(n27381) );
  XOR2XL U34787 ( .A(n41925), .B(n41312), .Y(n23186) );
  XOR2XL U34788 ( .A(n41842), .B(n36761), .Y(n20411) );
  XOR2XL U34789 ( .A(n41924), .B(n41316), .Y(n23146) );
  XOR2XL U34790 ( .A(n41921), .B(n41316), .Y(n23126) );
  XOR2XL U34791 ( .A(n41861), .B(n41311), .Y(n23716) );
  XOR2XL U34792 ( .A(n41860), .B(n41317), .Y(n23706) );
  XOR2XL U34793 ( .A(n41847), .B(n41318), .Y(n23847) );
  XOR2XL U34794 ( .A(n41905), .B(n41313), .Y(n23593) );
  XOR2XL U34795 ( .A(n41842), .B(n41310), .Y(n23787) );
  XOR2XL U34796 ( .A(n41846), .B(n41309), .Y(n23857) );
  XOR2XL U34797 ( .A(n41859), .B(n41310), .Y(n23736) );
  XOR2XL U34798 ( .A(n41853), .B(n41318), .Y(n23937) );
  XOR2XL U34799 ( .A(n41862), .B(n41318), .Y(n23766) );
  XOR2XL U34800 ( .A(n41858), .B(n41313), .Y(n23746) );
  XOR2XL U34801 ( .A(n41848), .B(n41310), .Y(n23837) );
  XOR2XL U34802 ( .A(n41849), .B(n41316), .Y(n23977) );
  XOR2XL U34803 ( .A(n41856), .B(n41311), .Y(n23987) );
  XOR2XL U34804 ( .A(n41851), .B(n41316), .Y(n23957) );
  XOR2XL U34805 ( .A(n41866), .B(n41314), .Y(n22459) );
  XOR2XL U34806 ( .A(n41863), .B(n41311), .Y(n23696) );
  XOR2XL U34807 ( .A(n41867), .B(n41317), .Y(n22449) );
  XOR2XL U34808 ( .A(n41872), .B(n41312), .Y(n22419) );
  XOR2XL U34809 ( .A(n41865), .B(n41311), .Y(n22469) );
  XOR2XL U34810 ( .A(n41893), .B(n41317), .Y(n24150) );
  XOR2XL U34811 ( .A(n41891), .B(n41316), .Y(n24109) );
  XOR2XL U34812 ( .A(n41888), .B(n41312), .Y(n24018) );
  XOR2XL U34813 ( .A(n41880), .B(n41311), .Y(n22319) );
  XOR2XL U34814 ( .A(n41896), .B(n41310), .Y(n24160) );
  XOR2XL U34815 ( .A(n41890), .B(n41313), .Y(n24119) );
  XOR2XL U34816 ( .A(n41873), .B(n41316), .Y(n22359) );
  XOR2XL U34817 ( .A(n41895), .B(n41311), .Y(n24139) );
  XOR2XL U34818 ( .A(n41883), .B(n41309), .Y(n24038) );
  XOR2XL U34819 ( .A(n41909), .B(n41309), .Y(n23471) );
  XOR2XL U34820 ( .A(n41884), .B(n41311), .Y(n24028) );
  XOR2XL U34821 ( .A(n41852), .B(n41318), .Y(n23947) );
  XOR2XL U34822 ( .A(n41874), .B(n41318), .Y(n22369) );
  XOR2XL U34823 ( .A(n41907), .B(n41313), .Y(n23571) );
  XOR2XL U34824 ( .A(n41864), .B(n41310), .Y(n23726) );
  XOR2XL U34825 ( .A(n41882), .B(n41318), .Y(n24048) );
  XOR2XL U34826 ( .A(n41881), .B(n41316), .Y(n24058) );
  XOR2XL U34827 ( .A(n41850), .B(n41316), .Y(n23967) );
  XOR2XL U34828 ( .A(n41870), .B(n36754), .Y(n19536) );
  XOR2XL U34829 ( .A(n41885), .B(n41317), .Y(n24078) );
  XOR2XL U34830 ( .A(n41906), .B(n41311), .Y(n23582) );
  XOR2XL U34831 ( .A(n41899), .B(n41318), .Y(n23531) );
  XOR2XL U34832 ( .A(n41904), .B(n41309), .Y(n23491) );
  XOR2XL U34833 ( .A(n41897), .B(n41311), .Y(n235510) );
  XOR2XL U34834 ( .A(n41877), .B(n41311), .Y(n22339) );
  XOR2XL U34835 ( .A(n41875), .B(n41311), .Y(n22379) );
  XOR2XL U34836 ( .A(n41846), .B(n36755), .Y(n20299) );
  XOR2XL U34837 ( .A(n41898), .B(n41317), .Y(n23541) );
  XOR2XL U34838 ( .A(n41894), .B(n41314), .Y(n24170) );
  XOR2XL U34839 ( .A(n41911), .B(n41317), .Y(n23451) );
  XOR2XL U34840 ( .A(n41876), .B(n41309), .Y(n22389) );
  XNOR2XL U34841 ( .A(n49516), .B(n36721), .Y(n20409) );
  XNOR2XL U34842 ( .A(n51143), .B(n41332), .Y(n23144) );
  XNOR2XL U34843 ( .A(n51146), .B(n41331), .Y(n23124) );
  XNOR2XL U34844 ( .A(n49513), .B(n42470), .Y(n20410) );
  XNOR2XL U34845 ( .A(n51435), .B(n42698), .Y(n28093) );
  XNOR2XL U34846 ( .A(n51366), .B(n42698), .Y(n28214) );
  XNOR2XL U34847 ( .A(n51365), .B(n42698), .Y(n28244) );
  XNOR2XL U34848 ( .A(n51368), .B(n42698), .Y(n28124) );
  XNOR2XL U34849 ( .A(n51407), .B(n42697), .Y(n29476) );
  XNOR2XL U34850 ( .A(n51359), .B(n42698), .Y(n28334) );
  XNOR2XL U34851 ( .A(n51371), .B(n42695), .Y(n24846) );
  XNOR2XL U34852 ( .A(n51354), .B(n42698), .Y(n28394) );
  XNOR2XL U34853 ( .A(n51361), .B(n42698), .Y(n28274) );
  XNOR2XL U34854 ( .A(n51360), .B(n42698), .Y(n28364) );
  XNOR2XL U34855 ( .A(n51351), .B(n42701), .Y(n31643) );
  XNOR2XL U34856 ( .A(n50715), .B(n36854), .Y(n23145) );
  XNOR2XL U34857 ( .A(n51404), .B(n42693), .Y(n29115) );
  XNOR2XL U34858 ( .A(n51411), .B(n42693), .Y(n29266) );
  XNOR2XL U34859 ( .A(n51408), .B(n42693), .Y(n29386) );
  XOR2XL U34860 ( .A(n41913), .B(n41313), .Y(n23226) );
  XOR2XL U34861 ( .A(n41917), .B(n41314), .Y(n23277) );
  XOR2XL U34862 ( .A(n41916), .B(n41317), .Y(n23236) );
  XNOR2XL U34863 ( .A(n49514), .B(n36793), .Y(n20408) );
  XNOR2XL U34864 ( .A(n50928), .B(n41295), .Y(n23183) );
  XNOR2XL U34865 ( .A(n50929), .B(n41293), .Y(n23143) );
  XNOR2XL U34866 ( .A(n50932), .B(n41296), .Y(n23123) );
  XOR2XL U34867 ( .A(n42061), .B(n42684), .Y(n43893) );
  XOR2XL U34868 ( .A(n42164), .B(n36882), .Y(n24937) );
  XOR2XL U34869 ( .A(n41905), .B(n36901), .Y(n24933) );
  XOR2XL U34870 ( .A(n42135), .B(n36880), .Y(n29116) );
  XOR2XL U34871 ( .A(n42136), .B(n42652), .Y(n29108) );
  XOR2XL U34872 ( .A(n42138), .B(n42652), .Y(n29018) );
  XOR2XL U34873 ( .A(n42165), .B(n42667), .Y(n24929) );
  XOR2XL U34874 ( .A(n41879), .B(n42601), .Y(n29014) );
  XOR2XL U34875 ( .A(n41877), .B(n42601), .Y(n29104) );
  XOR2XL U34876 ( .A(n41906), .B(n42605), .Y(n24925) );
  XOR2XL U34877 ( .A(n42153), .B(n36887), .Y(n27071) );
  XOR2XL U34878 ( .A(n41869), .B(n36901), .Y(n29263) );
  XOR2XL U34879 ( .A(n41878), .B(n36898), .Y(n29022) );
  XOR2XL U34880 ( .A(n42167), .B(n36882), .Y(n24757) );
  XOR2XL U34881 ( .A(n42144), .B(n36880), .Y(n26830) );
  XOR2XL U34882 ( .A(n41908), .B(n36897), .Y(n24753) );
  XOR2XL U34883 ( .A(n42137), .B(n36887), .Y(n29026) );
  XOR2XL U34884 ( .A(n42128), .B(n36887), .Y(n29267) );
  XOR2XL U34885 ( .A(n41870), .B(n42602), .Y(n29255) );
  XOR2XL U34886 ( .A(n41894), .B(n36892), .Y(n27067) );
  XOR2XL U34887 ( .A(n42166), .B(n36885), .Y(n24787) );
  XOR2XL U34888 ( .A(n41872), .B(n36895), .Y(n29383) );
  XOR2XL U34889 ( .A(n42132), .B(n42653), .Y(n29379) );
  XOR2XL U34890 ( .A(n41873), .B(n42602), .Y(n29375) );
  XOR2XL U34891 ( .A(n42168), .B(n42667), .Y(n24749) );
  XOR2XL U34892 ( .A(n41909), .B(n42608), .Y(n24745) );
  XOR2XL U34893 ( .A(n41885), .B(n36891), .Y(n26826) );
  XOR2XL U34894 ( .A(n42131), .B(n36886), .Y(n29387) );
  XOR2XL U34895 ( .A(n41895), .B(n42608), .Y(n27059) );
  XOR2XL U34896 ( .A(n42154), .B(n42662), .Y(n27063) );
  XOR2XL U34897 ( .A(n42169), .B(n36881), .Y(n24817) );
  XOR2XL U34898 ( .A(n41895), .B(n36895), .Y(n25083) );
  XOR2XL U34899 ( .A(n42154), .B(n36883), .Y(n25087) );
  XOR2XL U34900 ( .A(n41871), .B(n36898), .Y(n29413) );
  XOR2XL U34901 ( .A(n42155), .B(n36882), .Y(n25057) );
  XOR2XL U34902 ( .A(n41910), .B(n36893), .Y(n24813) );
  XOR2XL U34903 ( .A(n42130), .B(n36879), .Y(n29417) );
  XOR2XL U34904 ( .A(n42145), .B(n42661), .Y(n26822) );
  XOR2XL U34905 ( .A(n42131), .B(n42653), .Y(n29409) );
  XOR2XL U34906 ( .A(n41896), .B(n36891), .Y(n25053) );
  XOR2XL U34907 ( .A(n41886), .B(n42607), .Y(n26818) );
  XOR2XL U34908 ( .A(n41873), .B(n36892), .Y(n29473) );
  XOR2XL U34909 ( .A(n41872), .B(n42602), .Y(n29405) );
  XOR2XL U34910 ( .A(n41896), .B(n42607), .Y(n25075) );
  XOR2XL U34911 ( .A(n42155), .B(n42655), .Y(n25079) );
  XOR2XL U34912 ( .A(n42132), .B(n36881), .Y(n29477) );
  XOR2XL U34913 ( .A(n42133), .B(n42653), .Y(n29469) );
  XOR2XL U34914 ( .A(n41874), .B(n42602), .Y(n29465) );
  XOR2XL U34915 ( .A(n42170), .B(n42647), .Y(n24809) );
  XOR2XL U34916 ( .A(n42156), .B(n42667), .Y(n25049) );
  XOR2XL U34917 ( .A(n41911), .B(n36819), .Y(n24805) );
  XOR2XL U34918 ( .A(n41925), .B(n36901), .Y(n28421) );
  XOR2XL U34919 ( .A(n41897), .B(n42605), .Y(n25045) );
  XOR2XL U34920 ( .A(n42168), .B(n36880), .Y(n24847) );
  XOR2XL U34921 ( .A(n41925), .B(n42601), .Y(n28443) );
  XOR2XL U34922 ( .A(n42184), .B(n42652), .Y(n28447) );
  XOR2XL U34923 ( .A(n41924), .B(n36899), .Y(n28451) );
  XOR2XL U34924 ( .A(n42184), .B(n36883), .Y(n28425) );
  XOR2XL U34925 ( .A(n41909), .B(n36901), .Y(n24843) );
  XOR2XL U34926 ( .A(n41917), .B(n36891), .Y(n28571) );
  XOR2XL U34927 ( .A(n41926), .B(n36901), .Y(n28391) );
  XOR2XL U34928 ( .A(n42169), .B(n42663), .Y(n24839) );
  XOR2XL U34929 ( .A(n41918), .B(n42601), .Y(n28563) );
  XOR2XL U34930 ( .A(n42177), .B(n42652), .Y(n28567) );
  XOR2XL U34931 ( .A(n41910), .B(n36819), .Y(n24835) );
  XOR2XL U34932 ( .A(n42183), .B(n36882), .Y(n28455) );
  XOR2XL U34933 ( .A(n42176), .B(n36889), .Y(n28575) );
  XOR2XL U34934 ( .A(n42185), .B(n36887), .Y(n28395) );
  XOR2XL U34935 ( .A(n42150), .B(n36889), .Y(n27101) );
  XOR2XL U34936 ( .A(n41875), .B(n36901), .Y(n29082) );
  XOR2XL U34937 ( .A(n41876), .B(n42601), .Y(n29074) );
  XOR2XL U34938 ( .A(n42135), .B(n42652), .Y(n29078) );
  XOR2XL U34939 ( .A(n41916), .B(n36894), .Y(n28511) );
  XOR2XL U34940 ( .A(n42121), .B(n42662), .Y(n27364) );
  XOR2XL U34941 ( .A(n42134), .B(n36881), .Y(n29086) );
  XOR2XL U34942 ( .A(n42175), .B(n36879), .Y(n28515) );
  XOR2XL U34943 ( .A(n42176), .B(n42652), .Y(n28507) );
  XOR2XL U34944 ( .A(n41862), .B(n42608), .Y(n27360) );
  XOR2XL U34945 ( .A(n41917), .B(n42601), .Y(n28503) );
  XOR2XL U34946 ( .A(n41918), .B(n36897), .Y(n28541) );
  XOR2XL U34947 ( .A(n41891), .B(n36897), .Y(n27097) );
  XOR2XL U34948 ( .A(n42177), .B(n36885), .Y(n28545) );
  XOR2XL U34949 ( .A(n42178), .B(n42652), .Y(n28537) );
  XOR2XL U34950 ( .A(n41919), .B(n42601), .Y(n28533) );
  XOR2XL U34951 ( .A(n42151), .B(n42662), .Y(n27093) );
  XOR2XL U34952 ( .A(n41892), .B(n42608), .Y(n27089) );
  XOR2XL U34953 ( .A(n41923), .B(n36895), .Y(n28481) );
  XOR2XL U34954 ( .A(n42182), .B(n36882), .Y(n28485) );
  XOR2XL U34955 ( .A(n42183), .B(n42652), .Y(n28477) );
  XOR2XL U34956 ( .A(n42180), .B(n42652), .Y(n28357) );
  XOR2XL U34957 ( .A(n41921), .B(n42601), .Y(n28353) );
  XOR2XL U34958 ( .A(n41924), .B(n42601), .Y(n28473) );
  XOR2XL U34959 ( .A(n41929), .B(n36894), .Y(n31640) );
  XOR2XL U34960 ( .A(n42188), .B(n36882), .Y(n31644) );
  XOR2XL U34961 ( .A(n42189), .B(n42665), .Y(n31636) );
  XOR2XL U34962 ( .A(n41930), .B(n42608), .Y(n31632) );
  XOR2XL U34963 ( .A(n41927), .B(n36893), .Y(n31580) );
  XOR2XL U34964 ( .A(n42186), .B(n36880), .Y(n31584) );
  XOR2XL U34965 ( .A(n41934), .B(n36900), .Y(n31310) );
  XOR2XL U34966 ( .A(n42193), .B(n36888), .Y(n31314) );
  XOR2XL U34967 ( .A(n41935), .B(n36819), .Y(n31302) );
  XOR2XL U34968 ( .A(n42194), .B(n42656), .Y(n31306) );
  XOR2XL U34969 ( .A(n42187), .B(n42665), .Y(n31576) );
  XOR2XL U34970 ( .A(n41928), .B(n42608), .Y(n31572) );
  XOR2XL U34971 ( .A(n42104), .B(n36889), .Y(n28094) );
  XOR2XL U34972 ( .A(n41914), .B(n36900), .Y(n28211) );
  XOR2XL U34973 ( .A(n42173), .B(n36883), .Y(n28215) );
  XOR2XL U34974 ( .A(n41915), .B(n36900), .Y(n28241) );
  XOR2XL U34975 ( .A(n42174), .B(n36886), .Y(n28245) );
  XOR2XL U34976 ( .A(n41912), .B(n36893), .Y(n28121) );
  XOR2XL U34977 ( .A(n41921), .B(n36892), .Y(n28331) );
  XOR2XL U34978 ( .A(n42171), .B(n36886), .Y(n28125) );
  XOR2XL U34979 ( .A(n42180), .B(n36879), .Y(n28335) );
  XOR2XL U34980 ( .A(n41919), .B(n36895), .Y(n28271) );
  XOR2XL U34981 ( .A(n42178), .B(n36879), .Y(n28275) );
  XOR2XL U34982 ( .A(n41920), .B(n36892), .Y(n28361) );
  XOR2XL U34983 ( .A(n42179), .B(n36880), .Y(n28365) );
  XOR2XL U34984 ( .A(n42174), .B(n41286), .Y(n28207) );
  XOR2XL U34985 ( .A(n41915), .B(n42600), .Y(n28203) );
  XOR2XL U34986 ( .A(n41916), .B(n42600), .Y(n28233) );
  XOR2XL U34987 ( .A(n42175), .B(n41286), .Y(n28237) );
  XOR2XL U34988 ( .A(n42172), .B(n41286), .Y(n28117) );
  XOR2XL U34989 ( .A(n42181), .B(n41286), .Y(n28327) );
  XOR2XL U34990 ( .A(n41922), .B(n42600), .Y(n28323) );
  XOR2XL U34991 ( .A(n42185), .B(n41286), .Y(n28417) );
  XOR2XL U34992 ( .A(n41926), .B(n42600), .Y(n28413) );
  XOR2XL U34993 ( .A(n41927), .B(n42600), .Y(n28383) );
  XOR2XL U34994 ( .A(n42186), .B(n41286), .Y(n28387) );
  XOR2XL U34995 ( .A(n42179), .B(n41286), .Y(n28267) );
  XOR2XL U34996 ( .A(n41920), .B(n42600), .Y(n28263) );
  XNOR2XL U34997 ( .A(n51140), .B(n42554), .Y(n28401) );
  XNOR2XL U34998 ( .A(n51149), .B(n42554), .Y(n28491) );
  XNOR2XL U34999 ( .A(n51147), .B(n42554), .Y(n28521) );
  XNOR2XL U35000 ( .A(n51141), .B(n42554), .Y(n28431) );
  XNOR2XL U35001 ( .A(n50560), .B(n36780), .Y(n22471) );
  XNOR2XL U35002 ( .A(n51407), .B(n41300), .Y(n22361) );
  XNOR2XL U35003 ( .A(n50545), .B(n36783), .Y(n22321) );
  XNOR2XL U35004 ( .A(n51406), .B(n41302), .Y(n22371) );
  XNOR2XL U35005 ( .A(n51410), .B(n36741), .Y(n19538) );
  XNOR2XL U35006 ( .A(n51403), .B(n41304), .Y(n22341) );
  XNOR2XL U35007 ( .A(n51405), .B(n41299), .Y(n22381) );
  XNOR2XL U35008 ( .A(n51404), .B(n41302), .Y(n22391) );
  XOR2XL U35009 ( .A(n41902), .B(n42512), .Y(n25005) );
  XOR2XL U35010 ( .A(n41904), .B(n42525), .Y(n25155) );
  XOR2XL U35011 ( .A(n41860), .B(n42525), .Y(n27170) );
  XOR2XL U35012 ( .A(n41903), .B(n42525), .Y(n25185) );
  XOR2XL U35013 ( .A(n41905), .B(n42522), .Y(n24855) );
  XOR2XL U35014 ( .A(n41858), .B(n42525), .Y(n27230) );
  XOR2XL U35015 ( .A(n41859), .B(n42525), .Y(n27140) );
  XOR2XL U35016 ( .A(n41906), .B(n42522), .Y(n24885) );
  XOR2XL U35017 ( .A(n41862), .B(n42525), .Y(n27290) );
  XOR2XL U35018 ( .A(n41861), .B(n42525), .Y(n27200) );
  XOR2XL U35019 ( .A(n41857), .B(n42525), .Y(n27260) );
  XOR2XL U35020 ( .A(n41908), .B(n42512), .Y(n24945) );
  XOR2XL U35021 ( .A(n41894), .B(n42525), .Y(n27109) );
  XOR2XL U35022 ( .A(n41907), .B(n42528), .Y(n24915) );
  XOR2XL U35023 ( .A(n41897), .B(n42516), .Y(n25065) );
  XOR2XL U35024 ( .A(n41898), .B(n42525), .Y(n25035) );
  XOR2XL U35025 ( .A(n41896), .B(n42525), .Y(n27049) );
  XOR2XL U35026 ( .A(n41885), .B(n42522), .Y(n26838) );
  XOR2XL U35027 ( .A(n41869), .B(n42529), .Y(n29305) );
  XOR2XL U35028 ( .A(n41881), .B(n42522), .Y(n26778) );
  XOR2XL U35029 ( .A(n41883), .B(n42522), .Y(n26718) );
  XOR2XL U35030 ( .A(n41870), .B(n42529), .Y(n29335) );
  XOR2XL U35031 ( .A(n41879), .B(n42515), .Y(n29034) );
  XOR2XL U35032 ( .A(n41890), .B(n42522), .Y(n26929) );
  XOR2XL U35033 ( .A(n41891), .B(n42522), .Y(n26959) );
  XOR2XL U35034 ( .A(n41878), .B(n42515), .Y(n29094) );
  XOR2XL U35035 ( .A(n41872), .B(n42522), .Y(n29275) );
  XOR2XL U35036 ( .A(n41847), .B(n42522), .Y(n28072) );
  XOR2XL U35037 ( .A(n41886), .B(n42522), .Y(n26868) );
  XOR2XL U35038 ( .A(n41916), .B(n42522), .Y(n28193) );
  XOR2XL U35039 ( .A(n41892), .B(n42522), .Y(n26989) );
  XOR2XL U35040 ( .A(n41876), .B(n42516), .Y(n29425) );
  XOR2XL U35041 ( .A(n41895), .B(n42522), .Y(n27019) );
  XOR2XL U35042 ( .A(n41924), .B(n42518), .Y(n28283) );
  XOR2XL U35043 ( .A(n41912), .B(n42523), .Y(n24795) );
  XOR2XL U35044 ( .A(n41871), .B(n42516), .Y(n29245) );
  XOR2XL U35045 ( .A(n41914), .B(n42520), .Y(n28103) );
  XOR2XL U35046 ( .A(n41873), .B(n42516), .Y(n29395) );
  XOR2XL U35047 ( .A(n41880), .B(n42515), .Y(n29004) );
  XOR2XL U35048 ( .A(n41915), .B(n42522), .Y(n28163) );
  XOR2XL U35049 ( .A(n41887), .B(n42522), .Y(n26808) );
  XOR2XL U35050 ( .A(n41909), .B(n42523), .Y(n24765) );
  XOR2XL U35051 ( .A(n41910), .B(n42523), .Y(n24735) );
  XOR2XL U35052 ( .A(n41889), .B(n42522), .Y(n26899) );
  XOR2XL U35053 ( .A(n41874), .B(n42516), .Y(n29365) );
  XOR2XL U35054 ( .A(n41923), .B(n42518), .Y(n28313) );
  XOR2XL U35055 ( .A(n41875), .B(n42516), .Y(n29455) );
  XOR2XL U35056 ( .A(n41911), .B(n42523), .Y(n24825) );
  XOR2XL U35057 ( .A(n41863), .B(n42522), .Y(n27350) );
  XOR2XL U35058 ( .A(n41927), .B(n42515), .Y(n28403) );
  XOR2XL U35059 ( .A(n41918), .B(n42515), .Y(n28493) );
  XOR2XL U35060 ( .A(n41917), .B(n42522), .Y(n28223) );
  XOR2XL U35061 ( .A(n41921), .B(n42520), .Y(n28253) );
  XOR2XL U35062 ( .A(n41920), .B(n42515), .Y(n28523) );
  XOR2XL U35063 ( .A(n41928), .B(n42518), .Y(n28373) );
  XOR2XL U35064 ( .A(n41893), .B(n42522), .Y(n27079) );
  XOR2XL U35065 ( .A(n41877), .B(n42515), .Y(n29064) );
  XOR2XL U35066 ( .A(n41926), .B(n42515), .Y(n28433) );
  XOR2XL U35067 ( .A(n41919), .B(n42515), .Y(n28553) );
  XOR2XL U35068 ( .A(n41925), .B(n42515), .Y(n28463) );
  XOR2XL U35069 ( .A(n41922), .B(n42522), .Y(n28343) );
  XNOR2XL U35070 ( .A(n50935), .B(n42544), .Y(n28490) );
  XNOR2XL U35071 ( .A(n50925), .B(n42544), .Y(n28370) );
  XNOR2XL U35072 ( .A(n50933), .B(n42544), .Y(n28520) );
  XNOR2XL U35073 ( .A(n50927), .B(n42544), .Y(n28430) );
  XNOR2XL U35074 ( .A(n51206), .B(n41330), .Y(n23714) );
  XNOR2XL U35075 ( .A(n51207), .B(n41332), .Y(n23704) );
  XNOR2XL U35076 ( .A(n51220), .B(n41329), .Y(n23845) );
  XNOR2XL U35077 ( .A(n51162), .B(n36913), .Y(n23591) );
  XNOR2XL U35078 ( .A(n49516), .B(n41332), .Y(n23785) );
  XNOR2XL U35079 ( .A(n51208), .B(n41328), .Y(n23734) );
  XNOR2XL U35080 ( .A(n51221), .B(n41330), .Y(n23855) );
  XNOR2XL U35081 ( .A(n51214), .B(n41332), .Y(n23935) );
  XNOR2XL U35082 ( .A(n51205), .B(n41332), .Y(n23764) );
  XNOR2XL U35083 ( .A(n51209), .B(n41332), .Y(n23744) );
  XNOR2XL U35084 ( .A(n51218), .B(n41327), .Y(n23975) );
  XNOR2XL U35085 ( .A(n51216), .B(n41330), .Y(n23955) );
  XNOR2XL U35086 ( .A(n51201), .B(n41330), .Y(n22457) );
  XNOR2XL U35087 ( .A(n51219), .B(n41327), .Y(n23835) );
  XNOR2XL U35088 ( .A(n51204), .B(n36913), .Y(n23694) );
  XNOR2XL U35089 ( .A(n51211), .B(n41331), .Y(n23985) );
  XNOR2XL U35090 ( .A(n51196), .B(n41330), .Y(n22427) );
  XNOR2XL U35091 ( .A(n51200), .B(n36913), .Y(n22447) );
  XNOR2XL U35092 ( .A(n51174), .B(n36913), .Y(n24148) );
  XNOR2XL U35093 ( .A(n51176), .B(n41328), .Y(n24107) );
  XNOR2XL U35094 ( .A(n51195), .B(n41333), .Y(n22417) );
  XNOR2XL U35095 ( .A(n51224), .B(n41330), .Y(n23775) );
  XNOR2XL U35096 ( .A(n51202), .B(n41327), .Y(n22467) );
  XNOR2XL U35097 ( .A(n51187), .B(n41333), .Y(n22317) );
  XNOR2XL U35098 ( .A(n51179), .B(n36913), .Y(n24016) );
  XNOR2XL U35099 ( .A(n51171), .B(n41332), .Y(n24158) );
  XNOR2XL U35100 ( .A(n51197), .B(n41333), .Y(n22407) );
  XNOR2XL U35101 ( .A(n51194), .B(n41333), .Y(n22357) );
  XNOR2XL U35102 ( .A(n51172), .B(n41331), .Y(n24137) );
  XNOR2XL U35103 ( .A(n51177), .B(n41330), .Y(n24117) );
  XNOR2XL U35104 ( .A(n51184), .B(n41330), .Y(n24036) );
  XNOR2XL U35105 ( .A(n51183), .B(n41331), .Y(n24026) );
  XNOR2XL U35106 ( .A(n51160), .B(n41330), .Y(n23569) );
  XNOR2XL U35107 ( .A(n51215), .B(n41328), .Y(n23945) );
  XNOR2XL U35108 ( .A(n51193), .B(n41333), .Y(n22367) );
  XNOR2XL U35109 ( .A(n51185), .B(n41332), .Y(n24046) );
  XNOR2XL U35110 ( .A(n51203), .B(n41332), .Y(n23724) );
  XNOR2XL U35111 ( .A(n51197), .B(n36715), .Y(n19534) );
  XNOR2XL U35112 ( .A(n51186), .B(n41332), .Y(n24056) );
  XNOR2XL U35113 ( .A(n51217), .B(n36913), .Y(n23965) );
  XNOR2XL U35114 ( .A(n51182), .B(n41329), .Y(n24076) );
  XNOR2XL U35115 ( .A(n51190), .B(n41329), .Y(n22337) );
  XNOR2XL U35116 ( .A(n51161), .B(n41327), .Y(n23580) );
  XNOR2XL U35117 ( .A(n51168), .B(n41333), .Y(n23529) );
  XNOR2XL U35118 ( .A(n51163), .B(n41333), .Y(n23489) );
  XNOR2XL U35119 ( .A(n51170), .B(n41330), .Y(n23549) );
  XNOR2XL U35120 ( .A(n51192), .B(n41328), .Y(n22377) );
  XNOR2XL U35121 ( .A(n51169), .B(n41333), .Y(n23539) );
  XNOR2XL U35122 ( .A(n51156), .B(n41327), .Y(n23449) );
  XNOR2XL U35123 ( .A(n51173), .B(n41333), .Y(n24168) );
  XNOR2XL U35124 ( .A(n51191), .B(n41330), .Y(n22387) );
  XNOR2XL U35125 ( .A(n51167), .B(n41332), .Y(n235590) );
  XNOR2XL U35126 ( .A(n51181), .B(n41333), .Y(n24086) );
  XNOR2XL U35127 ( .A(n51205), .B(n36720), .Y(n20123) );
  XNOR2XL U35128 ( .A(n50778), .B(n36859), .Y(n23715) );
  XNOR2XL U35129 ( .A(n50779), .B(n36852), .Y(n23705) );
  XNOR2XL U35130 ( .A(n50792), .B(n36857), .Y(n23846) );
  XNOR2XL U35131 ( .A(n50734), .B(n36856), .Y(n23592) );
  XNOR2XL U35132 ( .A(n49513), .B(n36852), .Y(n23786) );
  XNOR2XL U35133 ( .A(n50793), .B(n36858), .Y(n23856) );
  XNOR2XL U35134 ( .A(n50780), .B(n36853), .Y(n23735) );
  XNOR2XL U35135 ( .A(n50786), .B(n36860), .Y(n23936) );
  XNOR2XL U35136 ( .A(n50777), .B(n36852), .Y(n23765) );
  XNOR2XL U35137 ( .A(n50781), .B(n36858), .Y(n23745) );
  XNOR2XL U35138 ( .A(n50790), .B(n36851), .Y(n23976) );
  XNOR2XL U35139 ( .A(n50791), .B(n36852), .Y(n23836) );
  XNOR2XL U35140 ( .A(n50788), .B(n36850), .Y(n23956) );
  XNOR2XL U35141 ( .A(n50773), .B(n36857), .Y(n22458) );
  XNOR2XL U35142 ( .A(n50783), .B(n36860), .Y(n23986) );
  XNOR2XL U35143 ( .A(n50776), .B(n36854), .Y(n23695) );
  XNOR2XL U35144 ( .A(n50768), .B(n36854), .Y(n22428) );
  XNOR2XL U35145 ( .A(n50772), .B(n36852), .Y(n22448) );
  XNOR2XL U35146 ( .A(n50767), .B(n36860), .Y(n22418) );
  XNOR2XL U35147 ( .A(n50746), .B(n36859), .Y(n24149) );
  XNOR2XL U35148 ( .A(n50748), .B(n36852), .Y(n24108) );
  XNOR2XL U35149 ( .A(n50796), .B(n36853), .Y(n23776) );
  XNOR2XL U35150 ( .A(n50774), .B(n36859), .Y(n22468) );
  XNOR2XL U35151 ( .A(n50759), .B(n36857), .Y(n22318) );
  XNOR2XL U35152 ( .A(n50751), .B(n36851), .Y(n24017) );
  XNOR2XL U35153 ( .A(n50769), .B(n36850), .Y(n22408) );
  XNOR2XL U35154 ( .A(n50743), .B(n36859), .Y(n24159) );
  XNOR2XL U35155 ( .A(n50749), .B(n36857), .Y(n24118) );
  XNOR2XL U35156 ( .A(n50766), .B(n36856), .Y(n22358) );
  XNOR2XL U35157 ( .A(n50744), .B(n36859), .Y(n24138) );
  XNOR2XL U35158 ( .A(n50756), .B(n36851), .Y(n24037) );
  XNOR2XL U35159 ( .A(n50755), .B(n36854), .Y(n24027) );
  XNOR2XL U35160 ( .A(n50787), .B(n36860), .Y(n23946) );
  XNOR2XL U35161 ( .A(n50732), .B(n36853), .Y(n23570) );
  XNOR2XL U35162 ( .A(n50765), .B(n36859), .Y(n22368) );
  XNOR2XL U35163 ( .A(n50757), .B(n36859), .Y(n24047) );
  XNOR2XL U35164 ( .A(n50775), .B(n36859), .Y(n23725) );
  XNOR2XL U35165 ( .A(n50758), .B(n36854), .Y(n24057) );
  XNOR2XL U35166 ( .A(n50769), .B(n42465), .Y(n19535) );
  XNOR2XL U35167 ( .A(n50789), .B(n36854), .Y(n23966) );
  XNOR2XL U35168 ( .A(n50754), .B(n36852), .Y(n24077) );
  XNOR2XL U35169 ( .A(n50733), .B(n36858), .Y(n23581) );
  XNOR2XL U35170 ( .A(n50740), .B(n36852), .Y(n23530) );
  XNOR2XL U35171 ( .A(n50735), .B(n36853), .Y(n23490) );
  XNOR2XL U35172 ( .A(n50742), .B(n36853), .Y(n23550) );
  XNOR2XL U35173 ( .A(n50762), .B(n36851), .Y(n22338) );
  XNOR2XL U35174 ( .A(n50764), .B(n36851), .Y(n22378) );
  XNOR2XL U35175 ( .A(n50741), .B(n36860), .Y(n23540) );
  XNOR2XL U35176 ( .A(n50745), .B(n36850), .Y(n24169) );
  XNOR2XL U35177 ( .A(n50728), .B(n36858), .Y(n23450) );
  XNOR2XL U35178 ( .A(n50763), .B(n36858), .Y(n22388) );
  XNOR2XL U35179 ( .A(n50753), .B(n36856), .Y(n24087) );
  XNOR2XL U35180 ( .A(n50358), .B(n42705), .Y(n29234) );
  XNOR2XL U35181 ( .A(n50351), .B(n42705), .Y(n29294) );
  XNOR2XL U35182 ( .A(n50345), .B(n42704), .Y(n29113) );
  XNOR2XL U35183 ( .A(n50352), .B(n42707), .Y(n29264) );
  XNOR2XL U35184 ( .A(n50349), .B(n41642), .Y(n29384) );
  XNOR2XL U35185 ( .A(n50350), .B(n42707), .Y(n29414) );
  XNOR2XL U35186 ( .A(n51009), .B(n42618), .Y(n27989) );
  XNOR2XL U35187 ( .A(n51002), .B(n36870), .Y(n27576) );
  XNOR2XL U35188 ( .A(n50369), .B(n42675), .Y(n27572) );
  XNOR2XL U35189 ( .A(n50963), .B(n42615), .Y(n26966) );
  XNOR2XL U35190 ( .A(n50959), .B(n42615), .Y(n27026) );
  XNOR2XL U35191 ( .A(n50319), .B(n36907), .Y(n25196) );
  XNOR2XL U35192 ( .A(n50999), .B(n42618), .Y(n27508) );
  XNOR2XL U35193 ( .A(n50332), .B(n42674), .Y(n26940) );
  XNOR2XL U35194 ( .A(n50965), .B(net219330), .Y(n26944) );
  XNOR2XL U35195 ( .A(n50316), .B(n42675), .Y(n24896) );
  XNOR2XL U35196 ( .A(n50997), .B(n42615), .Y(n27267) );
  XNOR2XL U35197 ( .A(n50930), .B(n42619), .Y(n28290) );
  XNOR2XL U35198 ( .A(n50962), .B(n42615), .Y(n26996) );
  XNOR2XL U35199 ( .A(n50949), .B(n40039), .Y(n24900) );
  XNOR2XL U35200 ( .A(n50993), .B(n42615), .Y(n27207) );
  XNOR2XL U35201 ( .A(n51010), .B(net219308), .Y(n27997) );
  XNOR2XL U35202 ( .A(n50965), .B(n36868), .Y(n26906) );
  XNOR2XL U35203 ( .A(n50377), .B(n42675), .Y(n27993) );
  XNOR2XL U35204 ( .A(n50328), .B(n42674), .Y(n27120) );
  XNOR2XL U35205 ( .A(n50961), .B(net219324), .Y(n27124) );
  XNOR2XL U35206 ( .A(n50939), .B(n42619), .Y(n28170) );
  XNOR2XL U35207 ( .A(n50990), .B(n42618), .Y(n27327) );
  XNOR2XL U35208 ( .A(n50331), .B(n42674), .Y(n26970) );
  XNOR2XL U35209 ( .A(n51007), .B(n42619), .Y(n28079) );
  XNOR2XL U35210 ( .A(n51000), .B(net219330), .Y(n27516) );
  XNOR2XL U35211 ( .A(n50367), .B(n42675), .Y(n27512) );
  XNOR2XL U35212 ( .A(n50327), .B(n42674), .Y(n27030) );
  XNOR2XL U35213 ( .A(n50960), .B(n40039), .Y(n27034) );
  XNOR2XL U35214 ( .A(n50964), .B(net219336), .Y(n26974) );
  XNOR2XL U35215 ( .A(n50998), .B(net219310), .Y(n27275) );
  XNOR2XL U35216 ( .A(n50365), .B(n42674), .Y(n27271) );
  XNOR2XL U35217 ( .A(n50966), .B(n36870), .Y(n26914) );
  XNOR2XL U35218 ( .A(n50298), .B(n42671), .Y(n28294) );
  XNOR2XL U35219 ( .A(n50330), .B(n42674), .Y(n27000) );
  XNOR2XL U35220 ( .A(n50963), .B(net219310), .Y(n27004) );
  XNOR2XL U35221 ( .A(n50299), .B(n42712), .Y(n28302) );
  XNOR2XL U35222 ( .A(n50969), .B(net219324), .Y(n26883) );
  XNOR2XL U35223 ( .A(n50333), .B(n42670), .Y(n26910) );
  XNOR2XL U35224 ( .A(n50361), .B(n42674), .Y(n27211) );
  XNOR2XL U35225 ( .A(n50994), .B(net219308), .Y(n27215) );
  XNOR2XL U35226 ( .A(n51005), .B(n42618), .Y(n27388) );
  XNOR2XL U35227 ( .A(n50307), .B(n42671), .Y(n28174) );
  XNOR2XL U35228 ( .A(n50358), .B(n42675), .Y(n27331) );
  XNOR2XL U35229 ( .A(n50991), .B(n36870), .Y(n27335) );
  XNOR2XL U35230 ( .A(n50938), .B(n42619), .Y(n28200) );
  XNOR2XL U35231 ( .A(n50308), .B(n42712), .Y(n28182) );
  XNOR2XL U35232 ( .A(n50375), .B(n42671), .Y(n28083) );
  XNOR2XL U35233 ( .A(n50947), .B(n40039), .Y(n24960) );
  XNOR2XL U35234 ( .A(n50376), .B(n42712), .Y(n28091) );
  XNOR2XL U35235 ( .A(n50958), .B(n42615), .Y(n27056) );
  XNOR2XL U35236 ( .A(n50948), .B(net219324), .Y(n24930) );
  XNOR2XL U35237 ( .A(n50937), .B(n42619), .Y(n28230) );
  XNOR2XL U35238 ( .A(n50967), .B(n36868), .Y(n26815) );
  XNOR2XL U35239 ( .A(n50940), .B(n42619), .Y(n28110) );
  XNOR2XL U35240 ( .A(n50931), .B(n42619), .Y(n28320) );
  XNOR2XL U35241 ( .A(n50307), .B(n42712), .Y(n28212) );
  XNOR2XL U35242 ( .A(n50957), .B(n42613), .Y(n25072) );
  XNOR2XL U35243 ( .A(n50373), .B(n42675), .Y(n27392) );
  XNOR2XL U35244 ( .A(n51006), .B(net219310), .Y(n27396) );
  XNOR2XL U35245 ( .A(n50306), .B(n42671), .Y(n28204) );
  XNOR2XL U35246 ( .A(n50956), .B(n42618), .Y(n25042) );
  XNOR2XL U35247 ( .A(n50945), .B(n42615), .Y(n24772) );
  XNOR2XL U35248 ( .A(n50326), .B(n42674), .Y(n27060) );
  XNOR2XL U35249 ( .A(n50959), .B(net219336), .Y(n27064) );
  XNOR2XL U35250 ( .A(n50968), .B(n40039), .Y(n26823) );
  XNOR2XL U35251 ( .A(n50927), .B(n42619), .Y(n28410) );
  XNOR2XL U35252 ( .A(n50305), .B(n36907), .Y(n28234) );
  XNOR2XL U35253 ( .A(n50300), .B(n42712), .Y(n28332) );
  XNOR2XL U35254 ( .A(n50306), .B(n42712), .Y(n28242) );
  XNOR2XL U35255 ( .A(n50308), .B(n42671), .Y(n28114) );
  XNOR2XL U35256 ( .A(n50299), .B(n42674), .Y(n28324) );
  XNOR2XL U35257 ( .A(n50942), .B(n42615), .Y(n24802) );
  XNOR2XL U35258 ( .A(n50979), .B(n42615), .Y(n29462) );
  XNOR2XL U35259 ( .A(n50957), .B(net219310), .Y(n25050) );
  XNOR2XL U35260 ( .A(n50325), .B(n42674), .Y(n25076) );
  XNOR2XL U35261 ( .A(n50958), .B(net219310), .Y(n25080) );
  XNOR2XL U35262 ( .A(n50324), .B(n42673), .Y(n25046) );
  XNOR2XL U35263 ( .A(n50991), .B(n42618), .Y(n27357) );
  XNOR2XL U35264 ( .A(n50946), .B(n40039), .Y(n24780) );
  XNOR2XL U35265 ( .A(n50943), .B(n42617), .Y(n24832) );
  XNOR2XL U35266 ( .A(n50933), .B(n42619), .Y(n28260) );
  XNOR2XL U35267 ( .A(n50295), .B(n42671), .Y(n28414) );
  XNOR2XL U35268 ( .A(n50348), .B(n42712), .Y(n29474) );
  XNOR2XL U35269 ( .A(n50961), .B(n42615), .Y(n27086) );
  XNOR2XL U35270 ( .A(n50347), .B(n42671), .Y(n29466) );
  XNOR2XL U35271 ( .A(n50295), .B(n42712), .Y(n28392) );
  XNOR2XL U35272 ( .A(n50992), .B(net219330), .Y(n27365) );
  XNOR2XL U35273 ( .A(n50302), .B(n42712), .Y(n28272) );
  XNOR2XL U35274 ( .A(n50359), .B(n42675), .Y(n27361) );
  XNOR2XL U35275 ( .A(n50301), .B(n42671), .Y(n28264) );
  XNOR2XL U35276 ( .A(n50312), .B(n42708), .Y(n24844) );
  XNOR2XL U35277 ( .A(n50944), .B(net219314), .Y(n24840) );
  XNOR2XL U35278 ( .A(n50962), .B(net258262), .Y(n27094) );
  XNOR2XL U35279 ( .A(n50932), .B(n42619), .Y(n28350) );
  XNOR2XL U35280 ( .A(n50329), .B(n42674), .Y(n27090) );
  XNOR2XL U35281 ( .A(n50300), .B(n42671), .Y(n28354) );
  XNOR2XL U35282 ( .A(n50301), .B(n42712), .Y(n28362) );
  XNOR2XL U35283 ( .A(n50923), .B(n42617), .Y(n31629) );
  XNOR2XL U35284 ( .A(n50920), .B(n42617), .Y(n31389) );
  XNOR2XL U35285 ( .A(n50291), .B(n42670), .Y(n31633) );
  XNOR2XL U35286 ( .A(n50989), .B(n41284), .Y(n29222) );
  XNOR2XL U35287 ( .A(n50356), .B(n42671), .Y(n29196) );
  XNOR2XL U35288 ( .A(n50985), .B(n41284), .Y(n29312) );
  XNOR2XL U35289 ( .A(n50352), .B(n42671), .Y(n29346) );
  XNOR2XL U35290 ( .A(n50357), .B(n42671), .Y(n29226) );
  XNOR2XL U35291 ( .A(n50982), .B(n41284), .Y(n29282) );
  XNOR2XL U35292 ( .A(n50353), .B(n42671), .Y(n29316) );
  XNOR2XL U35293 ( .A(n50350), .B(n42671), .Y(n29286) );
  XNOR2XL U35294 ( .A(n50976), .B(n41284), .Y(n29101) );
  XNOR2XL U35295 ( .A(n50983), .B(n41284), .Y(n29252) );
  XNOR2XL U35296 ( .A(n50980), .B(n41284), .Y(n29372) );
  XNOR2XL U35297 ( .A(n50344), .B(n36907), .Y(n29105) );
  XNOR2XL U35298 ( .A(n50981), .B(n41284), .Y(n29402) );
  XNOR2XL U35299 ( .A(n50351), .B(n42671), .Y(n29256) );
  XNOR2XL U35300 ( .A(n50348), .B(n42669), .Y(n29376) );
  XNOR2XL U35301 ( .A(n50349), .B(n42670), .Y(n29406) );
  XNOR2XL U35302 ( .A(n50992), .B(n41295), .Y(n23713) );
  XNOR2XL U35303 ( .A(n51006), .B(n41293), .Y(n23844) );
  XNOR2XL U35304 ( .A(n50993), .B(n41290), .Y(n23703) );
  XNOR2XL U35305 ( .A(n50948), .B(n41294), .Y(n23590) );
  XNOR2XL U35306 ( .A(n49514), .B(n41291), .Y(n23784) );
  XNOR2XL U35307 ( .A(n50994), .B(n41293), .Y(n23733) );
  XNOR2XL U35308 ( .A(n51007), .B(n41293), .Y(n23854) );
  XNOR2XL U35309 ( .A(n51000), .B(n41296), .Y(n23934) );
  XNOR2XL U35310 ( .A(n50991), .B(n41297), .Y(n23763) );
  XNOR2XL U35311 ( .A(n50995), .B(n41290), .Y(n23743) );
  XNOR2XL U35312 ( .A(n51004), .B(n41292), .Y(n23974) );
  XNOR2XL U35313 ( .A(n51002), .B(n41294), .Y(n23954) );
  XNOR2XL U35314 ( .A(n50987), .B(n41293), .Y(n22456) );
  XNOR2XL U35315 ( .A(n50990), .B(n41291), .Y(n23693) );
  XNOR2XL U35316 ( .A(n51005), .B(n41296), .Y(n23834) );
  XNOR2XL U35317 ( .A(n50982), .B(n41291), .Y(n22426) );
  XNOR2XL U35318 ( .A(n50997), .B(n41290), .Y(n23984) );
  XNOR2XL U35319 ( .A(n50986), .B(n41294), .Y(n22446) );
  XNOR2XL U35320 ( .A(n50960), .B(n41294), .Y(n24147) );
  XNOR2XL U35321 ( .A(n50962), .B(n41296), .Y(n24106) );
  XNOR2XL U35322 ( .A(n50981), .B(n41294), .Y(n22416) );
  XNOR2XL U35323 ( .A(n51010), .B(n36916), .Y(n23774) );
  XNOR2XL U35324 ( .A(n50988), .B(n41294), .Y(n22466) );
  XNOR2XL U35325 ( .A(n50973), .B(n41290), .Y(n22316) );
  XNOR2XL U35326 ( .A(n50965), .B(n41292), .Y(n24015) );
  XNOR2XL U35327 ( .A(n50957), .B(n41294), .Y(n24157) );
  XNOR2XL U35328 ( .A(n50983), .B(n41291), .Y(n22406) );
  XNOR2XL U35329 ( .A(n50980), .B(n41291), .Y(n22356) );
  XNOR2XL U35330 ( .A(n50958), .B(n41290), .Y(n24136) );
  XNOR2XL U35331 ( .A(n50963), .B(n41290), .Y(n24116) );
  XNOR2XL U35332 ( .A(n50970), .B(n41295), .Y(n24035) );
  XNOR2XL U35333 ( .A(n50946), .B(n41293), .Y(n23568) );
  XNOR2XL U35334 ( .A(n50969), .B(n41290), .Y(n24025) );
  XNOR2XL U35335 ( .A(n51001), .B(n41292), .Y(n23944) );
  XNOR2XL U35336 ( .A(n50971), .B(n41297), .Y(n24045) );
  XNOR2XL U35337 ( .A(n50979), .B(n41293), .Y(n22366) );
  XNOR2XL U35338 ( .A(n50983), .B(n36790), .Y(n19533) );
  XNOR2XL U35339 ( .A(n50989), .B(n41291), .Y(n23723) );
  XNOR2XL U35340 ( .A(n50972), .B(n41293), .Y(n24055) );
  XNOR2XL U35341 ( .A(n50968), .B(n41296), .Y(n24075) );
  XNOR2XL U35342 ( .A(n51003), .B(n41296), .Y(n23964) );
  XNOR2XL U35343 ( .A(n50976), .B(n41291), .Y(n22336) );
  XNOR2XL U35344 ( .A(n50954), .B(n41294), .Y(n23528) );
  XNOR2XL U35345 ( .A(n50947), .B(n41292), .Y(n23579) );
  XNOR2XL U35346 ( .A(n50949), .B(n41296), .Y(n23488) );
  XNOR2XL U35347 ( .A(n50956), .B(n41293), .Y(n23548) );
  XNOR2XL U35348 ( .A(n50978), .B(n41296), .Y(n22376) );
  XNOR2XL U35349 ( .A(n50955), .B(n41291), .Y(n23538) );
  XNOR2XL U35350 ( .A(n50942), .B(n41295), .Y(n23448) );
  XNOR2XL U35351 ( .A(n50959), .B(n41290), .Y(n24167) );
  XNOR2XL U35352 ( .A(n50953), .B(n41296), .Y(n235580) );
  XNOR2XL U35353 ( .A(n50977), .B(n41291), .Y(n22386) );
  XNOR2XL U35354 ( .A(n50991), .B(n36798), .Y(n20122) );
  XNOR2XL U35355 ( .A(n50967), .B(n41293), .Y(n24085) );
  XNOR2XL U35356 ( .A(n50554), .B(n42717), .Y(n29415) );
  XNOR2XL U35357 ( .A(n50975), .B(net258262), .Y(n29019) );
  XNOR2XL U35358 ( .A(n51189), .B(n41281), .Y(n29020) );
  XNOR2XL U35359 ( .A(n50761), .B(net219468), .Y(n29021) );
  XNOR2XL U35360 ( .A(n50750), .B(n36863), .Y(n26938) );
  XNOR2XL U35361 ( .A(n50740), .B(n36730), .Y(n25124) );
  XNOR2XL U35362 ( .A(n51422), .B(n42641), .Y(n27153) );
  XNOR2XL U35363 ( .A(n50738), .B(n36731), .Y(n24974) );
  XNOR2XL U35364 ( .A(n50734), .B(n36865), .Y(n24894) );
  XNOR2XL U35365 ( .A(n50737), .B(n36865), .Y(n25194) );
  XNOR2XL U35366 ( .A(n50755), .B(n36865), .Y(n26847) );
  XNOR2XL U35367 ( .A(n50777), .B(net219466), .Y(n27337) );
  XNOR2XL U35368 ( .A(n50746), .B(n36863), .Y(n27118) );
  XNOR2XL U35369 ( .A(n50734), .B(net258207), .Y(n24932) );
  XNOR2XL U35370 ( .A(n51428), .B(n42642), .Y(n27574) );
  XNOR2XL U35371 ( .A(n50795), .B(n42592), .Y(n27991) );
  XNOR2XL U35372 ( .A(n51391), .B(n42641), .Y(n26942) );
  XNOR2XL U35373 ( .A(n50745), .B(n36863), .Y(n27028) );
  XNOR2XL U35374 ( .A(n49511), .B(n36903), .Y(n27724) );
  XNOR2XL U35375 ( .A(n51378), .B(n36861), .Y(n25198) );
  XNOR2XL U35376 ( .A(n51396), .B(n36867), .Y(n26851) );
  XNOR2XL U35377 ( .A(n50749), .B(n36863), .Y(n26968) );
  XNOR2XL U35378 ( .A(n51375), .B(n36867), .Y(n24898) );
  XNOR2XL U35379 ( .A(n51213), .B(n42554), .Y(n27589) );
  XNOR2XL U35380 ( .A(n50785), .B(n42592), .Y(n27510) );
  XNOR2XL U35381 ( .A(n50716), .B(n42586), .Y(n28292) );
  XNOR2XL U35382 ( .A(n50748), .B(n36863), .Y(n26998) );
  XNOR2XL U35383 ( .A(n51387), .B(n42641), .Y(n27122) );
  XNOR2XL U35384 ( .A(n50754), .B(n36865), .Y(n26877) );
  XNOR2XL U35385 ( .A(n51165), .B(n42551), .Y(n25003) );
  XNOR2XL U35386 ( .A(n50779), .B(n36863), .Y(n27209) );
  XNOR2XL U35387 ( .A(n50745), .B(net219450), .Y(n27066) );
  XNOR2XL U35388 ( .A(n50783), .B(n36863), .Y(n27269) );
  XNOR2XL U35389 ( .A(n51163), .B(n42551), .Y(n25153) );
  XNOR2XL U35390 ( .A(n51436), .B(n42642), .Y(n27995) );
  XNOR2XL U35391 ( .A(n50754), .B(net219434), .Y(n26825) );
  XNOR2XL U35392 ( .A(n50725), .B(n42589), .Y(n28172) );
  XNOR2XL U35393 ( .A(n50776), .B(n42592), .Y(n27329) );
  XNOR2XL U35394 ( .A(n50751), .B(n36865), .Y(n26908) );
  XNOR2XL U35395 ( .A(n51386), .B(n42641), .Y(n27032) );
  XNOR2XL U35396 ( .A(n51390), .B(n42641), .Y(n26972) );
  XNOR2XL U35397 ( .A(n50793), .B(n42586), .Y(n28081) );
  XNOR2XL U35398 ( .A(n51221), .B(n42553), .Y(n28010) );
  XNOR2XL U35399 ( .A(n50744), .B(net258207), .Y(n25082) );
  XNOR2XL U35400 ( .A(n51426), .B(n42642), .Y(n27514) );
  XNOR2XL U35401 ( .A(n51179), .B(n42552), .Y(n26656) );
  XNOR2XL U35402 ( .A(n51182), .B(n42552), .Y(n26836) );
  XNOR2XL U35403 ( .A(n50743), .B(net258207), .Y(n25052) );
  XNOR2XL U35404 ( .A(n51357), .B(n42643), .Y(n28296) );
  XNOR2XL U35405 ( .A(n51389), .B(n42641), .Y(n27002) );
  XNOR2XL U35406 ( .A(n51214), .B(n42547), .Y(n27559) );
  XNOR2XL U35407 ( .A(n51420), .B(n42641), .Y(n27213) );
  XNOR2XL U35408 ( .A(n51424), .B(n42641), .Y(n27273) );
  XNOR2XL U35409 ( .A(n51392), .B(n36867), .Y(n26912) );
  XNOR2XL U35410 ( .A(n51417), .B(n42642), .Y(n27333) );
  XNOR2XL U35411 ( .A(n51366), .B(n42643), .Y(n28176) );
  XNOR2XL U35412 ( .A(n51434), .B(n42643), .Y(n28085) );
  XNOR2XL U35413 ( .A(n51186), .B(n42552), .Y(n26776) );
  XNOR2XL U35414 ( .A(n50730), .B(net219468), .Y(n24842) );
  XNOR2XL U35415 ( .A(n51208), .B(n42552), .Y(n27138) );
  XNOR2XL U35416 ( .A(n50724), .B(n36865), .Y(n28202) );
  XNOR2XL U35417 ( .A(n51212), .B(n42552), .Y(n27499) );
  XNOR2XL U35418 ( .A(n50744), .B(n36863), .Y(n27058) );
  XNOR2XL U35419 ( .A(n51164), .B(n42551), .Y(n25183) );
  XNOR2XL U35420 ( .A(n51374), .B(n42637), .Y(n24928) );
  XNOR2XL U35421 ( .A(n50723), .B(n36865), .Y(n28232) );
  XNOR2XL U35422 ( .A(n51162), .B(n42551), .Y(n24853) );
  XNOR2XL U35423 ( .A(n51184), .B(n42552), .Y(n26716) );
  XNOR2XL U35424 ( .A(n50778), .B(net219466), .Y(n27367) );
  XNOR2XL U35425 ( .A(n50753), .B(n36865), .Y(n26817) );
  XNOR2XL U35426 ( .A(n51222), .B(n42553), .Y(n27980) );
  XNOR2XL U35427 ( .A(n51183), .B(n42552), .Y(n26686) );
  XNOR2XL U35428 ( .A(n50743), .B(n42590), .Y(n25074) );
  XNOR2XL U35429 ( .A(n50726), .B(n34450), .Y(n28112) );
  XNOR2XL U35430 ( .A(n51177), .B(n42552), .Y(n26927) );
  XNOR2XL U35431 ( .A(n50717), .B(n42589), .Y(n28322) );
  XNOR2XL U35432 ( .A(n51365), .B(n42643), .Y(n28206) );
  XNOR2XL U35433 ( .A(n51205), .B(n42551), .Y(n27288) );
  XNOR2XL U35434 ( .A(n51406), .B(n42637), .Y(n29468) );
  XNOR2XL U35435 ( .A(n51385), .B(n42641), .Y(n27062) );
  XNOR2XL U35436 ( .A(n50748), .B(net219444), .Y(n27096) );
  XNOR2XL U35437 ( .A(n50742), .B(n36865), .Y(n25044) );
  XNOR2XL U35438 ( .A(n51176), .B(n42552), .Y(n26957) );
  XNOR2XL U35439 ( .A(n51364), .B(n42643), .Y(n28236) );
  XNOR2XL U35440 ( .A(n51161), .B(n42551), .Y(n24883) );
  XNOR2XL U35441 ( .A(n51197), .B(n42552), .Y(n29333) );
  XNOR2XL U35442 ( .A(n51394), .B(n36867), .Y(n26821) );
  XNOR2XL U35443 ( .A(n51206), .B(n36832), .Y(n27198) );
  XNOR2XL U35444 ( .A(n51210), .B(n36832), .Y(n27258) );
  XNOR2XL U35445 ( .A(n51175), .B(n42552), .Y(n26987) );
  XNOR2XL U35446 ( .A(n51173), .B(n42552), .Y(n27107) );
  XNOR2XL U35447 ( .A(n51384), .B(n36867), .Y(n25078) );
  XNOR2XL U35448 ( .A(n50713), .B(n42588), .Y(n28412) );
  XNOR2XL U35449 ( .A(n51181), .B(n42552), .Y(n26866) );
  XNOR2XL U35450 ( .A(n51358), .B(n42643), .Y(n28326) );
  XNOR2XL U35451 ( .A(n51220), .B(n42553), .Y(n28070) );
  XNOR2XL U35452 ( .A(n51203), .B(n36832), .Y(n27318) );
  XNOR2XL U35453 ( .A(n51383), .B(n36867), .Y(n25048) );
  XNOR2XL U35454 ( .A(n51188), .B(n42550), .Y(n29032) );
  XNOR2XL U35455 ( .A(n51172), .B(n42552), .Y(n27017) );
  XNOR2XL U35456 ( .A(n51151), .B(n42553), .Y(n28191) );
  XNOR2XL U35457 ( .A(n50765), .B(n42586), .Y(n29464) );
  XNOR2XL U35458 ( .A(n50777), .B(n42592), .Y(n27359) );
  XNOR2XL U35459 ( .A(n51143), .B(n42553), .Y(n28281) );
  XNOR2XL U35460 ( .A(n51159), .B(n42551), .Y(n24943) );
  XNOR2XL U35461 ( .A(n50729), .B(n36863), .Y(n24834) );
  XNOR2XL U35462 ( .A(n50719), .B(n36865), .Y(n28262) );
  XNOR2XL U35463 ( .A(n51354), .B(n42643), .Y(n28416) );
  XNOR2XL U35464 ( .A(n51195), .B(n42551), .Y(n29273) );
  XNOR2XL U35465 ( .A(n51189), .B(n42552), .Y(n29092) );
  XNOR2XL U35466 ( .A(n51160), .B(n42551), .Y(n24913) );
  XNOR2XL U35467 ( .A(n51153), .B(n42553), .Y(n28101) );
  XNOR2XL U35468 ( .A(n51152), .B(n42553), .Y(n28161) );
  XNOR2XL U35469 ( .A(n51191), .B(n36832), .Y(n29423) );
  XNOR2XL U35470 ( .A(n50747), .B(n36863), .Y(n27088) );
  XNOR2XL U35471 ( .A(n51180), .B(n42552), .Y(n26806) );
  XNOR2XL U35472 ( .A(n51218), .B(n36832), .Y(n27379) );
  XNOR2XL U35473 ( .A(n51418), .B(n42642), .Y(n27363) );
  XNOR2XL U35474 ( .A(n51360), .B(n42643), .Y(n28266) );
  XNOR2XL U35475 ( .A(n51178), .B(n42552), .Y(n26897) );
  XNOR2XL U35476 ( .A(n51170), .B(n42551), .Y(n25063) );
  XNOR2XL U35477 ( .A(n51171), .B(n42552), .Y(n27047) );
  XNOR2XL U35478 ( .A(n51169), .B(n42551), .Y(n25033) );
  XNOR2XL U35479 ( .A(n51196), .B(n42554), .Y(n29243) );
  XNOR2XL U35480 ( .A(n51194), .B(n42552), .Y(n29393) );
  XNOR2XL U35481 ( .A(n50718), .B(n42588), .Y(n28352) );
  XNOR2XL U35482 ( .A(n51155), .B(n42552), .Y(n24793) );
  XNOR2XL U35483 ( .A(n51388), .B(n42641), .Y(n27092) );
  XNOR2XL U35484 ( .A(n51144), .B(n42553), .Y(n28311) );
  XNOR2XL U35485 ( .A(n51204), .B(n42551), .Y(n27348) );
  XNOR2XL U35486 ( .A(n51157), .B(n42548), .Y(n24733) );
  XNOR2XL U35487 ( .A(n51193), .B(n42550), .Y(n29363) );
  XNOR2XL U35488 ( .A(n51150), .B(n42553), .Y(n28221) );
  XNOR2XL U35489 ( .A(n51158), .B(n42550), .Y(n24763) );
  XNOR2XL U35490 ( .A(n51359), .B(n42643), .Y(n28356) );
  XNOR2XL U35491 ( .A(n51139), .B(n42553), .Y(n28371) );
  XNOR2XL U35492 ( .A(n51146), .B(n42553), .Y(n28251) );
  XNOR2XL U35493 ( .A(n51174), .B(n42552), .Y(n27077) );
  XNOR2XL U35494 ( .A(n51156), .B(n42552), .Y(n24823) );
  XNOR2XL U35495 ( .A(n51350), .B(n36867), .Y(n31635) );
  XNOR2XL U35496 ( .A(n50709), .B(n42590), .Y(n31631) );
  XNOR2XL U35497 ( .A(n50706), .B(n42590), .Y(n31391) );
  XNOR2XL U35498 ( .A(n51347), .B(n42638), .Y(n31395) );
  XNOR2XL U35499 ( .A(n50774), .B(n36865), .Y(n29194) );
  XNOR2XL U35500 ( .A(n51412), .B(n36867), .Y(n29318) );
  XNOR2XL U35501 ( .A(n50770), .B(n34450), .Y(n29344) );
  XNOR2XL U35502 ( .A(n50775), .B(n34450), .Y(n29224) );
  XNOR2XL U35503 ( .A(n51409), .B(n36867), .Y(n29288) );
  XNOR2XL U35504 ( .A(n50771), .B(n42588), .Y(n29314) );
  XNOR2XL U35505 ( .A(n50768), .B(n36865), .Y(n29284) );
  XNOR2XL U35506 ( .A(n51410), .B(n42643), .Y(n29258) );
  XNOR2XL U35507 ( .A(n51407), .B(n36867), .Y(n29378) );
  XNOR2XL U35508 ( .A(n51408), .B(n42644), .Y(n29408) );
  XNOR2XL U35509 ( .A(n50769), .B(n42592), .Y(n29254) );
  XNOR2XL U35510 ( .A(n50766), .B(n36865), .Y(n29374) );
  XNOR2XL U35511 ( .A(n50767), .B(n42587), .Y(n29404) );
  XNOR2XL U35512 ( .A(n50573), .B(n36903), .Y(n27573) );
  XNOR2XL U35513 ( .A(n51177), .B(n42629), .Y(n26967) );
  XNOR2XL U35514 ( .A(n51173), .B(n42628), .Y(n27027) );
  XNOR2XL U35515 ( .A(n51168), .B(n42551), .Y(n25123) );
  XNOR2XL U35516 ( .A(n50536), .B(n36834), .Y(n26941) );
  XNOR2XL U35517 ( .A(n51166), .B(n41282), .Y(n25201) );
  XNOR2XL U35518 ( .A(n51166), .B(n42551), .Y(n24973) );
  XNOR2XL U35519 ( .A(n51179), .B(n41281), .Y(n26945) );
  XNOR2XL U35520 ( .A(n50523), .B(n41319), .Y(n25197) );
  XNOR2XL U35521 ( .A(n51213), .B(n42632), .Y(n27509) );
  XNOR2XL U35522 ( .A(n50520), .B(n36834), .Y(n24897) );
  XNOR2XL U35523 ( .A(n51144), .B(n42625), .Y(n28291) );
  XNOR2XL U35524 ( .A(n51176), .B(n42627), .Y(n26997) );
  XNOR2XL U35525 ( .A(n51163), .B(n41282), .Y(n24901) );
  XNOR2XL U35526 ( .A(n50503), .B(n42722), .Y(n28303) );
  XNOR2XL U35527 ( .A(n51207), .B(n41282), .Y(n27306) );
  XNOR2XL U35528 ( .A(n51207), .B(n42626), .Y(n27208) );
  XNOR2XL U35529 ( .A(n51211), .B(n42629), .Y(n27268) );
  XNOR2XL U35530 ( .A(n51224), .B(n41282), .Y(n27998) );
  XNOR2XL U35531 ( .A(n50532), .B(n36834), .Y(n27121) );
  XNOR2XL U35532 ( .A(n51175), .B(n41281), .Y(n27125) );
  XNOR2XL U35533 ( .A(n51179), .B(n42630), .Y(n26907) );
  XNOR2XL U35534 ( .A(n51153), .B(n42630), .Y(n28171) );
  XNOR2XL U35535 ( .A(n50581), .B(n36903), .Y(n27994) );
  XNOR2XL U35536 ( .A(n51204), .B(n42624), .Y(n27328) );
  XNOR2XL U35537 ( .A(n50512), .B(n42725), .Y(n28183) );
  XNOR2XL U35538 ( .A(n51160), .B(n42633), .Y(n24953) );
  XNOR2XL U35539 ( .A(n51164), .B(n41283), .Y(n24871) );
  XNOR2XL U35540 ( .A(n50535), .B(n36834), .Y(n26971) );
  XNOR2XL U35541 ( .A(n50580), .B(n42725), .Y(n28092) );
  XNOR2XL U35542 ( .A(n50531), .B(n36834), .Y(n27031) );
  XNOR2XL U35543 ( .A(n51174), .B(n41281), .Y(n27035) );
  XNOR2XL U35544 ( .A(n50571), .B(n36903), .Y(n27513) );
  XNOR2XL U35545 ( .A(n51178), .B(n41281), .Y(n26975) );
  XNOR2XL U35546 ( .A(n50785), .B(n36737), .Y(n27590) );
  XNOR2XL U35547 ( .A(n51212), .B(n41283), .Y(n27276) );
  XNOR2XL U35548 ( .A(n50779), .B(n42506), .Y(n27169) );
  XNOR2XL U35549 ( .A(n50502), .B(n41380), .Y(n28295) );
  XNOR2XL U35550 ( .A(n50534), .B(n36834), .Y(n27001) );
  XNOR2XL U35551 ( .A(n51177), .B(n41283), .Y(n27005) );
  XNOR2XL U35552 ( .A(n50569), .B(n36834), .Y(n27272) );
  XNOR2XL U35553 ( .A(n51161), .B(n42628), .Y(n24923) );
  XNOR2XL U35554 ( .A(n51183), .B(n41283), .Y(n26884) );
  XNOR2XL U35555 ( .A(n50737), .B(n36730), .Y(n25004) );
  XNOR2XL U35556 ( .A(n50565), .B(n36834), .Y(n27212) );
  XNOR2XL U35557 ( .A(n51208), .B(n41282), .Y(n27216) );
  XNOR2XL U35558 ( .A(n50537), .B(n41380), .Y(n26911) );
  XNOR2XL U35559 ( .A(n50735), .B(n36731), .Y(n25154) );
  XNOR2XL U35560 ( .A(n50511), .B(n42725), .Y(n28213) );
  XNOR2XL U35561 ( .A(n50511), .B(n41380), .Y(n28175) );
  XNOR2XL U35562 ( .A(n51438), .B(n42642), .Y(n27725) );
  XNOR2XL U35563 ( .A(n50562), .B(n36903), .Y(n27332) );
  XNOR2XL U35564 ( .A(n51205), .B(n41281), .Y(n27336) );
  XNOR2XL U35565 ( .A(n50579), .B(n41380), .Y(n28084) );
  XNOR2XL U35566 ( .A(n51161), .B(n41282), .Y(n24961) );
  XNOR2XL U35567 ( .A(n51152), .B(n34447), .Y(n28201) );
  XNOR2XL U35568 ( .A(n50754), .B(n42501), .Y(n26837) );
  XNOR2XL U35569 ( .A(n50793), .B(n36737), .Y(n28011) );
  XNOR2XL U35570 ( .A(n50751), .B(n42504), .Y(n26657) );
  XNOR2XL U35571 ( .A(n51172), .B(n42633), .Y(n27057) );
  XNOR2XL U35572 ( .A(n50786), .B(n36737), .Y(n27560) );
  XNOR2XL U35573 ( .A(n50552), .B(n42717), .Y(n29475) );
  XNOR2XL U35574 ( .A(n50726), .B(n42506), .Y(n28132) );
  XNOR2XL U35575 ( .A(n51151), .B(n42624), .Y(n28231) );
  XNOR2XL U35576 ( .A(n50513), .B(n36709), .Y(n28123) );
  XNOR2XL U35577 ( .A(n50510), .B(n42725), .Y(n28243) );
  XNOR2XL U35578 ( .A(n50504), .B(n36709), .Y(n28333) );
  XNOR2XL U35579 ( .A(n50519), .B(n36834), .Y(n24927) );
  XNOR2XL U35580 ( .A(n51181), .B(n34447), .Y(n26816) );
  XNOR2XL U35581 ( .A(n51154), .B(n42624), .Y(n28111) );
  XNOR2XL U35582 ( .A(n51145), .B(n42626), .Y(n28321) );
  XNOR2XL U35583 ( .A(n50758), .B(n42501), .Y(n26777) );
  XNOR2XL U35584 ( .A(n50781), .B(n42506), .Y(n27229) );
  XNOR2XL U35585 ( .A(n51171), .B(n42625), .Y(n25073) );
  XNOR2XL U35586 ( .A(n50577), .B(n36903), .Y(n27393) );
  XNOR2XL U35587 ( .A(n50516), .B(n41287), .Y(n24845) );
  XNOR2XL U35588 ( .A(n50510), .B(n41380), .Y(n28205) );
  XNOR2XL U35589 ( .A(n51170), .B(n42630), .Y(n25043) );
  XNOR2XL U35590 ( .A(n50780), .B(n42506), .Y(n27139) );
  XNOR2XL U35591 ( .A(n50784), .B(n36737), .Y(n27500) );
  XNOR2XL U35592 ( .A(n50530), .B(n36834), .Y(n27061) );
  XNOR2XL U35593 ( .A(n50736), .B(n36731), .Y(n25184) );
  XNOR2XL U35594 ( .A(n51173), .B(n41281), .Y(n27065) );
  XNOR2XL U35595 ( .A(n50789), .B(n36737), .Y(n27410) );
  XNOR2XL U35596 ( .A(n50509), .B(n41380), .Y(n28235) );
  XNOR2XL U35597 ( .A(n51182), .B(n41282), .Y(n26824) );
  XNOR2XL U35598 ( .A(n51141), .B(n42633), .Y(n28411) );
  XNOR2XL U35599 ( .A(n50512), .B(n41380), .Y(n28115) );
  XNOR2XL U35600 ( .A(n50503), .B(n41380), .Y(n28325) );
  XNOR2XL U35601 ( .A(n50499), .B(n36709), .Y(n28393) );
  XNOR2XL U35602 ( .A(n50755), .B(n42504), .Y(n26687) );
  XNOR2XL U35603 ( .A(n51193), .B(n42628), .Y(n29463) );
  XNOR2XL U35604 ( .A(n50529), .B(n36834), .Y(n25077) );
  XNOR2XL U35605 ( .A(n50749), .B(n42508), .Y(n26928) );
  XNOR2XL U35606 ( .A(n51172), .B(n41283), .Y(n25081) );
  XNOR2XL U35607 ( .A(n50506), .B(n36709), .Y(n28273) );
  XNOR2XL U35608 ( .A(n51171), .B(n41282), .Y(n25051) );
  XNOR2XL U35609 ( .A(n50777), .B(n42506), .Y(n27289) );
  XNOR2XL U35610 ( .A(n50528), .B(n36905), .Y(n25047) );
  XNOR2XL U35611 ( .A(n51205), .B(n42626), .Y(n27358) );
  XNOR2XL U35612 ( .A(n50748), .B(n42506), .Y(n26958) );
  XNOR2XL U35613 ( .A(n51157), .B(n42626), .Y(n24833) );
  XNOR2XL U35614 ( .A(n51147), .B(n42631), .Y(n28261) );
  XNOR2XL U35615 ( .A(n50733), .B(n42505), .Y(n24884) );
  XNOR2XL U35616 ( .A(n50778), .B(n42506), .Y(n27199) );
  XNOR2XL U35617 ( .A(n50499), .B(n41380), .Y(n28415) );
  XNOR2XL U35618 ( .A(n50782), .B(n36737), .Y(n27259) );
  XNOR2XL U35619 ( .A(n50753), .B(n42506), .Y(n26867) );
  XNOR2XL U35620 ( .A(n50747), .B(n42506), .Y(n26988) );
  XNOR2XL U35621 ( .A(n50745), .B(n42506), .Y(n27108) );
  XNOR2XL U35622 ( .A(n50792), .B(n36737), .Y(n28071) );
  XNOR2XL U35623 ( .A(n51175), .B(n42629), .Y(n27087) );
  XNOR2XL U35624 ( .A(n50551), .B(n36728), .Y(n29467) );
  XNOR2XL U35625 ( .A(n50775), .B(n36737), .Y(n27319) );
  XNOR2XL U35626 ( .A(n50760), .B(n42501), .Y(n29033) );
  XNOR2XL U35627 ( .A(n50744), .B(n42506), .Y(n27018) );
  XNOR2XL U35628 ( .A(n51206), .B(n41281), .Y(n27366) );
  XNOR2XL U35629 ( .A(n50563), .B(n36903), .Y(n27362) );
  XNOR2XL U35630 ( .A(n50505), .B(n41380), .Y(n28265) );
  XNOR2XL U35631 ( .A(n50731), .B(n36731), .Y(n24944) );
  XNOR2XL U35632 ( .A(n50761), .B(n42501), .Y(n29093) );
  XNOR2XL U35633 ( .A(n50767), .B(n42502), .Y(n29274) );
  XNOR2XL U35634 ( .A(n51158), .B(n41283), .Y(n24841) );
  XNOR2XL U35635 ( .A(n50732), .B(n42505), .Y(n24914) );
  XNOR2XL U35636 ( .A(n51146), .B(n42632), .Y(n28351) );
  XNOR2XL U35637 ( .A(n50505), .B(n41287), .Y(n28363) );
  XNOR2XL U35638 ( .A(n51176), .B(n41282), .Y(n27095) );
  XNOR2XL U35639 ( .A(n50752), .B(n42504), .Y(n26807) );
  XNOR2XL U35640 ( .A(n50533), .B(n36834), .Y(n27091) );
  XNOR2XL U35641 ( .A(n50727), .B(n42505), .Y(n24794) );
  XNOR2XL U35642 ( .A(n50763), .B(n42502), .Y(n29424) );
  XNOR2XL U35643 ( .A(n50790), .B(n36737), .Y(n27380) );
  XNOR2XL U35644 ( .A(n50750), .B(n42504), .Y(n26898) );
  XNOR2XL U35645 ( .A(n50715), .B(n42501), .Y(n28282) );
  XNOR2XL U35646 ( .A(n50742), .B(n36731), .Y(n25064) );
  XNOR2XL U35647 ( .A(n50496), .B(n36875), .Y(n31642) );
  XNOR2XL U35648 ( .A(n50743), .B(n42506), .Y(n27048) );
  XNOR2XL U35649 ( .A(n50741), .B(n36730), .Y(n25034) );
  XNOR2XL U35650 ( .A(n50768), .B(n42502), .Y(n29244) );
  XNOR2XL U35651 ( .A(n50766), .B(n42502), .Y(n29394) );
  XNOR2XL U35652 ( .A(n50729), .B(n42505), .Y(n24734) );
  XNOR2XL U35653 ( .A(n50730), .B(n42505), .Y(n24764) );
  XNOR2XL U35654 ( .A(n50504), .B(n41380), .Y(n28355) );
  XNOR2XL U35655 ( .A(n50759), .B(n42501), .Y(n29003) );
  XNOR2XL U35656 ( .A(n50494), .B(n42718), .Y(n31402) );
  XNOR2XL U35657 ( .A(n50776), .B(n36737), .Y(n27349) );
  XNOR2XL U35658 ( .A(n50765), .B(n42502), .Y(n29364) );
  XNOR2XL U35659 ( .A(n50728), .B(n42505), .Y(n24824) );
  XNOR2XL U35660 ( .A(n50746), .B(n42506), .Y(n27078) );
  XNOR2XL U35661 ( .A(n51137), .B(n42625), .Y(n31630) );
  XNOR2XL U35662 ( .A(n51134), .B(n42628), .Y(n31390) );
  XNOR2XL U35663 ( .A(n50764), .B(n42502), .Y(n29454) );
  XNOR2XL U35664 ( .A(n50722), .B(n42501), .Y(n28222) );
  XNOR2XL U35665 ( .A(n50712), .B(n42501), .Y(n28402) );
  XNOR2XL U35666 ( .A(n50718), .B(n42501), .Y(n28252) );
  XNOR2XL U35667 ( .A(n50719), .B(n42501), .Y(n28522) );
  XNOR2XL U35668 ( .A(n50493), .B(n41380), .Y(n31394) );
  XNOR2XL U35669 ( .A(n50495), .B(n41380), .Y(n31634) );
  XNOR2XL U35670 ( .A(n51154), .B(n41332), .Y(n23224) );
  XNOR2XL U35671 ( .A(n51150), .B(n41329), .Y(n23275) );
  XNOR2XL U35672 ( .A(n51151), .B(n41328), .Y(n23234) );
  XNOR2XL U35673 ( .A(n51149), .B(n41331), .Y(n23264) );
  XNOR2XL U35674 ( .A(n50561), .B(n41319), .Y(n29227) );
  XNOR2XL U35675 ( .A(n50557), .B(n36905), .Y(n29317) );
  XNOR2XL U35676 ( .A(n50554), .B(n41379), .Y(n29287) );
  XNOR2XL U35677 ( .A(n50548), .B(n41379), .Y(n29106) );
  XNOR2XL U35678 ( .A(n50555), .B(n36903), .Y(n29257) );
  XNOR2XL U35679 ( .A(n50552), .B(n41319), .Y(n29377) );
  XNOR2XL U35680 ( .A(n50553), .B(n36903), .Y(n29407) );
  XNOR2XL U35681 ( .A(n51203), .B(n42629), .Y(n29223) );
  XNOR2XL U35682 ( .A(n51199), .B(n42624), .Y(n29313) );
  XNOR2XL U35683 ( .A(n51196), .B(n42628), .Y(n29283) );
  XNOR2XL U35684 ( .A(n51197), .B(n42633), .Y(n29253) );
  XNOR2XL U35685 ( .A(n51194), .B(n42632), .Y(n29373) );
  XNOR2XL U35686 ( .A(n51195), .B(n42625), .Y(n29403) );
  XNOR2XL U35687 ( .A(n50726), .B(n36851), .Y(n23225) );
  XNOR2XL U35688 ( .A(n50722), .B(n36853), .Y(n23276) );
  XNOR2XL U35689 ( .A(n50723), .B(n36856), .Y(n23235) );
  XNOR2XL U35690 ( .A(n50721), .B(n36858), .Y(n23265) );
  XNOR2XL U35691 ( .A(n50723), .B(n36731), .Y(n28192) );
  XNOR2XL U35692 ( .A(n50716), .B(n36730), .Y(n28312) );
  XNOR2XL U35693 ( .A(n50721), .B(n36731), .Y(n28492) );
  XNOR2XL U35694 ( .A(n50711), .B(n36730), .Y(n28372) );
  XNOR2XL U35695 ( .A(n51198), .B(n41283), .Y(n29261) );
  XNOR2XL U35696 ( .A(n50770), .B(net219468), .Y(n29262) );
  XNOR2XL U35697 ( .A(n50932), .B(net219310), .Y(n28328) );
  XNOR2XL U35698 ( .A(n51146), .B(n41282), .Y(n28329) );
  XNOR2XL U35699 ( .A(n50718), .B(net219468), .Y(n28330) );
  XNOR2XL U35700 ( .A(n50980), .B(net219308), .Y(n29470) );
  XNOR2XL U35701 ( .A(n51194), .B(n41283), .Y(n29471) );
  XNOR2XL U35702 ( .A(n50766), .B(net219450), .Y(n29472) );
  XNOR2XL U35703 ( .A(n50934), .B(net219310), .Y(n28268) );
  XNOR2XL U35704 ( .A(n51148), .B(n41283), .Y(n28269) );
  XNOR2XL U35705 ( .A(n50720), .B(net219468), .Y(n28270) );
  NOR4X2 U35706 ( .A(n31547), .B(n31548), .C(n31549), .D(n31550), .Y(n43220)
         );
  XNOR2XL U35707 ( .A(n50712), .B(net219450), .Y(n31579) );
  XNOR2XL U35708 ( .A(n50922), .B(net219310), .Y(n31367) );
  XNOR2XL U35709 ( .A(n51136), .B(n41282), .Y(n31368) );
  XNOR2XL U35710 ( .A(n50708), .B(net219450), .Y(n31369) );
  XNOR2XL U35711 ( .A(n50928), .B(net219310), .Y(n28418) );
  XNOR2XL U35712 ( .A(n51142), .B(n41283), .Y(n28419) );
  XNOR2XL U35713 ( .A(n50714), .B(net219468), .Y(n28420) );
  XNOR2XL U35714 ( .A(n50930), .B(net219330), .Y(n28478) );
  XNOR2XL U35715 ( .A(n51144), .B(n41281), .Y(n28479) );
  XNOR2XL U35716 ( .A(n50716), .B(net219468), .Y(n28480) );
  XOR2XL U35717 ( .A(n42084), .B(n41321), .Y(n44876) );
  XOR2XL U35718 ( .A(n42091), .B(n41323), .Y(n44725) );
  XOR2XL U35719 ( .A(n42083), .B(n41321), .Y(n45339) );
  XOR2XL U35720 ( .A(n42079), .B(n36873), .Y(n45515) );
  XOR2XL U35721 ( .A(n42078), .B(n36877), .Y(n45488) );
  XNOR2XL U35722 ( .A(n51355), .B(n42702), .Y(n28424) );
  XNOR2XL U35723 ( .A(n51356), .B(n42701), .Y(n28454) );
  XNOR2XL U35724 ( .A(n51363), .B(n42698), .Y(n28574) );
  XNOR2XL U35725 ( .A(n51364), .B(n42701), .Y(n28514) );
  XNOR2XL U35726 ( .A(n51362), .B(n42702), .Y(n28544) );
  XNOR2XL U35727 ( .A(n51357), .B(n42701), .Y(n28484) );
  XOR2XL U35728 ( .A(n42103), .B(n36877), .Y(n27683) );
  XOR2XL U35729 ( .A(n42112), .B(n36801), .Y(n27562) );
  XOR2XL U35730 ( .A(n42102), .B(n41321), .Y(n27713) );
  XOR2XL U35731 ( .A(n42114), .B(n36873), .Y(n27502) );
  XOR2XL U35732 ( .A(n42104), .B(n36873), .Y(n27983) );
  XOR2XL U35733 ( .A(n42123), .B(n36877), .Y(n27321) );
  XOR2XL U35734 ( .A(n42108), .B(n36877), .Y(n27382) );
  XOR2XL U35735 ( .A(n42184), .B(n36815), .Y(n23187) );
  XOR2XL U35736 ( .A(n42101), .B(n42493), .Y(n20412) );
  XOR2XL U35737 ( .A(n42183), .B(n36817), .Y(n23147) );
  XOR2XL U35738 ( .A(n42180), .B(n36813), .Y(n23127) );
  XNOR2XL U35739 ( .A(n50344), .B(n42707), .Y(n29053) );
  XNOR2XL U35740 ( .A(n50296), .B(n42707), .Y(n28422) );
  XNOR2XL U35741 ( .A(n50297), .B(n42707), .Y(n28452) );
  XNOR2XL U35742 ( .A(n50304), .B(n42709), .Y(n28572) );
  XNOR2XL U35743 ( .A(n50305), .B(n42707), .Y(n28512) );
  XNOR2XL U35744 ( .A(n50303), .B(n42707), .Y(n28542) );
  XNOR2XL U35745 ( .A(n50298), .B(n42707), .Y(n28482) );
  XOR2XL U35746 ( .A(n42103), .B(n36815), .Y(n23808) );
  XOR2XL U35747 ( .A(n42119), .B(n36814), .Y(n23707) );
  XOR2XL U35748 ( .A(n42120), .B(n36810), .Y(n23717) );
  XOR2XL U35749 ( .A(n42106), .B(n36810), .Y(n23848) );
  XOR2XL U35750 ( .A(n42164), .B(n36816), .Y(n23594) );
  XOR2XL U35751 ( .A(n42101), .B(n36809), .Y(n23788) );
  XOR2XL U35752 ( .A(n42105), .B(n36814), .Y(n23858) );
  XOR2XL U35753 ( .A(n42138), .B(n36808), .Y(n22350) );
  XOR2XL U35754 ( .A(n42112), .B(n36815), .Y(n23938) );
  XOR2XL U35755 ( .A(n42121), .B(n36817), .Y(n23767) );
  XOR2XL U35756 ( .A(n42117), .B(n36808), .Y(n23747) );
  XOR2XL U35757 ( .A(n42118), .B(n36817), .Y(n23737) );
  XOR2XL U35758 ( .A(n42114), .B(n36815), .Y(n24008) );
  XOR2XL U35759 ( .A(n42107), .B(n36813), .Y(n23838) );
  XOR2XL U35760 ( .A(n42115), .B(n36817), .Y(n23988) );
  XOR2XL U35761 ( .A(n42108), .B(n36817), .Y(n23978) );
  XOR2XL U35762 ( .A(n42126), .B(n36808), .Y(n22450) );
  XOR2XL U35763 ( .A(n42110), .B(n36817), .Y(n23958) );
  XOR2XL U35764 ( .A(n42122), .B(n36811), .Y(n23697) );
  XOR2XL U35765 ( .A(n42125), .B(n36807), .Y(n22460) );
  XOR2XL U35766 ( .A(n42124), .B(n36809), .Y(n22470) );
  XOR2XL U35767 ( .A(n42147), .B(n36814), .Y(n24019) );
  XOR2XL U35768 ( .A(n42150), .B(n36808), .Y(n24110) );
  XOR2XL U35769 ( .A(n42152), .B(n36811), .Y(n24151) );
  XOR2XL U35770 ( .A(n42149), .B(n36815), .Y(n24120) );
  XOR2XL U35771 ( .A(n42139), .B(n36808), .Y(n22320) );
  XOR2XL U35772 ( .A(n42154), .B(n36810), .Y(n24140) );
  XOR2XL U35773 ( .A(n42142), .B(n36808), .Y(n24039) );
  XOR2XL U35774 ( .A(n42155), .B(n36817), .Y(n24161) );
  XOR2XL U35775 ( .A(n42132), .B(n36811), .Y(n22360) );
  XOR2XL U35776 ( .A(n42168), .B(n36814), .Y(n23472) );
  XOR2XL U35777 ( .A(n42143), .B(n36808), .Y(n24029) );
  XOR2XL U35778 ( .A(n42111), .B(n36817), .Y(n23948) );
  XOR2XL U35779 ( .A(n42133), .B(n36814), .Y(n22370) );
  XOR2XL U35780 ( .A(n42123), .B(n36814), .Y(n23727) );
  XOR2XL U35781 ( .A(n42140), .B(n36816), .Y(n24059) );
  XOR2XL U35782 ( .A(n42166), .B(n36807), .Y(n23572) );
  XOR2XL U35783 ( .A(n42109), .B(n36807), .Y(n23968) );
  XOR2XL U35784 ( .A(n42141), .B(n36810), .Y(n24049) );
  XOR2XL U35785 ( .A(n42158), .B(n36810), .Y(n23532) );
  XOR2XL U35786 ( .A(n42129), .B(n42480), .Y(n19537) );
  XOR2XL U35787 ( .A(n42165), .B(n36816), .Y(n23583) );
  XOR2XL U35788 ( .A(n42120), .B(n42492), .Y(n20115) );
  XOR2XL U35789 ( .A(n42156), .B(n36813), .Y(n235520) );
  XOR2XL U35790 ( .A(n42163), .B(n36813), .Y(n23492) );
  XOR2XL U35791 ( .A(n42144), .B(n36815), .Y(n24079) );
  XOR2XL U35792 ( .A(n42104), .B(n42479), .Y(n20290) );
  XOR2XL U35793 ( .A(n42136), .B(n36813), .Y(n22340) );
  XOR2XL U35794 ( .A(n42134), .B(n36809), .Y(n22380) );
  XOR2XL U35795 ( .A(n42105), .B(n42480), .Y(n20300) );
  XNOR2XL U35796 ( .A(n50507), .B(n42584), .Y(n28495) );
  XNOR2XL U35797 ( .A(n50505), .B(n42584), .Y(n28525) );
  XNOR2XL U35798 ( .A(n50497), .B(n42584), .Y(n28375) );
  XNOR2XL U35799 ( .A(n50499), .B(n42584), .Y(n28435) );
  XNOR2XL U35800 ( .A(n50343), .B(n36907), .Y(n29045) );
  XNOR2XL U35801 ( .A(n50342), .B(n36907), .Y(n29015) );
  XNOR2XL U35802 ( .A(n50926), .B(n42620), .Y(n28380) );
  XNOR2XL U35803 ( .A(n50935), .B(n42620), .Y(n28560) );
  XNOR2XL U35804 ( .A(n50296), .B(n36907), .Y(n28444) );
  XNOR2XL U35805 ( .A(n50934), .B(n42620), .Y(n28530) );
  XNOR2XL U35806 ( .A(n50294), .B(n36907), .Y(n28384) );
  XNOR2XL U35807 ( .A(n50303), .B(n36907), .Y(n28564) );
  XNOR2XL U35808 ( .A(n50304), .B(n36907), .Y(n28504) );
  XNOR2XL U35809 ( .A(n50929), .B(n42620), .Y(n28470) );
  XNOR2XL U35810 ( .A(n50302), .B(n36907), .Y(n28534) );
  XNOR2XL U35811 ( .A(n50297), .B(n36907), .Y(n28474) );
  XNOR2XL U35812 ( .A(n50526), .B(n42580), .Y(n25127) );
  XNOR2XL U35813 ( .A(n50524), .B(n42580), .Y(n24977) );
  XNOR2XL U35814 ( .A(n51009), .B(n42542), .Y(n27679) );
  XNOR2XL U35815 ( .A(n50379), .B(n42675), .Y(n27723) );
  XNOR2XL U35816 ( .A(n50999), .B(n42542), .Y(n27588) );
  XNOR2XL U35817 ( .A(n50951), .B(n42539), .Y(n25002) );
  XNOR2XL U35818 ( .A(n50949), .B(n42539), .Y(n25152) );
  XNOR2XL U35819 ( .A(n51007), .B(n42543), .Y(n28009) );
  XNOR2XL U35820 ( .A(n50965), .B(n42540), .Y(n26655) );
  XNOR2XL U35821 ( .A(n50968), .B(n42540), .Y(n26835) );
  XNOR2XL U35822 ( .A(n51000), .B(n42542), .Y(n27558) );
  XNOR2XL U35823 ( .A(n51010), .B(n42542), .Y(n27709) );
  XNOR2XL U35824 ( .A(n51005), .B(n42543), .Y(n28039) );
  XNOR2XL U35825 ( .A(n50972), .B(n42540), .Y(n26775) );
  XNOR2XL U35826 ( .A(n50994), .B(n42541), .Y(n27137) );
  XNOR2XL U35827 ( .A(n50998), .B(n42542), .Y(n27498) );
  XNOR2XL U35828 ( .A(n51003), .B(n42542), .Y(n27408) );
  XNOR2XL U35829 ( .A(n50950), .B(n42539), .Y(n25182) );
  XNOR2XL U35830 ( .A(n50969), .B(n42540), .Y(n26685) );
  XNOR2XL U35831 ( .A(n51008), .B(n42542), .Y(n27979) );
  XNOR2XL U35832 ( .A(n50963), .B(n42541), .Y(n26926) );
  XNOR2XL U35833 ( .A(n50991), .B(n42541), .Y(n27287) );
  XNOR2XL U35834 ( .A(n50962), .B(n42541), .Y(n26956) );
  XNOR2XL U35835 ( .A(n50948), .B(n42536), .Y(n24852) );
  XNOR2XL U35836 ( .A(n50947), .B(n42539), .Y(n24882) );
  XNOR2XL U35837 ( .A(n50983), .B(n42535), .Y(n29332) );
  XNOR2XL U35838 ( .A(n50992), .B(n42541), .Y(n27197) );
  XNOR2XL U35839 ( .A(n50961), .B(n42541), .Y(n26986) );
  XNOR2XL U35840 ( .A(n50996), .B(n42541), .Y(n27257) );
  XNOR2XL U35841 ( .A(n50959), .B(n42541), .Y(n27106) );
  XNOR2XL U35842 ( .A(n50967), .B(n42540), .Y(n26865) );
  XNOR2XL U35843 ( .A(n51006), .B(n42543), .Y(n28069) );
  XNOR2XL U35844 ( .A(n50989), .B(n42542), .Y(n27317) );
  XNOR2XL U35845 ( .A(n50958), .B(n42541), .Y(n27016) );
  XNOR2XL U35846 ( .A(n50937), .B(n42543), .Y(n28190) );
  XNOR2XL U35847 ( .A(n50929), .B(n42543), .Y(n28280) );
  XNOR2XL U35848 ( .A(n50945), .B(n42539), .Y(n24942) );
  XNOR2XL U35849 ( .A(n50981), .B(n42535), .Y(n29272) );
  XNOR2XL U35850 ( .A(n50946), .B(n42539), .Y(n24912) );
  XNOR2XL U35851 ( .A(n50939), .B(n42543), .Y(n28100) );
  XNOR2XL U35852 ( .A(n50938), .B(n42543), .Y(n28160) );
  XNOR2XL U35853 ( .A(n50977), .B(n42535), .Y(n29422) );
  XNOR2XL U35854 ( .A(n51004), .B(n42542), .Y(n27378) );
  XNOR2XL U35855 ( .A(n50966), .B(n42540), .Y(n26805) );
  XNOR2XL U35856 ( .A(n50956), .B(n42539), .Y(n25062) );
  XNOR2XL U35857 ( .A(n50957), .B(n42541), .Y(n27046) );
  XNOR2XL U35858 ( .A(n50964), .B(n42540), .Y(n26896) );
  XNOR2XL U35859 ( .A(n50955), .B(n42539), .Y(n25032) );
  XNOR2XL U35860 ( .A(n50982), .B(n42535), .Y(n29242) );
  XNOR2XL U35861 ( .A(n50980), .B(n42535), .Y(n29392) );
  XNOR2XL U35862 ( .A(n50941), .B(n42536), .Y(n24792) );
  XNOR2XL U35863 ( .A(n50930), .B(n42543), .Y(n28310) );
  XNOR2XL U35864 ( .A(n50990), .B(n42542), .Y(n27347) );
  XNOR2XL U35865 ( .A(n50943), .B(n42543), .Y(n24732) );
  XNOR2XL U35866 ( .A(n50979), .B(n42535), .Y(n29362) );
  XNOR2XL U35867 ( .A(n50936), .B(n42543), .Y(n28220) );
  XNOR2XL U35868 ( .A(n50944), .B(n42544), .Y(n24762) );
  XNOR2XL U35869 ( .A(n50926), .B(n42543), .Y(n28400) );
  XNOR2XL U35870 ( .A(n50932), .B(n42543), .Y(n28250) );
  XNOR2XL U35871 ( .A(n50960), .B(n42541), .Y(n27076) );
  XNOR2XL U35872 ( .A(n50978), .B(n42535), .Y(n29452) );
  XNOR2XL U35873 ( .A(n50942), .B(n42541), .Y(n24822) );
  XNOR2XL U35874 ( .A(n50940), .B(n41291), .Y(n23223) );
  XNOR2XL U35875 ( .A(n50936), .B(n41293), .Y(n23274) );
  XNOR2XL U35876 ( .A(n50937), .B(n41293), .Y(n23233) );
  XNOR2XL U35877 ( .A(n50935), .B(n36916), .Y(n23263) );
  XNOR2XL U35878 ( .A(n50973), .B(n42534), .Y(n29001) );
  XNOR2XL U35879 ( .A(n50547), .B(n42725), .Y(n29024) );
  XNOR2XL U35880 ( .A(n50500), .B(n42725), .Y(n28423) );
  XNOR2XL U35881 ( .A(n50501), .B(n42725), .Y(n28453) );
  XNOR2XL U35882 ( .A(n50508), .B(n42725), .Y(n28573) );
  XNOR2XL U35883 ( .A(n50509), .B(n42725), .Y(n28513) );
  XNOR2XL U35884 ( .A(n50507), .B(n42725), .Y(n28543) );
  XNOR2XL U35885 ( .A(n50502), .B(n42725), .Y(n28483) );
  XNOR2XL U35886 ( .A(n50513), .B(n42579), .Y(n24797) );
  XNOR2XL U35887 ( .A(n50516), .B(n42579), .Y(n24767) );
  XNOR2XL U35888 ( .A(n50515), .B(n42579), .Y(n24737) );
  XNOR2XL U35889 ( .A(n50514), .B(n42579), .Y(n24827) );
  XNOR2XL U35890 ( .A(n50714), .B(n42592), .Y(n28442) );
  XNOR2XL U35891 ( .A(n50712), .B(n42592), .Y(n28382) );
  XNOR2XL U35892 ( .A(n50721), .B(n42592), .Y(n28562) );
  XNOR2XL U35893 ( .A(n50763), .B(n42592), .Y(n29073) );
  XNOR2XL U35894 ( .A(n50722), .B(n42592), .Y(n28502) );
  XNOR2XL U35895 ( .A(n50720), .B(n42592), .Y(n28532) );
  XNOR2XL U35896 ( .A(n50715), .B(n42592), .Y(n28472) );
  XNOR2XL U35897 ( .A(n50546), .B(n36905), .Y(n29016) );
  XNOR2XL U35898 ( .A(n50500), .B(n36905), .Y(n28445) );
  XNOR2XL U35899 ( .A(n50498), .B(n36903), .Y(n28385) );
  XNOR2XL U35900 ( .A(n50507), .B(n36728), .Y(n28565) );
  XNOR2XL U35901 ( .A(n50508), .B(n36905), .Y(n28505) );
  XNOR2XL U35902 ( .A(n50506), .B(n41380), .Y(n28535) );
  XNOR2XL U35903 ( .A(n50501), .B(n36903), .Y(n28475) );
  XNOR2XL U35904 ( .A(n51142), .B(n42628), .Y(n28441) );
  XNOR2XL U35905 ( .A(n51140), .B(n42627), .Y(n28381) );
  XNOR2XL U35906 ( .A(n51149), .B(n42628), .Y(n28561) );
  XNOR2XL U35907 ( .A(n51191), .B(n42626), .Y(n29072) );
  XNOR2XL U35908 ( .A(n51150), .B(n42628), .Y(n28501) );
  XNOR2XL U35909 ( .A(n51148), .B(n42627), .Y(n28531) );
  XNOR2XL U35910 ( .A(n51143), .B(n42624), .Y(n28471) );
  XOR2XL U35911 ( .A(n42172), .B(n36816), .Y(n23227) );
  XOR2XL U35912 ( .A(n42176), .B(n36809), .Y(n23278) );
  XOR2XL U35913 ( .A(n42175), .B(n36814), .Y(n23237) );
  XNOR2XL U35914 ( .A(n51435), .B(n41300), .Y(n23819) );
  XNOR2XL U35915 ( .A(n51436), .B(n41305), .Y(n23809) );
  XNOR2XL U35916 ( .A(n51433), .B(n41301), .Y(n23849) );
  XNOR2XL U35917 ( .A(n51438), .B(n41302), .Y(n23789) );
  XNOR2XL U35918 ( .A(n50533), .B(n36779), .Y(n24101) );
  XNOR2XL U35919 ( .A(n51434), .B(n41299), .Y(n23859) );
  XNOR2XL U35920 ( .A(n51427), .B(n41302), .Y(n23939) );
  XNOR2XL U35921 ( .A(n51425), .B(n41302), .Y(n24009) );
  XNOR2XL U35922 ( .A(n50563), .B(n36780), .Y(n23768) );
  XNOR2XL U35923 ( .A(n51426), .B(n41299), .Y(n23999) );
  XNOR2XL U35924 ( .A(n50566), .B(n36783), .Y(n23738) );
  XNOR2XL U35925 ( .A(n50567), .B(n36778), .Y(n23748) );
  XNOR2XL U35926 ( .A(n51424), .B(n41302), .Y(n23989) );
  XNOR2XL U35927 ( .A(n51429), .B(n41301), .Y(n23959) );
  XNOR2XL U35928 ( .A(n50577), .B(n36780), .Y(n23839) );
  XNOR2XL U35929 ( .A(n51437), .B(n41305), .Y(n23779) );
  XNOR2XL U35930 ( .A(n50576), .B(n36779), .Y(n23979) );
  XNOR2XL U35931 ( .A(n51365), .B(n41305), .Y(n23208) );
  XNOR2XL U35932 ( .A(n50562), .B(n36786), .Y(n23698) );
  XNOR2XL U35933 ( .A(n51392), .B(n41300), .Y(n24020) );
  XNOR2XL U35934 ( .A(n51372), .B(n41301), .Y(n23605) );
  XNOR2XL U35935 ( .A(n51410), .B(n41299), .Y(n22411) );
  XNOR2XL U35936 ( .A(n51363), .B(n41303), .Y(n23279) );
  XNOR2XL U35937 ( .A(n50534), .B(n36785), .Y(n24111) );
  XNOR2XL U35938 ( .A(n50532), .B(n36783), .Y(n24152) );
  XNOR2XL U35939 ( .A(n51397), .B(n36918), .Y(n24040) );
  XNOR2XL U35940 ( .A(n50535), .B(n36784), .Y(n24121) );
  XNOR2XL U35941 ( .A(n51371), .B(n41305), .Y(n23473) );
  XNOR2XL U35942 ( .A(n50530), .B(n36782), .Y(n24142) );
  XNOR2XL U35943 ( .A(n51396), .B(n41299), .Y(n24030) );
  XNOR2XL U35944 ( .A(n51428), .B(n41305), .Y(n23949) );
  XNOR2XL U35945 ( .A(n51373), .B(n36918), .Y(n23574) );
  XNOR2XL U35946 ( .A(n51398), .B(n41304), .Y(n24050) );
  XNOR2XL U35947 ( .A(n50501), .B(n36776), .Y(n23148) );
  XNOR2XL U35948 ( .A(n50564), .B(n36771), .Y(n20117) );
  XNOR2XL U35949 ( .A(n51430), .B(n41301), .Y(n23969) );
  XNOR2XL U35950 ( .A(n50561), .B(n36777), .Y(n23728) );
  XNOR2XL U35951 ( .A(n50544), .B(n36783), .Y(n24060) );
  XNOR2XL U35952 ( .A(n51381), .B(n41302), .Y(n23533) );
  XNOR2XL U35953 ( .A(n51374), .B(n41302), .Y(n23585) );
  XNOR2XL U35954 ( .A(n51435), .B(n36740), .Y(n20291) );
  XNOR2XL U35955 ( .A(n51376), .B(n41300), .Y(n23493) );
  XNOR2XL U35956 ( .A(n51395), .B(n41299), .Y(n24080) );
  XNOR2XL U35957 ( .A(n51434), .B(n36742), .Y(n20301) );
  XNOR2XL U35958 ( .A(n51364), .B(n41300), .Y(n23238) );
  XNOR2XL U35959 ( .A(n50512), .B(n36784), .Y(n23228) );
  XNOR2XL U35960 ( .A(n50504), .B(n36778), .Y(n23128) );
  XNOR2XL U35961 ( .A(n51375), .B(n36871), .Y(n24936) );
  XNOR2XL U35962 ( .A(n51373), .B(n42695), .Y(n24786) );
  XNOR2XL U35963 ( .A(n50325), .B(n42707), .Y(n25054) );
  XNOR2XL U35964 ( .A(n50529), .B(n36709), .Y(n25055) );
  XNOR2XL U35965 ( .A(n51384), .B(n42697), .Y(n25056) );
  XNOR2XL U35966 ( .A(n50311), .B(n42672), .Y(n24836) );
  XNOR2XL U35967 ( .A(n50515), .B(n36905), .Y(n24837) );
  XNOR2XL U35968 ( .A(n51370), .B(n42641), .Y(n24838) );
  XNOR2XL U35969 ( .A(n50569), .B(n42582), .Y(n27533) );
  XNOR2XL U35970 ( .A(n50581), .B(n42582), .Y(n27684) );
  XNOR2XL U35971 ( .A(n50571), .B(n42582), .Y(n27593) );
  XNOR2XL U35972 ( .A(n50986), .B(n42535), .Y(n29152) );
  XNOR2XL U35973 ( .A(n50523), .B(n42580), .Y(n25007) );
  XNOR2XL U35974 ( .A(n50521), .B(n42580), .Y(n25157) );
  XNOR2XL U35975 ( .A(n50540), .B(n42576), .Y(n26840) );
  XNOR2XL U35976 ( .A(n50987), .B(n42535), .Y(n29182) );
  XNOR2XL U35977 ( .A(n50572), .B(n42582), .Y(n27563) );
  XNOR2XL U35978 ( .A(n50579), .B(n42583), .Y(n28014) );
  XNOR2XL U35979 ( .A(n50582), .B(n42582), .Y(n27714) );
  XNOR2XL U35980 ( .A(n50537), .B(n42576), .Y(n26660) );
  XNOR2XL U35981 ( .A(n50544), .B(n42576), .Y(n26780) );
  XNOR2XL U35982 ( .A(n50566), .B(n42581), .Y(n27142) );
  XNOR2XL U35983 ( .A(n50570), .B(n42582), .Y(n27503) );
  XNOR2XL U35984 ( .A(n50522), .B(n42580), .Y(n25187) );
  XNOR2XL U35985 ( .A(n50577), .B(n42583), .Y(n28044) );
  XNOR2XL U35986 ( .A(n50575), .B(n42582), .Y(n27413) );
  XNOR2XL U35987 ( .A(n50580), .B(n42582), .Y(n27984) );
  XNOR2XL U35988 ( .A(n50556), .B(n42577), .Y(n29307) );
  XNOR2XL U35989 ( .A(n50541), .B(n42576), .Y(n26690) );
  XNOR2XL U35990 ( .A(n50534), .B(n42581), .Y(n26961) );
  XNOR2XL U35991 ( .A(n50535), .B(n42581), .Y(n26931) );
  XNOR2XL U35992 ( .A(n50564), .B(n42581), .Y(n27202) );
  XNOR2XL U35993 ( .A(n50568), .B(n42581), .Y(n27262) );
  XNOR2XL U35994 ( .A(n50519), .B(n42580), .Y(n24887) );
  XNOR2XL U35995 ( .A(n50555), .B(n42577), .Y(n29337) );
  XNOR2XL U35996 ( .A(n50578), .B(n42583), .Y(n28074) );
  XNOR2XL U35997 ( .A(n50531), .B(n42581), .Y(n27111) );
  XNOR2XL U35998 ( .A(n50533), .B(n42581), .Y(n26991) );
  XNOR2XL U35999 ( .A(n50509), .B(n42583), .Y(n28195) );
  XNOR2XL U36000 ( .A(n50539), .B(n42576), .Y(n26870) );
  XNOR2XL U36001 ( .A(n50530), .B(n42581), .Y(n27021) );
  XNOR2XL U36002 ( .A(n50561), .B(n42582), .Y(n27322) );
  XNOR2XL U36003 ( .A(n50518), .B(n42580), .Y(n24917) );
  XNOR2XL U36004 ( .A(n50501), .B(n42583), .Y(n28285) );
  XNOR2XL U36005 ( .A(n50517), .B(n42580), .Y(n24947) );
  XNOR2XL U36006 ( .A(n50511), .B(n42583), .Y(n28105) );
  XNOR2XL U36007 ( .A(n50553), .B(n42577), .Y(n29277) );
  XNOR2XL U36008 ( .A(n50538), .B(n42576), .Y(n26810) );
  XNOR2XL U36009 ( .A(n50510), .B(n42583), .Y(n28165) );
  XNOR2XL U36010 ( .A(n50576), .B(n42582), .Y(n27383) );
  XNOR2XL U36011 ( .A(n50549), .B(n42577), .Y(n29427) );
  XNOR2XL U36012 ( .A(n50536), .B(n42576), .Y(n26901) );
  XNOR2XL U36013 ( .A(n50527), .B(n42580), .Y(n25037) );
  XNOR2XL U36014 ( .A(n50529), .B(n42581), .Y(n27051) );
  XNOR2XL U36015 ( .A(n50554), .B(n42577), .Y(n29247) );
  XNOR2XL U36016 ( .A(n50552), .B(n42577), .Y(n29397) );
  XNOR2XL U36017 ( .A(n50528), .B(n42580), .Y(n25067) );
  XNOR2XL U36018 ( .A(n50502), .B(n42583), .Y(n28315) );
  XNOR2XL U36019 ( .A(n50562), .B(n42582), .Y(n27352) );
  XNOR2XL U36020 ( .A(n50498), .B(n42583), .Y(n28405) );
  XNOR2XL U36021 ( .A(n50504), .B(n42583), .Y(n28255) );
  XNOR2XL U36022 ( .A(n50532), .B(n42581), .Y(n27081) );
  XNOR2XL U36023 ( .A(n50508), .B(n42583), .Y(n28225) );
  XNOR2XL U36024 ( .A(n50551), .B(n42577), .Y(n29367) );
  XNOR2XL U36025 ( .A(n50550), .B(n42577), .Y(n29457) );
  XNOR2XL U36026 ( .A(n51413), .B(n41303), .Y(n22451) );
  XNOR2XL U36027 ( .A(n51408), .B(n41300), .Y(n22421) );
  XNOR2XL U36028 ( .A(n51409), .B(n41302), .Y(n22431) );
  XNOR2XL U36029 ( .A(n50546), .B(n42576), .Y(n29036) );
  XNOR2XL U36030 ( .A(n50547), .B(n42576), .Y(n29096) );
  XNOR2XL U36031 ( .A(n50545), .B(n42576), .Y(n29006) );
  XOR2XL U36032 ( .A(n42494), .B(n42073), .Y(n47648) );
  XOR2XL U36033 ( .A(n42494), .B(n42095), .Y(n47504) );
  XOR2XL U36034 ( .A(n42161), .B(n41321), .Y(n25006) );
  XOR2XL U36035 ( .A(n42163), .B(n41323), .Y(n25156) );
  XOR2XL U36036 ( .A(n42113), .B(n41321), .Y(n27592) );
  XOR2XL U36037 ( .A(n42119), .B(n36877), .Y(n27171) );
  XOR2XL U36038 ( .A(n42105), .B(n36877), .Y(n28013) );
  XOR2XL U36039 ( .A(n42162), .B(n36801), .Y(n25186) );
  XOR2XL U36040 ( .A(n42164), .B(n41323), .Y(n24856) );
  XOR2XL U36041 ( .A(n42117), .B(n36873), .Y(n27231) );
  XOR2XL U36042 ( .A(n42118), .B(n41321), .Y(n27141) );
  XOR2XL U36043 ( .A(n42165), .B(n41323), .Y(n24886) );
  XOR2XL U36044 ( .A(n42120), .B(n41321), .Y(n27201) );
  XOR2XL U36045 ( .A(n42121), .B(n41323), .Y(n27291) );
  XOR2XL U36046 ( .A(n42116), .B(n36877), .Y(n27261) );
  XOR2XL U36047 ( .A(n42166), .B(n36873), .Y(n24916) );
  XOR2XL U36048 ( .A(n42167), .B(n36873), .Y(n24946) );
  XOR2XL U36049 ( .A(n42153), .B(n41323), .Y(n27110) );
  XOR2XL U36050 ( .A(n42157), .B(n41322), .Y(n25036) );
  XOR2XL U36051 ( .A(n42156), .B(n36801), .Y(n25066) );
  XOR2XL U36052 ( .A(n42155), .B(n36877), .Y(n27050) );
  XOR2XL U36053 ( .A(n42144), .B(n36877), .Y(n26839) );
  XOR2XL U36054 ( .A(n42128), .B(n36873), .Y(n29306) );
  XOR2XL U36055 ( .A(n42140), .B(n36877), .Y(n26779) );
  XOR2XL U36056 ( .A(n42142), .B(n41323), .Y(n26719) );
  XOR2XL U36057 ( .A(n42129), .B(n36801), .Y(n29336) );
  XOR2XL U36058 ( .A(n42138), .B(n36801), .Y(n29035) );
  XOR2XL U36059 ( .A(n42143), .B(n36877), .Y(n26689) );
  XOR2XL U36060 ( .A(n42150), .B(n41323), .Y(n26960) );
  XOR2XL U36061 ( .A(n42137), .B(n41321), .Y(n29095) );
  XOR2XL U36062 ( .A(n42149), .B(n36801), .Y(n26930) );
  XOR2XL U36063 ( .A(n42106), .B(n41321), .Y(n28073) );
  XOR2XL U36064 ( .A(n42175), .B(n41322), .Y(n28194) );
  XOR2XL U36065 ( .A(n42131), .B(n36801), .Y(n29276) );
  XOR2XL U36066 ( .A(n42145), .B(n36877), .Y(n26869) );
  XOR2XL U36067 ( .A(n42151), .B(n36877), .Y(n26990) );
  XOR2XL U36068 ( .A(n42135), .B(n41321), .Y(n29426) );
  XOR2XL U36069 ( .A(n42171), .B(n36877), .Y(n24796) );
  XOR2XL U36070 ( .A(n42154), .B(n41323), .Y(n27020) );
  XOR2XL U36071 ( .A(n42130), .B(n36801), .Y(n29246) );
  XOR2XL U36072 ( .A(n42183), .B(n36873), .Y(n28284) );
  XOR2XL U36073 ( .A(n42132), .B(n41321), .Y(n29396) );
  XOR2XL U36074 ( .A(n42173), .B(n36801), .Y(n28104) );
  XOR2XL U36075 ( .A(n42139), .B(n36877), .Y(n29005) );
  XOR2XL U36076 ( .A(n42174), .B(n36877), .Y(n28164) );
  XOR2XL U36077 ( .A(n42146), .B(n36801), .Y(n26809) );
  XOR2XL U36078 ( .A(n42168), .B(n41323), .Y(n24766) );
  XOR2XL U36079 ( .A(n42169), .B(n41323), .Y(n24736) );
  XOR2XL U36080 ( .A(n42148), .B(n36877), .Y(n26900) );
  XOR2XL U36081 ( .A(n42182), .B(n41322), .Y(n28314) );
  XOR2XL U36082 ( .A(n42133), .B(n36873), .Y(n29366) );
  XOR2XL U36083 ( .A(n42134), .B(n41322), .Y(n29456) );
  XOR2XL U36084 ( .A(n42170), .B(n41323), .Y(n24826) );
  XOR2XL U36085 ( .A(n42122), .B(n36877), .Y(n27351) );
  XOR2XL U36086 ( .A(n42186), .B(n36801), .Y(n28404) );
  XOR2XL U36087 ( .A(n42177), .B(n36873), .Y(n28494) );
  XOR2XL U36088 ( .A(n42180), .B(n36877), .Y(n28254) );
  XOR2XL U36089 ( .A(n42179), .B(n41322), .Y(n28524) );
  XOR2XL U36090 ( .A(n42176), .B(n41321), .Y(n28224) );
  XOR2XL U36091 ( .A(n42152), .B(n41323), .Y(n27080) );
  XOR2XL U36092 ( .A(n42187), .B(n41321), .Y(n28374) );
  XOR2XL U36093 ( .A(n42136), .B(n41321), .Y(n29065) );
  XOR2XL U36094 ( .A(n42185), .B(n36801), .Y(n28434) );
  XOR2XL U36095 ( .A(n42178), .B(n41322), .Y(n28554) );
  XOR2XL U36096 ( .A(n42184), .B(n36801), .Y(n28464) );
  XOR2XL U36097 ( .A(n42181), .B(n36877), .Y(n28344) );
  XNOR2XL U36098 ( .A(n51355), .B(n42644), .Y(n28446) );
  XNOR2XL U36099 ( .A(n51353), .B(n42644), .Y(n28386) );
  XNOR2XL U36100 ( .A(n51362), .B(n42644), .Y(n28566) );
  XNOR2XL U36101 ( .A(n51404), .B(n42644), .Y(n29077) );
  XNOR2XL U36102 ( .A(n51363), .B(n42644), .Y(n28506) );
  XNOR2XL U36103 ( .A(n51361), .B(n42644), .Y(n28536) );
  XNOR2XL U36104 ( .A(n51356), .B(n42644), .Y(n28476) );
  XNOR2XL U36105 ( .A(n50791), .B(n42508), .Y(n28041) );
  XNOR2XL U36106 ( .A(n50794), .B(n42508), .Y(n27981) );
  XNOR2XL U36107 ( .A(n50725), .B(n42508), .Y(n28102) );
  XNOR2XL U36108 ( .A(n50559), .B(n42577), .Y(n29187) );
  XNOR2XL U36109 ( .A(n51201), .B(n42554), .Y(n29183) );
  XOR2XL U36110 ( .A(n42495), .B(n42093), .Y(n47482) );
  XOR2XL U36111 ( .A(n36817), .B(n42072), .Y(n46547) );
  XOR2XL U36112 ( .A(n36808), .B(n42071), .Y(n46492) );
  XOR2XL U36113 ( .A(n36807), .B(n42073), .Y(n46536) );
  XOR2XL U36114 ( .A(n36809), .B(n42074), .Y(n46514) );
  XOR2XL U36115 ( .A(n36816), .B(n42086), .Y(n46448) );
  XOR2XL U36116 ( .A(n36811), .B(n42096), .Y(n46297) );
  XOR2XL U36117 ( .A(n36815), .B(n42087), .Y(n46437) );
  XOR2XL U36118 ( .A(n36807), .B(n42088), .Y(n46426) );
  XOR2XL U36119 ( .A(n42494), .B(n42070), .Y(n47604) );
  XOR2XL U36120 ( .A(n36808), .B(n42083), .Y(n46379) );
  XOR2XL U36121 ( .A(n36810), .B(n42080), .Y(n46357) );
  XOR2XL U36122 ( .A(n36811), .B(n42075), .Y(n46525) );
  XOR2XL U36123 ( .A(n36814), .B(n42100), .Y(n46213) );
  XOR2XL U36124 ( .A(n42494), .B(n42072), .Y(n47637) );
  XOR2XL U36125 ( .A(n36816), .B(n42095), .Y(n46263) );
  XOR2XL U36126 ( .A(n36813), .B(n42090), .Y(n46404) );
  XOR2XL U36127 ( .A(n36759), .B(n41814), .Y(n47645) );
  XOR2XL U36128 ( .A(n42494), .B(n42071), .Y(n47626) );
  XOR2XL U36129 ( .A(n36807), .B(n42081), .Y(n46368) );
  XOR2XL U36130 ( .A(n36814), .B(n42079), .Y(n46335) );
  XOR2XL U36131 ( .A(n36815), .B(n42078), .Y(n46324) );
  XOR2XL U36132 ( .A(n36815), .B(n42091), .Y(n46415) );
  XOR2XL U36133 ( .A(n36807), .B(n42082), .Y(n46386) );
  XOR2XL U36134 ( .A(n36810), .B(n42085), .Y(n46466) );
  XOR2XL U36135 ( .A(n36813), .B(n42094), .Y(n46252) );
  XOR2XL U36136 ( .A(n36807), .B(n42084), .Y(n46459) );
  XOR2XL U36137 ( .A(n36811), .B(n42097), .Y(n46224) );
  XOR2XL U36138 ( .A(n36759), .B(n41836), .Y(n47501) );
  XOR2XL U36139 ( .A(n42494), .B(n42075), .Y(n47582) );
  XOR2XL U36140 ( .A(n36817), .B(n42089), .Y(n46393) );
  XOR2XL U36141 ( .A(n42494), .B(n42094), .Y(n47493) );
  XOR2XL U36142 ( .A(n42495), .B(n42087), .Y(n47460) );
  XOR2XL U36143 ( .A(n36809), .B(n42092), .Y(n46235) );
  XOR2XL U36144 ( .A(n42494), .B(n42097), .Y(n47513) );
  XOR2XL U36145 ( .A(n42495), .B(n42086), .Y(n47449) );
  XOR2XL U36146 ( .A(n42495), .B(n42088), .Y(n47383) );
  XOR2XL U36147 ( .A(n42495), .B(n42089), .Y(n47394) );
  XOR2XL U36148 ( .A(n42495), .B(n42082), .Y(n47372) );
  XOR2XL U36149 ( .A(n36761), .B(n41818), .Y(n47304) );
  XOR2XL U36150 ( .A(n42493), .B(n42076), .Y(n47296) );
  XOR2XL U36151 ( .A(n42494), .B(n42074), .Y(n47593) );
  XOR2XL U36152 ( .A(n42494), .B(n42096), .Y(n47524) );
  XOR2XL U36153 ( .A(n42495), .B(n42091), .Y(n47416) );
  XOR2XL U36154 ( .A(n42495), .B(n42079), .Y(n47328) );
  XOR2XL U36155 ( .A(n42495), .B(n42092), .Y(n47471) );
  XOR2XL U36156 ( .A(n42495), .B(n42083), .Y(n47361) );
  XOR2XL U36157 ( .A(n42495), .B(n42085), .Y(n47438) );
  XOR2XL U36158 ( .A(n42495), .B(n42090), .Y(n47405) );
  XOR2XL U36159 ( .A(n42496), .B(n42078), .Y(n47317) );
  XOR2XL U36160 ( .A(n36816), .B(n42098), .Y(n46274) );
  XOR2XL U36161 ( .A(n36813), .B(n42099), .Y(n46285) );
  XOR2XL U36162 ( .A(n42494), .B(n42098), .Y(n47535) );
  XOR2XL U36163 ( .A(n36814), .B(n42070), .Y(n46506) );
  XOR2XL U36164 ( .A(n42494), .B(n42064), .Y(n47669) );
  XNOR2XL U36165 ( .A(n41316), .B(n41810), .Y(n46481) );
  XNOR2XL U36166 ( .A(n41309), .B(n41811), .Y(n46472) );
  XNOR2XL U36167 ( .A(n42496), .B(n42068), .Y(n47655) );
  XNOR2XL U36168 ( .A(n36816), .B(n42093), .Y(n46244) );
  XNOR2XL U36169 ( .A(n41316), .B(n41834), .Y(n46245) );
  XNOR2XL U36170 ( .A(n41317), .B(n41812), .Y(n46504) );
  XOR2XL U36171 ( .A(n36791), .B(n41803), .Y(n47667) );
  NOR3X2 U36172 ( .A(n29137), .B(n29141), .C(n29127), .Y(n43611) );
  XOR2XL U36173 ( .A(n41305), .B(n41799), .Y(n46286) );
  XOR2XL U36174 ( .A(n36779), .B(n42061), .Y(n46287) );
  XOR2XL U36175 ( .A(n41328), .B(n41801), .Y(n46273) );
  XOR2XL U36176 ( .A(n41333), .B(n41802), .Y(n46284) );
  XOR2XL U36177 ( .A(n36793), .B(n41805), .Y(n47545) );
  XOR2XL U36178 ( .A(n36746), .B(n41799), .Y(n47544) );
  XOR2XL U36179 ( .A(n41296), .B(n41805), .Y(n46283) );
  NAND3XL U36180 ( .A(n12387), .B(n11085), .C(n11208), .Y(n48504) );
  NAND2XL U36181 ( .A(n11094), .B(n11092), .Y(n48505) );
  NAND4XL U36182 ( .A(net209225), .B(n12303), .C(n10846), .D(n10847), .Y(
        n48506) );
  NAND4XL U36183 ( .A(n12144), .B(n12794), .C(n10566), .D(n12079), .Y(n48208)
         );
  NAND2XL U36184 ( .A(n12795), .B(n12146), .Y(n48206) );
  NAND2XL U36185 ( .A(net209249), .B(n12324), .Y(n48486) );
  NAND3XL U36186 ( .A(n11200), .B(n12384), .C(n11131), .Y(n48487) );
  XOR2XL U36187 ( .A(n36753), .B(n41841), .Y(n47567) );
  XOR2XL U36188 ( .A(n41309), .B(n41840), .Y(n46282) );
  NAND4XL U36189 ( .A(n11379), .B(n12929), .C(net210099), .D(n11386), .Y(
        n48080) );
  NAND4XL U36190 ( .A(n12723), .B(n10554), .C(n12065), .D(n12063), .Y(n48215)
         );
  XOR2XL U36191 ( .A(n36755), .B(n41826), .Y(n47435) );
  NAND3XL U36192 ( .A(n12954), .B(n13015), .C(n12959), .Y(n48060) );
  NAND2XL U36193 ( .A(n10553), .B(n10606), .Y(n48213) );
  NAND2XL U36194 ( .A(n12741), .B(n12793), .Y(n48194) );
  NAND4BXL U36195 ( .AN(n48226), .B(n48225), .C(n10543), .D(n12708), .Y(n48230) );
  NAND4XL U36196 ( .A(n41776), .B(n12033), .C(n12035), .D(n48228), .Y(n48229)
         );
  NAND2XL U36197 ( .A(n12049), .B(n12151), .Y(n48226) );
  NAND3XL U36198 ( .A(n11075), .B(n11073), .C(n12388), .Y(n48512) );
  NAND2XL U36199 ( .A(n11117), .B(n11115), .Y(n48493) );
  NAND2XL U36200 ( .A(n10852), .B(n10853), .Y(n48494) );
  NAND2XL U36201 ( .A(n11138), .B(n10870), .Y(n48477) );
  NAND2XL U36202 ( .A(n48057), .B(n11423), .Y(n48059) );
  NAND2XL U36203 ( .A(net209268), .B(n11140), .Y(n48476) );
  OR2X4 U36204 ( .A(n29132), .B(n29123), .Y(n43620) );
  INVXL U36205 ( .A(n12035), .Y(net209964) );
  INVXL U36206 ( .A(net209927), .Y(net209926) );
  INVXL U36207 ( .A(n11389), .Y(net210100) );
  AND3XL U36208 ( .A(n12087), .B(n12747), .C(n12089), .Y(n48196) );
  AND2XL U36209 ( .A(net209202), .B(n12287), .Y(n48511) );
  XOR2XL U36210 ( .A(n41927), .B(n41314), .Y(n23166) );
  XOR2XL U36211 ( .A(n41844), .B(n36759), .Y(n20391) );
  XOR2XL U36212 ( .A(n41843), .B(n36760), .Y(n20401) );
  XOR2XL U36213 ( .A(n41922), .B(n41312), .Y(n23136) );
  XOR2XL U36214 ( .A(n41923), .B(n41311), .Y(n23156) );
  XOR2XL U36215 ( .A(n41886), .B(n41311), .Y(n24088) );
  XOR2XL U36216 ( .A(n41900), .B(n41316), .Y(n235610) );
  XOR2XL U36217 ( .A(n41849), .B(n36759), .Y(n20217) );
  XOR2XL U36218 ( .A(n41862), .B(n36755), .Y(n20125) );
  XOR2XL U36219 ( .A(n41859), .B(n36761), .Y(n20165) );
  XOR2XL U36220 ( .A(n41857), .B(n36756), .Y(n20145) );
  XOR2XL U36221 ( .A(n41912), .B(n41311), .Y(n23481) );
  XOR2XL U36222 ( .A(n41848), .B(n36761), .Y(n20279) );
  XOR2XL U36223 ( .A(n41847), .B(n36755), .Y(n20269) );
  XOR2XL U36224 ( .A(n41860), .B(n36755), .Y(n20175) );
  XOR2XL U36225 ( .A(n41910), .B(n41309), .Y(n23461) );
  XOR2XL U36226 ( .A(n41903), .B(n41309), .Y(n23521) );
  XOR2XL U36227 ( .A(n41901), .B(n41309), .Y(n23501) );
  XOR2XL U36228 ( .A(n41872), .B(n36760), .Y(n19556) );
  XOR2XL U36229 ( .A(n41850), .B(n36755), .Y(n20207) );
  XOR2XL U36230 ( .A(n41854), .B(n36757), .Y(n20247) );
  XOR2XL U36231 ( .A(n41878), .B(n41318), .Y(n22329) );
  XOR2XL U36232 ( .A(n41871), .B(n36756), .Y(n19566) );
  XOR2XL U36233 ( .A(n41892), .B(n36753), .Y(n19779) );
  XOR2XL U36234 ( .A(n41894), .B(n36754), .Y(n19759) );
  XOR2XL U36235 ( .A(n41863), .B(n36760), .Y(n20135) );
  XOR2XL U36236 ( .A(n41856), .B(n36759), .Y(n20227) );
  XOR2XL U36237 ( .A(n41887), .B(n41318), .Y(n24068) );
  XOR2XL U36238 ( .A(n41852), .B(n36760), .Y(n20186) );
  XOR2XL U36239 ( .A(n41885), .B(n36759), .Y(n19728) );
  XOR2XL U36240 ( .A(n41864), .B(n36753), .Y(n20104) );
  XOR2XL U36241 ( .A(n41874), .B(n36761), .Y(n19626) );
  XOR2XL U36242 ( .A(n41926), .B(n41312), .Y(n23196) );
  XOR2XL U36243 ( .A(n41853), .B(n36754), .Y(n20257) );
  XOR2XL U36244 ( .A(n41851), .B(n36753), .Y(n20197) );
  XOR2XL U36245 ( .A(n41875), .B(n36759), .Y(n19646) );
  XOR2XL U36246 ( .A(n41910), .B(n36760), .Y(n21090) );
  XOR2XL U36247 ( .A(n41895), .B(n36754), .Y(n19769) );
  XOR2XL U36248 ( .A(n41855), .B(n36756), .Y(n20237) );
  XOR2XL U36249 ( .A(n41902), .B(n41310), .Y(n23511) );
  XOR2XL U36250 ( .A(n41886), .B(n36757), .Y(n19718) );
  XOR2XL U36251 ( .A(n41932), .B(n41318), .Y(n22976) );
  XOR2XL U36252 ( .A(n41877), .B(n36757), .Y(n19849) );
  XOR2XL U36253 ( .A(n41896), .B(n36756), .Y(n19749) );
  XOR2XL U36254 ( .A(n41887), .B(n36760), .Y(n19708) );
  XOR2XL U36255 ( .A(n41898), .B(n36757), .Y(n21019) );
  XOR2XL U36256 ( .A(n41930), .B(n41316), .Y(n22956) );
  XOR2XL U36257 ( .A(n41876), .B(n36755), .Y(n19636) );
  XOR2XL U36258 ( .A(n41911), .B(n36759), .Y(n21120) );
  XOR2XL U36259 ( .A(n41878), .B(n36755), .Y(n19819) );
  XOR2XL U36260 ( .A(n41880), .B(n36757), .Y(n19839) );
  XOR2XL U36261 ( .A(n41933), .B(n41317), .Y(n22996) );
  XOR2XL U36262 ( .A(n41883), .B(n36755), .Y(n19668) );
  XOR2XL U36263 ( .A(n41912), .B(n36753), .Y(n21110) );
  XOR2XL U36264 ( .A(n41913), .B(n36759), .Y(n19960) );
  XOR2XL U36265 ( .A(n41935), .B(n41314), .Y(n23016) );
  XOR2XL U36266 ( .A(n41899), .B(n36754), .Y(n21040) );
  XOR2XL U36267 ( .A(n41900), .B(n36759), .Y(n21029) );
  XOR2XL U36268 ( .A(n41882), .B(n36756), .Y(n19678) );
  XOR2XL U36269 ( .A(n41884), .B(n36759), .Y(n19657) );
  XOR2XL U36270 ( .A(n41868), .B(n36755), .Y(n19576) );
  XOR2XL U36271 ( .A(n41928), .B(n36754), .Y(n19990) );
  XOR2XL U36272 ( .A(n41930), .B(n36755), .Y(n21594) );
  XOR2XL U36273 ( .A(n41867), .B(n36753), .Y(n19586) );
  XOR2XL U36274 ( .A(n41927), .B(n36753), .Y(n19980) );
  XOR2XL U36275 ( .A(n41937), .B(n41311), .Y(n22926) );
  XOR2XL U36276 ( .A(n41879), .B(n36761), .Y(n19829) );
  XOR2XL U36277 ( .A(n41902), .B(n36760), .Y(n20968) );
  XOR2XL U36278 ( .A(n41934), .B(n41318), .Y(n23006) );
  XOR2XL U36279 ( .A(n41914), .B(n36753), .Y(n19950) );
  XOR2XL U36280 ( .A(n41881), .B(n36760), .Y(n19688) );
  XOR2XL U36281 ( .A(n41901), .B(n36754), .Y(n20978) );
  XOR2XL U36282 ( .A(n41931), .B(n36761), .Y(n21584) );
  XOR2XL U36283 ( .A(n41888), .B(n36760), .Y(n19698) );
  XOR2XL U36284 ( .A(n41936), .B(n41310), .Y(n22986) );
  XOR2XL U36285 ( .A(n41915), .B(n36755), .Y(n19940) );
  XOR2XL U36286 ( .A(n41932), .B(n36761), .Y(n21574) );
  XOR2XL U36287 ( .A(n41917), .B(n36759), .Y(n19910) );
  XOR2XL U36288 ( .A(n41934), .B(n36759), .Y(n21494) );
  XOR2XL U36289 ( .A(n41904), .B(n36753), .Y(n20999) );
  XOR2XL U36290 ( .A(n41903), .B(n36757), .Y(n20989) );
  XOR2XL U36291 ( .A(n41936), .B(n36757), .Y(n21524) );
  XOR2XL U36292 ( .A(n41916), .B(n36759), .Y(n19930) );
  XNOR2XL U36293 ( .A(n51224), .B(n36716), .Y(n20399) );
  XNOR2XL U36294 ( .A(n51140), .B(n41331), .Y(n23164) );
  XNOR2XL U36295 ( .A(n51145), .B(n41329), .Y(n23134) );
  XNOR2XL U36296 ( .A(n51144), .B(n41327), .Y(n23154) );
  XNOR2XL U36297 ( .A(n50796), .B(n42470), .Y(n20400) );
  XNOR2XL U36298 ( .A(n51347), .B(n42694), .Y(n31343) );
  XNOR2XL U36299 ( .A(n51344), .B(n42694), .Y(n31433) );
  XNOR2XL U36300 ( .A(n51345), .B(n42691), .Y(n31463) );
  XNOR2XL U36301 ( .A(n51339), .B(n42702), .Y(n31193) );
  XNOR2XL U36302 ( .A(n51341), .B(n42691), .Y(n31283) );
  XNOR2XL U36303 ( .A(n51342), .B(n42701), .Y(n31493) );
  XNOR2XL U36304 ( .A(n51343), .B(n42701), .Y(n31523) );
  XNOR2XL U36305 ( .A(n51340), .B(n42702), .Y(n31253) );
  XNOR2XL U36306 ( .A(n51338), .B(n42697), .Y(n31223) );
  XNOR2XL U36307 ( .A(n50712), .B(n36859), .Y(n23165) );
  XNOR2XL U36308 ( .A(n50716), .B(n36856), .Y(n23155) );
  XOR2XL U36309 ( .A(n41918), .B(n41312), .Y(n23266) );
  XOR2XL U36310 ( .A(n41919), .B(n41318), .Y(n23256) );
  XOR2XL U36311 ( .A(n41920), .B(n41311), .Y(n23246) );
  XNOR2XL U36312 ( .A(n51010), .B(n36791), .Y(n20398) );
  XNOR2XL U36313 ( .A(n50926), .B(n41293), .Y(n23163) );
  XNOR2XL U36314 ( .A(n50931), .B(n41294), .Y(n23133) );
  XNOR2XL U36315 ( .A(n50930), .B(n41294), .Y(n23153) );
  XOR2XL U36316 ( .A(n42191), .B(n42656), .Y(n31366) );
  XOR2XL U36317 ( .A(n41933), .B(n36898), .Y(n31340) );
  XOR2XL U36318 ( .A(n42192), .B(n36886), .Y(n31344) );
  XOR2XL U36319 ( .A(n42193), .B(n42656), .Y(n31336) );
  XOR2XL U36320 ( .A(n41934), .B(n42608), .Y(n31332) );
  XOR2XL U36321 ( .A(n41936), .B(n36901), .Y(n31430) );
  XOR2XL U36322 ( .A(n42195), .B(n36880), .Y(n31434) );
  XOR2XL U36323 ( .A(n41937), .B(n42605), .Y(n31422) );
  XOR2XL U36324 ( .A(n42196), .B(n42656), .Y(n31426) );
  XOR2XL U36325 ( .A(n41935), .B(n36895), .Y(n31460) );
  XOR2XL U36326 ( .A(n41941), .B(n36900), .Y(n31190) );
  XOR2XL U36327 ( .A(n42194), .B(n36882), .Y(n31464) );
  XOR2XL U36328 ( .A(n42200), .B(n36881), .Y(n31194) );
  XOR2XL U36329 ( .A(n42201), .B(n42656), .Y(n31186) );
  XOR2XL U36330 ( .A(n41942), .B(n42608), .Y(n31182) );
  XOR2XL U36331 ( .A(n42195), .B(n42656), .Y(n31456) );
  XOR2XL U36332 ( .A(n41936), .B(n42607), .Y(n31452) );
  XOR2XL U36333 ( .A(n41939), .B(n36892), .Y(n31280) );
  XOR2XL U36334 ( .A(n42198), .B(n36879), .Y(n31284) );
  XOR2XL U36335 ( .A(n41940), .B(n42607), .Y(n31272) );
  XOR2XL U36336 ( .A(n42199), .B(n42656), .Y(n31276) );
  XOR2XL U36337 ( .A(n41938), .B(n36894), .Y(n31490) );
  XOR2XL U36338 ( .A(n42197), .B(n36883), .Y(n31494) );
  XOR2XL U36339 ( .A(n41939), .B(n42607), .Y(n31482) );
  XOR2XL U36340 ( .A(n42198), .B(n42656), .Y(n31486) );
  XOR2XL U36341 ( .A(n41937), .B(n36891), .Y(n31520) );
  XOR2XL U36342 ( .A(n41940), .B(n36893), .Y(n31250) );
  XOR2XL U36343 ( .A(n42196), .B(n36889), .Y(n31524) );
  XOR2XL U36344 ( .A(n42199), .B(n36881), .Y(n31254) );
  XOR2XL U36345 ( .A(n42200), .B(n42656), .Y(n31246) );
  XOR2XL U36346 ( .A(n41941), .B(n42607), .Y(n31242) );
  XOR2XL U36347 ( .A(n42197), .B(n42656), .Y(n31516) );
  XOR2XL U36348 ( .A(n41942), .B(n36898), .Y(n31220) );
  XOR2XL U36349 ( .A(n41938), .B(n42607), .Y(n31512) );
  XOR2XL U36350 ( .A(n42201), .B(n36887), .Y(n31224) );
  XOR2XL U36351 ( .A(n41943), .B(n42607), .Y(n31212) );
  XOR2XL U36352 ( .A(n42202), .B(n42656), .Y(n31216) );
  XNOR2XL U36353 ( .A(n51142), .B(n42554), .Y(n28461) );
  XNOR2XL U36354 ( .A(n51145), .B(n42554), .Y(n28341) );
  XNOR2XL U36355 ( .A(n50534), .B(n36765), .Y(n19791) );
  XNOR2XL U36356 ( .A(n50533), .B(n36770), .Y(n19781) );
  XNOR2XL U36357 ( .A(n50560), .B(n36773), .Y(n19608) );
  XNOR2XL U36358 ( .A(n50529), .B(n36765), .Y(n19751) );
  XNOR2XL U36359 ( .A(n51402), .B(n36918), .Y(n22331) );
  XNOR2XL U36360 ( .A(n51409), .B(n36742), .Y(n19568) );
  XNOR2XL U36361 ( .A(n51408), .B(n36750), .Y(n19558) );
  XNOR2XL U36362 ( .A(n51407), .B(n36743), .Y(n19618) );
  XNOR2XL U36363 ( .A(n51406), .B(n36748), .Y(n19628) );
  XNOR2XL U36364 ( .A(n51414), .B(n36747), .Y(n19598) );
  XNOR2XL U36365 ( .A(n51413), .B(n36748), .Y(n19588) );
  XNOR2XL U36366 ( .A(n51412), .B(n36743), .Y(n19578) );
  XOR2XL U36367 ( .A(n41929), .B(n42519), .Y(n31562) );
  XOR2XL U36368 ( .A(n41934), .B(n42519), .Y(n31382) );
  XOR2XL U36369 ( .A(n41933), .B(n42519), .Y(n31352) );
  XOR2XL U36370 ( .A(n41935), .B(n42519), .Y(n31322) );
  XOR2XL U36371 ( .A(n41937), .B(n42519), .Y(n31442) );
  XOR2XL U36372 ( .A(n41938), .B(n42519), .Y(n31412) );
  XOR2XL U36373 ( .A(n41943), .B(n42518), .Y(n31172) );
  XNOR2XL U36374 ( .A(n50928), .B(n42544), .Y(n28460) );
  XNOR2XL U36375 ( .A(n51219), .B(n36716), .Y(n20277) );
  XNOR2XL U36376 ( .A(n51208), .B(n36722), .Y(n20163) );
  XNOR2XL U36377 ( .A(n51210), .B(n36714), .Y(n20143) );
  XNOR2XL U36378 ( .A(n51155), .B(n41327), .Y(n23479) );
  XNOR2XL U36379 ( .A(n51207), .B(n36714), .Y(n20173) );
  XNOR2XL U36380 ( .A(n51220), .B(n36714), .Y(n20267) );
  XNOR2XL U36381 ( .A(n51166), .B(n41330), .Y(n23499) );
  XNOR2XL U36382 ( .A(n51195), .B(n36717), .Y(n19554) );
  XNOR2XL U36383 ( .A(n51217), .B(n36716), .Y(n20205) );
  XNOR2XL U36384 ( .A(n51164), .B(n41331), .Y(n23519) );
  XNOR2XL U36385 ( .A(n51157), .B(n41333), .Y(n23459) );
  XNOR2XL U36386 ( .A(n51213), .B(n36715), .Y(n20245) );
  XNOR2XL U36387 ( .A(n51189), .B(n41327), .Y(n22327) );
  XNOR2XL U36388 ( .A(n51196), .B(n36717), .Y(n19564) );
  XNOR2XL U36389 ( .A(n51175), .B(n36720), .Y(n19777) );
  XNOR2XL U36390 ( .A(n51173), .B(n36721), .Y(n19757) );
  XNOR2XL U36391 ( .A(n51211), .B(n36716), .Y(n20225) );
  XNOR2XL U36392 ( .A(n51215), .B(n36722), .Y(n20184) );
  XNOR2XL U36393 ( .A(n51204), .B(n36718), .Y(n20133) );
  XNOR2XL U36394 ( .A(n51180), .B(n41331), .Y(n24066) );
  XNOR2XL U36395 ( .A(n51203), .B(n36715), .Y(n20102) );
  XNOR2XL U36396 ( .A(n51182), .B(n36718), .Y(n19726) );
  XNOR2XL U36397 ( .A(n51193), .B(n36722), .Y(n19624) );
  XNOR2XL U36398 ( .A(n51223), .B(n36716), .Y(n20389) );
  XNOR2XL U36399 ( .A(n51141), .B(n41332), .Y(n23194) );
  XNOR2XL U36400 ( .A(n51214), .B(n36721), .Y(n20255) );
  XNOR2XL U36401 ( .A(n51216), .B(n36716), .Y(n20195) );
  XNOR2XL U36402 ( .A(n51192), .B(n36721), .Y(n19644) );
  XNOR2XL U36403 ( .A(n51157), .B(n36715), .Y(n21088) );
  XNOR2XL U36404 ( .A(n51165), .B(n41332), .Y(n23509) );
  XNOR2XL U36405 ( .A(n51172), .B(n36716), .Y(n19767) );
  XNOR2XL U36406 ( .A(n51181), .B(n36718), .Y(n19716) );
  XNOR2XL U36407 ( .A(n51212), .B(n36717), .Y(n20235) );
  XNOR2XL U36408 ( .A(n51135), .B(n41332), .Y(n22974) );
  XNOR2XL U36409 ( .A(n51171), .B(n36714), .Y(n19747) );
  XNOR2XL U36410 ( .A(n51190), .B(n36722), .Y(n19847) );
  XNOR2XL U36411 ( .A(n51180), .B(n36720), .Y(n19706) );
  XNOR2XL U36412 ( .A(n51169), .B(n36715), .Y(n21017) );
  XNOR2XL U36413 ( .A(n51191), .B(n36722), .Y(n19634) );
  XNOR2XL U36414 ( .A(n51137), .B(n41330), .Y(n22954) );
  XNOR2XL U36415 ( .A(n51156), .B(n36720), .Y(n21118) );
  XNOR2XL U36416 ( .A(n51189), .B(n36716), .Y(n19817) );
  XNOR2XL U36417 ( .A(n51187), .B(n36721), .Y(n19837) );
  XNOR2XL U36418 ( .A(n51134), .B(n41329), .Y(n22994) );
  XNOR2XL U36419 ( .A(n51155), .B(n36720), .Y(n21108) );
  XNOR2XL U36420 ( .A(n51184), .B(n36717), .Y(n19666) );
  XNOR2XL U36421 ( .A(n51132), .B(n41331), .Y(n23014) );
  XNOR2XL U36422 ( .A(n51154), .B(n36715), .Y(n19958) );
  XNOR2XL U36423 ( .A(n51167), .B(n36715), .Y(n21027) );
  XNOR2XL U36424 ( .A(n51168), .B(n36720), .Y(n21038) );
  XNOR2XL U36425 ( .A(n51185), .B(n36718), .Y(n19676) );
  XNOR2XL U36426 ( .A(n51183), .B(n36718), .Y(n19655) );
  XNOR2XL U36427 ( .A(n51199), .B(n36720), .Y(n19574) );
  XNOR2XL U36428 ( .A(n51139), .B(n36720), .Y(n19988) );
  XNOR2XL U36429 ( .A(n51137), .B(n36721), .Y(n21592) );
  XNOR2XL U36430 ( .A(n51130), .B(n41327), .Y(n22924) );
  XNOR2XL U36431 ( .A(n51165), .B(n36714), .Y(n20966) );
  XNOR2XL U36432 ( .A(n51200), .B(n36720), .Y(n19584) );
  XNOR2XL U36433 ( .A(n51140), .B(n36717), .Y(n19978) );
  XNOR2XL U36434 ( .A(n51153), .B(n36717), .Y(n19948) );
  XNOR2XL U36435 ( .A(n51188), .B(n36714), .Y(n19827) );
  XNOR2XL U36436 ( .A(n51133), .B(n41327), .Y(n23004) );
  XNOR2XL U36437 ( .A(n51186), .B(n36722), .Y(n19686) );
  XNOR2XL U36438 ( .A(n51166), .B(n36717), .Y(n20976) );
  XNOR2XL U36439 ( .A(n51179), .B(n36720), .Y(n19696) );
  XNOR2XL U36440 ( .A(n51136), .B(n36718), .Y(n21582) );
  XNOR2XL U36441 ( .A(n51135), .B(n36722), .Y(n21572) );
  XNOR2XL U36442 ( .A(n51131), .B(n41330), .Y(n22984) );
  XNOR2XL U36443 ( .A(n51152), .B(n36718), .Y(n19938) );
  XNOR2XL U36444 ( .A(n51150), .B(n36718), .Y(n19908) );
  XNOR2XL U36445 ( .A(n51133), .B(n36716), .Y(n21492) );
  XNOR2XL U36446 ( .A(n51163), .B(n36721), .Y(n20997) );
  XNOR2XL U36447 ( .A(n51131), .B(n36715), .Y(n21522) );
  XNOR2XL U36448 ( .A(n51151), .B(n36721), .Y(n19928) );
  XNOR2XL U36449 ( .A(n51164), .B(n36714), .Y(n20987) );
  XNOR2XL U36450 ( .A(n51147), .B(n36717), .Y(n19888) );
  XNOR2XL U36451 ( .A(n51149), .B(n36721), .Y(n19918) );
  XNOR2XL U36452 ( .A(n50739), .B(n36858), .Y(n235600) );
  XNOR2XL U36453 ( .A(n50777), .B(n42468), .Y(n20124) );
  XNOR2XL U36454 ( .A(n50791), .B(n42469), .Y(n20278) );
  XNOR2XL U36455 ( .A(n50780), .B(n42468), .Y(n20164) );
  XNOR2XL U36456 ( .A(n50782), .B(n42468), .Y(n20144) );
  XNOR2XL U36457 ( .A(n50727), .B(n36858), .Y(n23480) );
  XNOR2XL U36458 ( .A(n50792), .B(n42469), .Y(n20268) );
  XNOR2XL U36459 ( .A(n50779), .B(n42468), .Y(n20174) );
  XNOR2XL U36460 ( .A(n50738), .B(n36858), .Y(n23500) );
  XNOR2XL U36461 ( .A(n50729), .B(n36853), .Y(n23460) );
  XNOR2XL U36462 ( .A(n50736), .B(n36857), .Y(n23520) );
  XNOR2XL U36463 ( .A(n50767), .B(n42465), .Y(n19555) );
  XNOR2XL U36464 ( .A(n50789), .B(n42469), .Y(n20206) );
  XNOR2XL U36465 ( .A(n50785), .B(n42469), .Y(n20246) );
  XNOR2XL U36466 ( .A(n50761), .B(n36860), .Y(n22328) );
  XNOR2XL U36467 ( .A(n50768), .B(n42465), .Y(n19565) );
  XNOR2XL U36468 ( .A(n50747), .B(n42468), .Y(n19778) );
  XNOR2XL U36469 ( .A(n50745), .B(n42468), .Y(n19758) );
  XNOR2XL U36470 ( .A(n50783), .B(n42469), .Y(n20226) );
  XNOR2XL U36471 ( .A(n50776), .B(n42468), .Y(n20134) );
  XNOR2XL U36472 ( .A(n50752), .B(n36857), .Y(n24067) );
  XNOR2XL U36473 ( .A(n50787), .B(n42469), .Y(n20185) );
  XNOR2XL U36474 ( .A(n50754), .B(n42468), .Y(n19727) );
  XNOR2XL U36475 ( .A(n50775), .B(n42468), .Y(n20103) );
  XNOR2XL U36476 ( .A(n50765), .B(n42465), .Y(n19625) );
  XNOR2XL U36477 ( .A(n50713), .B(n36860), .Y(n23195) );
  XNOR2XL U36478 ( .A(n50786), .B(n42469), .Y(n20256) );
  XNOR2XL U36479 ( .A(n50795), .B(n42469), .Y(n20390) );
  XNOR2XL U36480 ( .A(n50788), .B(n42469), .Y(n20196) );
  XNOR2XL U36481 ( .A(n50764), .B(n42465), .Y(n19645) );
  XNOR2XL U36482 ( .A(n50729), .B(n42460), .Y(n21089) );
  XNOR2XL U36483 ( .A(n50744), .B(n42456), .Y(n19768) );
  XNOR2XL U36484 ( .A(n50737), .B(n36854), .Y(n23510) );
  XNOR2XL U36485 ( .A(n50784), .B(n42469), .Y(n20236) );
  XNOR2XL U36486 ( .A(n50753), .B(n42468), .Y(n19717) );
  XNOR2XL U36487 ( .A(n50707), .B(n36851), .Y(n22975) );
  XNOR2XL U36488 ( .A(n50762), .B(n42466), .Y(n19848) );
  XNOR2XL U36489 ( .A(n50743), .B(n42468), .Y(n19748) );
  XNOR2XL U36490 ( .A(n50752), .B(n42466), .Y(n19707) );
  XNOR2XL U36491 ( .A(n50741), .B(n42459), .Y(n21018) );
  XNOR2XL U36492 ( .A(n50709), .B(n36850), .Y(n22955) );
  XNOR2XL U36493 ( .A(n50763), .B(n42465), .Y(n19635) );
  XNOR2XL U36494 ( .A(n50728), .B(n42460), .Y(n21119) );
  XNOR2XL U36495 ( .A(n50761), .B(n42466), .Y(n19818) );
  XNOR2XL U36496 ( .A(n50759), .B(n42466), .Y(n19838) );
  XNOR2XL U36497 ( .A(n50706), .B(n36859), .Y(n22995) );
  XNOR2XL U36498 ( .A(n50727), .B(n42460), .Y(n21109) );
  XNOR2XL U36499 ( .A(n50756), .B(n42465), .Y(n19667) );
  XNOR2XL U36500 ( .A(n50704), .B(n36850), .Y(n23015) );
  XNOR2XL U36501 ( .A(n50726), .B(n42467), .Y(n19959) );
  XNOR2XL U36502 ( .A(n50740), .B(n42459), .Y(n21039) );
  XNOR2XL U36503 ( .A(n50739), .B(n42459), .Y(n21028) );
  XNOR2XL U36504 ( .A(n50757), .B(n42465), .Y(n19677) );
  XNOR2XL U36505 ( .A(n50755), .B(n42465), .Y(n19656) );
  XNOR2XL U36506 ( .A(n50771), .B(n42465), .Y(n19575) );
  XNOR2XL U36507 ( .A(n50711), .B(n42467), .Y(n19989) );
  XNOR2XL U36508 ( .A(n50709), .B(n42466), .Y(n21593) );
  XNOR2XL U36509 ( .A(n50702), .B(n36851), .Y(n22925) );
  XNOR2XL U36510 ( .A(n50772), .B(n42465), .Y(n19585) );
  XNOR2XL U36511 ( .A(n50712), .B(n42467), .Y(n19979) );
  XNOR2XL U36512 ( .A(n50737), .B(n42459), .Y(n20967) );
  XNOR2XL U36513 ( .A(n50760), .B(n42466), .Y(n19828) );
  XNOR2XL U36514 ( .A(n50705), .B(n36854), .Y(n23005) );
  XNOR2XL U36515 ( .A(n50725), .B(n42467), .Y(n19949) );
  XNOR2XL U36516 ( .A(n50758), .B(n42465), .Y(n19687) );
  XNOR2XL U36517 ( .A(n50738), .B(n42459), .Y(n20977) );
  XNOR2XL U36518 ( .A(n50708), .B(n42466), .Y(n21583) );
  XNOR2XL U36519 ( .A(n50751), .B(n42456), .Y(n19697) );
  XNOR2XL U36520 ( .A(n50703), .B(n36853), .Y(n22985) );
  XNOR2XL U36521 ( .A(n50724), .B(n42467), .Y(n19939) );
  XNOR2XL U36522 ( .A(n50707), .B(n42466), .Y(n21573) );
  XNOR2XL U36523 ( .A(n50722), .B(n42466), .Y(n19909) );
  XNOR2XL U36524 ( .A(n50705), .B(n42459), .Y(n21493) );
  XNOR2XL U36525 ( .A(n50735), .B(n42459), .Y(n20998) );
  XNOR2XL U36526 ( .A(n50736), .B(n42459), .Y(n20988) );
  XNOR2XL U36527 ( .A(n50703), .B(n42459), .Y(n21523) );
  XNOR2XL U36528 ( .A(n50723), .B(n42467), .Y(n19929) );
  XNOR2XL U36529 ( .A(n50719), .B(n42466), .Y(n19889) );
  XNOR2XL U36530 ( .A(n50721), .B(n42466), .Y(n19919) );
  XNOR2XL U36531 ( .A(n50288), .B(n42670), .Y(n31393) );
  XNOR2XL U36532 ( .A(n50289), .B(n42711), .Y(n31401) );
  XNOR2XL U36533 ( .A(n50919), .B(n42616), .Y(n31329) );
  XNOR2XL U36534 ( .A(n50290), .B(n42711), .Y(n31371) );
  XNOR2XL U36535 ( .A(n50288), .B(n42704), .Y(n31341) );
  XNOR2XL U36536 ( .A(n50287), .B(n42676), .Y(n31333) );
  XNOR2XL U36537 ( .A(n50916), .B(n42617), .Y(n31419) );
  XNOR2XL U36538 ( .A(n50284), .B(n42670), .Y(n31423) );
  XNOR2XL U36539 ( .A(n50285), .B(n42711), .Y(n31431) );
  XNOR2XL U36540 ( .A(n50917), .B(n42617), .Y(n31449) );
  XNOR2XL U36541 ( .A(n50911), .B(n42616), .Y(n31179) );
  XNOR2XL U36542 ( .A(n50286), .B(n42711), .Y(n31461) );
  XNOR2XL U36543 ( .A(n50285), .B(n42670), .Y(n31453) );
  XNOR2XL U36544 ( .A(n50279), .B(n42670), .Y(n31183) );
  XNOR2XL U36545 ( .A(n50280), .B(n42704), .Y(n31191) );
  XNOR2XL U36546 ( .A(n50913), .B(n42616), .Y(n31269) );
  XNOR2XL U36547 ( .A(n50914), .B(n42617), .Y(n31479) );
  XNOR2XL U36548 ( .A(n50281), .B(n42671), .Y(n31273) );
  XNOR2XL U36549 ( .A(n50282), .B(n42704), .Y(n31281) );
  XNOR2XL U36550 ( .A(n50282), .B(n42670), .Y(n31483) );
  XNOR2XL U36551 ( .A(n50283), .B(n42711), .Y(n31491) );
  XNOR2XL U36552 ( .A(n50915), .B(n42617), .Y(n31509) );
  XNOR2XL U36553 ( .A(n51005), .B(n36799), .Y(n20276) );
  XNOR2XL U36554 ( .A(n50994), .B(n36793), .Y(n20162) );
  XNOR2XL U36555 ( .A(n50996), .B(n36789), .Y(n20142) );
  XNOR2XL U36556 ( .A(n50941), .B(n41296), .Y(n23478) );
  XNOR2XL U36557 ( .A(n50963), .B(n36792), .Y(n19806) );
  XNOR2XL U36558 ( .A(n50993), .B(n36796), .Y(n20172) );
  XNOR2XL U36559 ( .A(n51006), .B(n36790), .Y(n20266) );
  XNOR2XL U36560 ( .A(n50952), .B(n41295), .Y(n23498) );
  XNOR2XL U36561 ( .A(n50981), .B(n36790), .Y(n19553) );
  XNOR2XL U36562 ( .A(n51003), .B(n36798), .Y(n20204) );
  XNOR2XL U36563 ( .A(n50999), .B(n36790), .Y(n20244) );
  XNOR2XL U36564 ( .A(n50950), .B(n41296), .Y(n23518) );
  XNOR2XL U36565 ( .A(n50943), .B(n41297), .Y(n23458) );
  XNOR2XL U36566 ( .A(n50961), .B(n36795), .Y(n19776) );
  XNOR2XL U36567 ( .A(n50975), .B(n41295), .Y(n22326) );
  XNOR2XL U36568 ( .A(n50982), .B(n36793), .Y(n19563) );
  XNOR2XL U36569 ( .A(n50980), .B(n36797), .Y(n19613) );
  XNOR2XL U36570 ( .A(n50959), .B(n36792), .Y(n19756) );
  XNOR2XL U36571 ( .A(n50997), .B(n36797), .Y(n20224) );
  XNOR2XL U36572 ( .A(n51001), .B(n36793), .Y(n20183) );
  XNOR2XL U36573 ( .A(n50990), .B(n36797), .Y(n20132) );
  XNOR2XL U36574 ( .A(n50966), .B(n41295), .Y(n24065) );
  XNOR2XL U36575 ( .A(n50989), .B(n36789), .Y(n20101) );
  XNOR2XL U36576 ( .A(n50968), .B(n36792), .Y(n19725) );
  XNOR2XL U36577 ( .A(n50979), .B(n36796), .Y(n19623) );
  XNOR2XL U36578 ( .A(n51009), .B(n36795), .Y(n20388) );
  XNOR2XL U36579 ( .A(n50927), .B(n41296), .Y(n23193) );
  XNOR2XL U36580 ( .A(n51000), .B(n36792), .Y(n20254) );
  XNOR2XL U36581 ( .A(n50987), .B(n36790), .Y(n19593) );
  XNOR2XL U36582 ( .A(n51002), .B(n36799), .Y(n20194) );
  XNOR2XL U36583 ( .A(n50978), .B(n36797), .Y(n19643) );
  XNOR2XL U36584 ( .A(n50943), .B(n36789), .Y(n21087) );
  XNOR2XL U36585 ( .A(n50951), .B(n41294), .Y(n23508) );
  XNOR2XL U36586 ( .A(n50988), .B(n36789), .Y(n19603) );
  XNOR2XL U36587 ( .A(n50967), .B(n36799), .Y(n19715) );
  XNOR2XL U36588 ( .A(n50958), .B(n36795), .Y(n19766) );
  XNOR2XL U36589 ( .A(n50998), .B(n36796), .Y(n20234) );
  XNOR2XL U36590 ( .A(n50921), .B(n41293), .Y(n22973) );
  XNOR2XL U36591 ( .A(n50957), .B(n36795), .Y(n19746) );
  XNOR2XL U36592 ( .A(n50976), .B(n36790), .Y(n19846) );
  XNOR2XL U36593 ( .A(n50966), .B(n36791), .Y(n19705) );
  XNOR2XL U36594 ( .A(n50955), .B(n36793), .Y(n21016) );
  XNOR2XL U36595 ( .A(n50977), .B(n36798), .Y(n19633) );
  XNOR2XL U36596 ( .A(n50923), .B(n41294), .Y(n22953) );
  XNOR2XL U36597 ( .A(n50956), .B(n36798), .Y(n21006) );
  XNOR2XL U36598 ( .A(n50942), .B(n36797), .Y(n21117) );
  XNOR2XL U36599 ( .A(n50975), .B(n36796), .Y(n19816) );
  XNOR2XL U36600 ( .A(n50973), .B(n36795), .Y(n19836) );
  XNOR2XL U36601 ( .A(n50920), .B(n41293), .Y(n22993) );
  XNOR2XL U36602 ( .A(n50941), .B(n36789), .Y(n21107) );
  XNOR2XL U36603 ( .A(n50970), .B(n36791), .Y(n19665) );
  XNOR2XL U36604 ( .A(n50918), .B(n41295), .Y(n23013) );
  XNOR2XL U36605 ( .A(n50940), .B(n36791), .Y(n19957) );
  XNOR2XL U36606 ( .A(n50953), .B(n36795), .Y(n21026) );
  XNOR2XL U36607 ( .A(n50954), .B(n36792), .Y(n21037) );
  XNOR2XL U36608 ( .A(n50971), .B(n36798), .Y(n19675) );
  XNOR2XL U36609 ( .A(n50969), .B(n36796), .Y(n19654) );
  XNOR2XL U36610 ( .A(n50985), .B(n36799), .Y(n19573) );
  XNOR2XL U36611 ( .A(n50925), .B(n36798), .Y(n19987) );
  XNOR2XL U36612 ( .A(n50923), .B(n36799), .Y(n21591) );
  XNOR2XL U36613 ( .A(n50916), .B(n41292), .Y(n22923) );
  XNOR2XL U36614 ( .A(n50951), .B(n36790), .Y(n20965) );
  XNOR2XL U36615 ( .A(n50986), .B(n36798), .Y(n19583) );
  XNOR2XL U36616 ( .A(n50926), .B(n36795), .Y(n19977) );
  XNOR2XL U36617 ( .A(n50939), .B(n36796), .Y(n19947) );
  XNOR2XL U36618 ( .A(n50974), .B(n36795), .Y(n19826) );
  XNOR2XL U36619 ( .A(n50919), .B(n41297), .Y(n23003) );
  XNOR2XL U36620 ( .A(n50972), .B(n36799), .Y(n19685) );
  XNOR2XL U36621 ( .A(n50952), .B(n36797), .Y(n20975) );
  XNOR2XL U36622 ( .A(n50965), .B(n36790), .Y(n19695) );
  XNOR2XL U36623 ( .A(n50922), .B(n36793), .Y(n21581) );
  XNOR2XL U36624 ( .A(n50921), .B(n36789), .Y(n21571) );
  XNOR2XL U36625 ( .A(n50917), .B(n41291), .Y(n22983) );
  XNOR2XL U36626 ( .A(n50938), .B(n36797), .Y(n19937) );
  XNOR2XL U36627 ( .A(n50936), .B(n36798), .Y(n19907) );
  XNOR2XL U36628 ( .A(n50919), .B(n36798), .Y(n21491) );
  XNOR2XL U36629 ( .A(n50949), .B(n36791), .Y(n20996) );
  XNOR2XL U36630 ( .A(n50917), .B(n36790), .Y(n21521) );
  XNOR2XL U36631 ( .A(n50937), .B(n36791), .Y(n19927) );
  XNOR2XL U36632 ( .A(n50950), .B(n36793), .Y(n20986) );
  XNOR2XL U36633 ( .A(n50933), .B(n36793), .Y(n19887) );
  XNOR2XL U36634 ( .A(n50935), .B(n36797), .Y(n19917) );
  XNOR2XL U36635 ( .A(n51352), .B(n36867), .Y(n31575) );
  XNOR2XL U36636 ( .A(n50711), .B(n42590), .Y(n31571) );
  XNOR2XL U36637 ( .A(n51138), .B(n42550), .Y(n31560) );
  XNOR2XL U36638 ( .A(n51133), .B(n42550), .Y(n31380) );
  XNOR2XL U36639 ( .A(n51348), .B(n42644), .Y(n31365) );
  XNOR2XL U36640 ( .A(n51346), .B(n42637), .Y(n31335) );
  XNOR2XL U36641 ( .A(n50705), .B(n42588), .Y(n31331) );
  XNOR2XL U36642 ( .A(n50702), .B(n34450), .Y(n31421) );
  XNOR2XL U36643 ( .A(n51343), .B(n42639), .Y(n31425) );
  XNOR2XL U36644 ( .A(n51132), .B(n42552), .Y(n31320) );
  XNOR2XL U36645 ( .A(n51338), .B(n42641), .Y(n31185) );
  XNOR2XL U36646 ( .A(n51344), .B(n42639), .Y(n31455) );
  XNOR2XL U36647 ( .A(n50697), .B(n42588), .Y(n31181) );
  XNOR2XL U36648 ( .A(n50703), .B(n42590), .Y(n31451) );
  XNOR2XL U36649 ( .A(n50699), .B(n42588), .Y(n31271) );
  XNOR2XL U36650 ( .A(n51340), .B(n42638), .Y(n31275) );
  XNOR2XL U36651 ( .A(n50700), .B(n42590), .Y(n31481) );
  XNOR2XL U36652 ( .A(n51341), .B(n42639), .Y(n31485) );
  XNOR2XL U36653 ( .A(n51130), .B(n42550), .Y(n31440) );
  XNOR2XL U36654 ( .A(n51129), .B(n42550), .Y(n31410) );
  XNOR2XL U36655 ( .A(n50762), .B(n42502), .Y(n29063) );
  XNOR2XL U36656 ( .A(n50720), .B(n42502), .Y(n28552) );
  XNOR2XL U36657 ( .A(n37251), .B(n36875), .Y(n31372) );
  XNOR2XL U36658 ( .A(n50493), .B(n42720), .Y(n31342) );
  XNOR2XL U36659 ( .A(n50714), .B(n42501), .Y(n28462) );
  XNOR2XL U36660 ( .A(n50717), .B(n42501), .Y(n28342) );
  XNOR2XL U36661 ( .A(n50710), .B(n42499), .Y(n31561) );
  XNOR2XL U36662 ( .A(n51133), .B(n42626), .Y(n31330) );
  XNOR2XL U36663 ( .A(n50490), .B(n42717), .Y(n31432) );
  XNOR2XL U36664 ( .A(n50703), .B(n42508), .Y(n31291) );
  XNOR2XL U36665 ( .A(n50492), .B(n36728), .Y(n31334) );
  XNOR2XL U36666 ( .A(n51130), .B(n42633), .Y(n31420) );
  XNOR2XL U36667 ( .A(n50491), .B(n42717), .Y(n31462) );
  XNOR2XL U36668 ( .A(n50486), .B(n42720), .Y(n31192) );
  XNOR2XL U36669 ( .A(n50489), .B(n36903), .Y(n31424) );
  XNOR2XL U36670 ( .A(n37252), .B(n42720), .Y(n31282) );
  XNOR2XL U36671 ( .A(n51131), .B(n42626), .Y(n31450) );
  XNOR2XL U36672 ( .A(n51125), .B(n42633), .Y(n31180) );
  XNOR2XL U36673 ( .A(n50704), .B(n42505), .Y(n31321) );
  XNOR2XL U36674 ( .A(n50488), .B(n42717), .Y(n31492) );
  XNOR2XL U36675 ( .A(n50485), .B(n42680), .Y(n31184) );
  XNOR2XL U36676 ( .A(n50490), .B(n41380), .Y(n31454) );
  XNOR2XL U36677 ( .A(n51127), .B(n42628), .Y(n31270) );
  XNOR2XL U36678 ( .A(n50487), .B(n42680), .Y(n31274) );
  XNOR2XL U36679 ( .A(n50489), .B(n41287), .Y(n31522) );
  XNOR2XL U36680 ( .A(n51128), .B(n42633), .Y(n31480) );
  XNOR2XL U36681 ( .A(n50487), .B(n42720), .Y(n31252) );
  XNOR2XL U36682 ( .A(n50485), .B(n42720), .Y(n31222) );
  XNOR2XL U36683 ( .A(n37252), .B(n36903), .Y(n31484) );
  XNOR2XL U36684 ( .A(n50702), .B(n42505), .Y(n31441) );
  XNOR2XL U36685 ( .A(n50701), .B(n42505), .Y(n31411) );
  XNOR2XL U36686 ( .A(n51129), .B(n42628), .Y(n31510) );
  XNOR2XL U36687 ( .A(n51126), .B(n42630), .Y(n31240) );
  XNOR2XL U36688 ( .A(n51148), .B(n41333), .Y(n23254) );
  XNOR2XL U36689 ( .A(n51147), .B(n41331), .Y(n23244) );
  XNOR2XL U36690 ( .A(n50720), .B(n36856), .Y(n23255) );
  XNOR2XL U36691 ( .A(n50719), .B(n36860), .Y(n23245) );
  XNOR2XL U36692 ( .A(n51190), .B(n42549), .Y(n29062) );
  XNOR2XL U36693 ( .A(n50713), .B(n36730), .Y(n28432) );
  XNOR2XL U36694 ( .A(n50920), .B(net219330), .Y(n31337) );
  XNOR2XL U36695 ( .A(n51134), .B(n41283), .Y(n31338) );
  XNOR2XL U36696 ( .A(n50706), .B(net219450), .Y(n31339) );
  XNOR2XL U36697 ( .A(n50918), .B(net219310), .Y(n31457) );
  XNOR2XL U36698 ( .A(n51132), .B(n41281), .Y(n31458) );
  XNOR2XL U36699 ( .A(n50704), .B(net219450), .Y(n31459) );
  XNOR2XL U36700 ( .A(n50916), .B(net219330), .Y(n31517) );
  XNOR2XL U36701 ( .A(n51130), .B(n41281), .Y(n31518) );
  XNOR2XL U36702 ( .A(n50702), .B(net219450), .Y(n31519) );
  XOR2XL U36703 ( .A(n42186), .B(n36809), .Y(n23167) );
  XOR2XL U36704 ( .A(n42103), .B(n42493), .Y(n20392) );
  XOR2XL U36705 ( .A(n42102), .B(n42493), .Y(n20402) );
  XOR2XL U36706 ( .A(n42181), .B(n36807), .Y(n23137) );
  XOR2XL U36707 ( .A(n42182), .B(n36814), .Y(n23157) );
  XOR2XL U36708 ( .A(n42153), .B(n36811), .Y(n24171) );
  XOR2XL U36709 ( .A(n42157), .B(n36811), .Y(n23542) );
  XOR2XL U36710 ( .A(n42135), .B(n36816), .Y(n22390) );
  XOR2XL U36711 ( .A(n42145), .B(n36816), .Y(n24089) );
  XOR2XL U36712 ( .A(n42170), .B(n36811), .Y(n23452) );
  XOR2XL U36713 ( .A(n42108), .B(n42480), .Y(n20218) );
  XOR2XL U36714 ( .A(n42118), .B(n42492), .Y(n20166) );
  XOR2XL U36715 ( .A(n42116), .B(n42492), .Y(n20146) );
  XOR2XL U36716 ( .A(n42159), .B(n36815), .Y(n235620) );
  XOR2XL U36717 ( .A(n42171), .B(n36813), .Y(n23482) );
  XOR2XL U36718 ( .A(n42121), .B(n42492), .Y(n20126) );
  XOR2XL U36719 ( .A(n42106), .B(n42480), .Y(n20270) );
  XOR2XL U36720 ( .A(n42107), .B(n42480), .Y(n20280) );
  XOR2XL U36721 ( .A(n42119), .B(n42492), .Y(n20176) );
  XOR2XL U36722 ( .A(n42162), .B(n36807), .Y(n23522) );
  XOR2XL U36723 ( .A(n42169), .B(n36816), .Y(n23462) );
  XOR2XL U36724 ( .A(n42137), .B(n36811), .Y(n22330) );
  XOR2XL U36725 ( .A(n42130), .B(n42480), .Y(n19567) );
  XOR2XL U36726 ( .A(n42160), .B(n36814), .Y(n23502) );
  XOR2XL U36727 ( .A(n42132), .B(n42478), .Y(n19617) );
  XOR2XL U36728 ( .A(n42131), .B(n42480), .Y(n19557) );
  XOR2XL U36729 ( .A(n42109), .B(n42480), .Y(n20208) );
  XOR2XL U36730 ( .A(n42113), .B(n42480), .Y(n20248) );
  XOR2XL U36731 ( .A(n42122), .B(n42492), .Y(n20136) );
  XOR2XL U36732 ( .A(n42146), .B(n36810), .Y(n24069) );
  XOR2XL U36733 ( .A(n42151), .B(n42489), .Y(n19780) );
  XOR2XL U36734 ( .A(n42153), .B(n42489), .Y(n19760) );
  XOR2XL U36735 ( .A(n42115), .B(n42480), .Y(n20228) );
  XOR2XL U36736 ( .A(n42144), .B(n42489), .Y(n19729) );
  XOR2XL U36737 ( .A(n42111), .B(n42480), .Y(n20187) );
  XOR2XL U36738 ( .A(n42123), .B(n42492), .Y(n20105) );
  XOR2XL U36739 ( .A(n42112), .B(n42480), .Y(n20258) );
  XOR2XL U36740 ( .A(n42185), .B(n36809), .Y(n23197) );
  XOR2XL U36741 ( .A(n42133), .B(n42478), .Y(n19627) );
  XOR2XL U36742 ( .A(n42110), .B(n42480), .Y(n20198) );
  XOR2XL U36743 ( .A(n42134), .B(n42480), .Y(n19647) );
  XOR2XL U36744 ( .A(n42124), .B(n42492), .Y(n19607) );
  XOR2XL U36745 ( .A(n42125), .B(n42492), .Y(n19597) );
  XOR2XL U36746 ( .A(n42154), .B(n42489), .Y(n19770) );
  XOR2XL U36747 ( .A(n42169), .B(n42484), .Y(n21091) );
  XOR2XL U36748 ( .A(n42114), .B(n42480), .Y(n20238) );
  XOR2XL U36749 ( .A(n42191), .B(n36811), .Y(n22977) );
  XOR2XL U36750 ( .A(n42184), .B(n42491), .Y(n20012) );
  XOR2XL U36751 ( .A(n42136), .B(n42490), .Y(n19850) );
  XOR2XL U36752 ( .A(n42161), .B(n36807), .Y(n23512) );
  XOR2XL U36753 ( .A(n42145), .B(n42489), .Y(n19719) );
  XOR2XL U36754 ( .A(n42146), .B(n42489), .Y(n19709) );
  XOR2XL U36755 ( .A(n42155), .B(n42489), .Y(n19750) );
  XOR2XL U36756 ( .A(n42189), .B(n36810), .Y(n22957) );
  XOR2XL U36757 ( .A(n42157), .B(n42483), .Y(n21020) );
  XOR2XL U36758 ( .A(n42156), .B(n42484), .Y(n21010) );
  XOR2XL U36759 ( .A(n42170), .B(n42484), .Y(n21121) );
  XOR2XL U36760 ( .A(n42135), .B(n42480), .Y(n19637) );
  XOR2XL U36761 ( .A(n42137), .B(n42490), .Y(n19820) );
  XOR2XL U36762 ( .A(n42139), .B(n42490), .Y(n19840) );
  XOR2XL U36763 ( .A(n42142), .B(n42489), .Y(n19669) );
  XOR2XL U36764 ( .A(n42192), .B(n36810), .Y(n22997) );
  XOR2XL U36765 ( .A(n42172), .B(n42491), .Y(n19961) );
  XOR2XL U36766 ( .A(n42171), .B(n42484), .Y(n21111) );
  XOR2XL U36767 ( .A(n42194), .B(n36808), .Y(n23017) );
  XOR2XL U36768 ( .A(n42158), .B(n42483), .Y(n21041) );
  XOR2XL U36769 ( .A(n42159), .B(n42483), .Y(n21030) );
  XOR2XL U36770 ( .A(n42141), .B(n42489), .Y(n19679) );
  XOR2XL U36771 ( .A(n42126), .B(n42480), .Y(n19587) );
  XOR2XL U36772 ( .A(n42186), .B(n42491), .Y(n19981) );
  XOR2XL U36773 ( .A(n42143), .B(n42492), .Y(n19658) );
  XOR2XL U36774 ( .A(n42127), .B(n42479), .Y(n19577) );
  XOR2XL U36775 ( .A(n42187), .B(n42491), .Y(n19991) );
  XOR2XL U36776 ( .A(n42138), .B(n42490), .Y(n19830) );
  XOR2XL U36777 ( .A(n42193), .B(n36817), .Y(n23007) );
  XOR2XL U36778 ( .A(n42189), .B(n42483), .Y(n21595) );
  XOR2XL U36779 ( .A(n42196), .B(n36809), .Y(n22927) );
  XOR2XL U36780 ( .A(n42140), .B(n42489), .Y(n19689) );
  XOR2XL U36781 ( .A(n42161), .B(n42483), .Y(n20969) );
  XOR2XL U36782 ( .A(n42173), .B(n42491), .Y(n19951) );
  XOR2XL U36783 ( .A(n42160), .B(n42483), .Y(n20979) );
  XOR2XL U36784 ( .A(n42190), .B(n42490), .Y(n21585) );
  XOR2XL U36785 ( .A(n42147), .B(n42489), .Y(n19699) );
  XOR2XL U36786 ( .A(n42195), .B(n36816), .Y(n22987) );
  XOR2XL U36787 ( .A(n42174), .B(n42491), .Y(n19941) );
  XOR2XL U36788 ( .A(n42191), .B(n42486), .Y(n21575) );
  XOR2XL U36789 ( .A(n42176), .B(n42490), .Y(n19911) );
  XOR2XL U36790 ( .A(n42193), .B(n42486), .Y(n21495) );
  XOR2XL U36791 ( .A(n42163), .B(n42483), .Y(n21000) );
  XOR2XL U36792 ( .A(n42162), .B(n42483), .Y(n20990) );
  XNOR2XL U36793 ( .A(n50500), .B(n42584), .Y(n28465) );
  XNOR2XL U36794 ( .A(n50931), .B(n42543), .Y(n28340) );
  XNOR2XL U36795 ( .A(n50924), .B(n42538), .Y(n31559) );
  XNOR2XL U36796 ( .A(n50917), .B(n42537), .Y(n31289) );
  XNOR2XL U36797 ( .A(n50918), .B(n42537), .Y(n31319) );
  XNOR2XL U36798 ( .A(n50916), .B(n42538), .Y(n31439) );
  XNOR2XL U36799 ( .A(n50915), .B(n42538), .Y(n31409) );
  XNOR2XL U36800 ( .A(n50934), .B(n41291), .Y(n23253) );
  XNOR2XL U36801 ( .A(n50933), .B(n41293), .Y(n23243) );
  XNOR2XL U36802 ( .A(n50976), .B(n42534), .Y(n29061) );
  XOR2XL U36803 ( .A(n42178), .B(n36814), .Y(n23257) );
  XOR2XL U36804 ( .A(n42177), .B(n36813), .Y(n23267) );
  XOR2XL U36805 ( .A(n42179), .B(n36813), .Y(n23247) );
  XNOR2XL U36806 ( .A(n51382), .B(n41300), .Y(n23543) );
  XNOR2XL U36807 ( .A(n51394), .B(n41300), .Y(n24090) );
  XNOR2XL U36808 ( .A(n50531), .B(n36784), .Y(n24173) );
  XNOR2XL U36809 ( .A(n50563), .B(n36766), .Y(n20127) );
  XNOR2XL U36810 ( .A(n50506), .B(n36785), .Y(n23258) );
  XNOR2XL U36811 ( .A(n51380), .B(n41300), .Y(n23563) );
  XNOR2XL U36812 ( .A(n50507), .B(n36776), .Y(n23269) );
  XNOR2XL U36813 ( .A(n50514), .B(n36785), .Y(n23453) );
  XNOR2XL U36814 ( .A(n50578), .B(n36767), .Y(n20271) );
  XNOR2XL U36815 ( .A(n50565), .B(n36767), .Y(n20177) );
  XNOR2XL U36816 ( .A(n50513), .B(n36782), .Y(n23483) );
  XNOR2XL U36817 ( .A(n51377), .B(n41303), .Y(n23523) );
  XNOR2XL U36818 ( .A(n50515), .B(n36778), .Y(n23463) );
  XNOR2XL U36819 ( .A(n51430), .B(n36741), .Y(n20209) );
  XNOR2XL U36820 ( .A(n51426), .B(n36749), .Y(n20249) );
  XNOR2XL U36821 ( .A(n51379), .B(n41302), .Y(n23503) );
  XNOR2XL U36822 ( .A(n50562), .B(n36774), .Y(n20137) );
  XNOR2XL U36823 ( .A(n51424), .B(n36744), .Y(n20229) );
  XNOR2XL U36824 ( .A(n50498), .B(n36778), .Y(n23168) );
  XNOR2XL U36825 ( .A(n51393), .B(n41302), .Y(n24070) );
  XNOR2XL U36826 ( .A(n51428), .B(n36749), .Y(n20189) );
  XNOR2XL U36827 ( .A(n50531), .B(n36764), .Y(n19761) );
  XNOR2XL U36828 ( .A(n50561), .B(n36771), .Y(n20106) );
  XNOR2XL U36829 ( .A(n51427), .B(n36744), .Y(n20260) );
  XNOR2XL U36830 ( .A(n51373), .B(n36740), .Y(n21062) );
  XNOR2XL U36831 ( .A(n51429), .B(n36744), .Y(n20199) );
  XNOR2XL U36832 ( .A(n51436), .B(n36750), .Y(n20393) );
  XNOR2XL U36833 ( .A(n50499), .B(n36783), .Y(n23198) );
  XNOR2XL U36834 ( .A(n51437), .B(n36743), .Y(n20403) );
  XNOR2XL U36835 ( .A(n50503), .B(n36779), .Y(n23138) );
  XNOR2XL U36836 ( .A(n51425), .B(n36747), .Y(n20239) );
  XNOR2XL U36837 ( .A(n51372), .B(n36749), .Y(n21052) );
  XNOR2XL U36838 ( .A(n50530), .B(n36773), .Y(n19771) );
  XNOR2XL U36839 ( .A(n50515), .B(n36773), .Y(n21092) );
  XNOR2XL U36840 ( .A(n51348), .B(n41302), .Y(n22978) );
  XNOR2XL U36841 ( .A(n50500), .B(n36765), .Y(n20014) );
  XNOR2XL U36842 ( .A(n51403), .B(n36749), .Y(n19851) );
  XNOR2XL U36843 ( .A(n50499), .B(n36774), .Y(n20003) );
  XNOR2XL U36844 ( .A(n51378), .B(n41303), .Y(n23513) );
  XNOR2XL U36845 ( .A(n51350), .B(n41303), .Y(n22958) );
  XNOR2XL U36846 ( .A(n51382), .B(n36750), .Y(n21021) );
  XNOR2XL U36847 ( .A(n51402), .B(n36750), .Y(n19821) );
  XNOR2XL U36848 ( .A(n50545), .B(n36770), .Y(n19841) );
  XNOR2XL U36849 ( .A(n51404), .B(n36750), .Y(n19638) );
  XNOR2XL U36850 ( .A(n51347), .B(n41299), .Y(n22998) );
  XNOR2XL U36851 ( .A(n50512), .B(n36772), .Y(n19962) );
  XNOR2XL U36852 ( .A(n51345), .B(n41303), .Y(n23018) );
  XNOR2XL U36853 ( .A(n50513), .B(n36770), .Y(n21112) );
  XNOR2XL U36854 ( .A(n51381), .B(n36747), .Y(n21042) );
  XNOR2XL U36855 ( .A(n50498), .B(n36767), .Y(n19982) );
  XNOR2XL U36856 ( .A(n50497), .B(n36770), .Y(n19993) );
  XNOR2XL U36857 ( .A(n50546), .B(n36770), .Y(n19831) );
  XNOR2XL U36858 ( .A(n51346), .B(n41304), .Y(n23008) );
  XNOR2XL U36859 ( .A(n51380), .B(n36742), .Y(n21032) );
  XNOR2XL U36860 ( .A(n51343), .B(n41300), .Y(n22928) );
  XNOR2XL U36861 ( .A(n51366), .B(n36750), .Y(n19952) );
  XNOR2XL U36862 ( .A(n51378), .B(n36746), .Y(n20970) );
  XNOR2XL U36863 ( .A(n50544), .B(n36773), .Y(n19690) );
  XNOR2XL U36864 ( .A(n51379), .B(n36748), .Y(n20981) );
  XNOR2XL U36865 ( .A(n51349), .B(n36748), .Y(n21586) );
  XNOR2XL U36866 ( .A(n51344), .B(n41303), .Y(n22988) );
  XNOR2XL U36867 ( .A(n51365), .B(n36741), .Y(n19942) );
  XNOR2XL U36868 ( .A(n51347), .B(n36742), .Y(n21506) );
  XNOR2XL U36869 ( .A(n51363), .B(n36740), .Y(n19912) );
  XNOR2XL U36870 ( .A(n51348), .B(n36744), .Y(n21576) );
  XNOR2XL U36871 ( .A(n51346), .B(n36749), .Y(n21496) );
  XNOR2XL U36872 ( .A(n51376), .B(n36749), .Y(n21001) );
  XNOR2XL U36873 ( .A(n51377), .B(n36749), .Y(n20991) );
  XNOR2XL U36874 ( .A(n51364), .B(n36741), .Y(n19932) );
  XNOR2XL U36875 ( .A(n50497), .B(n36785), .Y(n23178) );
  XNOR2XL U36876 ( .A(n50505), .B(n36786), .Y(n23248) );
  XNOR2XL U36877 ( .A(n50502), .B(n36777), .Y(n23158) );
  XOR2XL U36878 ( .A(n41873), .B(n36757), .Y(n19616) );
  XNOR2XL U36879 ( .A(n50766), .B(n42465), .Y(n19615) );
  XNOR2XL U36880 ( .A(n51194), .B(n36722), .Y(n19614) );
  XOR2XL U36881 ( .A(n41865), .B(n36756), .Y(n19606) );
  XNOR2XL U36882 ( .A(n50774), .B(n42465), .Y(n19605) );
  XNOR2XL U36883 ( .A(n51202), .B(n36717), .Y(n19604) );
  XOR2XL U36884 ( .A(n41897), .B(n36755), .Y(n21009) );
  XNOR2XL U36885 ( .A(n50742), .B(n42460), .Y(n21008) );
  XNOR2XL U36886 ( .A(n51170), .B(n36718), .Y(n21007) );
  XNOR2XL U36887 ( .A(n51405), .B(n36742), .Y(n19648) );
  XNOR2XL U36888 ( .A(n51394), .B(n36750), .Y(n19720) );
  XNOR2XL U36889 ( .A(n51393), .B(n36744), .Y(n19710) );
  XNOR2XL U36890 ( .A(n51397), .B(n36749), .Y(n19670) );
  XNOR2XL U36891 ( .A(n51398), .B(n36747), .Y(n19680) );
  XNOR2XL U36892 ( .A(n51396), .B(n36747), .Y(n19660) );
  XNOR2XL U36893 ( .A(n51392), .B(n36744), .Y(n19700) );
  XNOR2XL U36894 ( .A(n50503), .B(n42583), .Y(n28345) );
  XNOR2XL U36895 ( .A(n50490), .B(n42578), .Y(n31294) );
  XNOR2XL U36896 ( .A(n50491), .B(n42583), .Y(n31324) );
  XNOR2XL U36897 ( .A(n50548), .B(n42576), .Y(n29066) );
  XOR2XL U36898 ( .A(n42188), .B(n36873), .Y(n31563) );
  XOR2XL U36899 ( .A(n42193), .B(n41323), .Y(n31383) );
  XOR2XL U36900 ( .A(n42192), .B(n41321), .Y(n31353) );
  XOR2XL U36901 ( .A(n42194), .B(n41322), .Y(n31323) );
  XOR2XL U36902 ( .A(n42196), .B(n36873), .Y(n31443) );
  XOR2XL U36903 ( .A(n42197), .B(n41323), .Y(n31413) );
  XOR2XL U36904 ( .A(n42202), .B(n36801), .Y(n31173) );
  NAND2XL U36905 ( .A(n10863), .B(n11132), .Y(n11129) );
  XOR2XL U36906 ( .A(n42494), .B(n42100), .Y(n47570) );
  NAND2XL U36907 ( .A(n11990), .B(n11991), .Y(n11987) );
  NAND2XL U36908 ( .A(n10853), .B(n10854), .Y(n11107) );
  NAND2XL U36909 ( .A(n11017), .B(n11018), .Y(n11014) );
  NAND2XL U36910 ( .A(n10553), .B(n10556), .Y(n12055) );
  NAND2XL U36911 ( .A(n11388), .B(n11389), .Y(n11385) );
  INVXL U36912 ( .A(n11984), .Y(net151495) );
  AND2XL U36913 ( .A(n11515), .B(n11516), .Y(n11318) );
  INVXL U36914 ( .A(n12893), .Y(net151448) );
  AOI211X2 U36915 ( .A0(n11998), .A1(n11999), .B0(net171132), .C0(net171134),
        .Y(n11996) );
  NAND2XL U36916 ( .A(n12034), .B(n12035), .Y(n12031) );
  NAND2XL U36917 ( .A(n11074), .B(n11075), .Y(n11071) );
  NAND2XL U36918 ( .A(n12025), .B(n12026), .Y(n12023) );
  NAND2XL U36919 ( .A(n11416), .B(n11417), .Y(n11413) );
  NOR2XL U36920 ( .A(net171550), .B(n37253), .Y(n11400) );
  NAND2XL U36921 ( .A(n11094), .B(n11095), .Y(n11091) );
  NAND2XL U36922 ( .A(n10567), .B(n10566), .Y(n12077) );
  NAND2XL U36923 ( .A(n10845), .B(n10847), .Y(n11101) );
  AND2XL U36924 ( .A(n11204), .B(n40396), .Y(n11102) );
  NAND2XL U36925 ( .A(n10565), .B(n10559), .Y(n12071) );
  AND2XL U36926 ( .A(n12144), .B(n12145), .Y(n12074) );
  INVXL U36927 ( .A(n11052), .Y(net171462) );
  INVXL U36928 ( .A(n12922), .Y(n50103) );
  AND2XL U36929 ( .A(n11509), .B(n11510), .Y(n11361) );
  NAND3XL U36930 ( .A(n10529), .B(net209800), .C(n12026), .Y(n48237) );
  INVXL U36931 ( .A(n12156), .Y(net209784) );
  INVXL U36932 ( .A(n12391), .Y(net171471) );
  AND2XL U36933 ( .A(n11054), .B(n12274), .Y(n48524) );
  XOR2XL U36934 ( .A(n41920), .B(n36761), .Y(n19890) );
  XOR2XL U36935 ( .A(n41918), .B(n36756), .Y(n19920) );
  XOR2XL U36936 ( .A(n41938), .B(n41314), .Y(n22916) );
  XOR2XL U36937 ( .A(n41935), .B(n36754), .Y(n21514) );
  XOR2XL U36938 ( .A(n41919), .B(n36754), .Y(n19900) );
  XOR2XL U36939 ( .A(n41938), .B(n36753), .Y(n21454) );
  XOR2XL U36940 ( .A(n41924), .B(n36755), .Y(n19870) );
  XOR2XL U36941 ( .A(n41922), .B(n36759), .Y(n19880) );
  XOR2XL U36942 ( .A(n41921), .B(n36756), .Y(n19860) );
  XOR2XL U36943 ( .A(n41939), .B(n41311), .Y(n22906) );
  XOR2XL U36944 ( .A(n41923), .B(n36760), .Y(n19970) );
  XOR2XL U36945 ( .A(n41944), .B(n41309), .Y(n22896) );
  XOR2XL U36946 ( .A(n41941), .B(n41311), .Y(n23026) );
  XOR2XL U36947 ( .A(n41939), .B(n36757), .Y(n21484) );
  XOR2XL U36948 ( .A(n41940), .B(n41312), .Y(n22936) );
  XOR2XL U36949 ( .A(n41945), .B(n41313), .Y(n22824) );
  XOR2XL U36950 ( .A(n41943), .B(n41316), .Y(n23036) );
  XOR2XL U36951 ( .A(n41940), .B(n36753), .Y(n21474) );
  XOR2XL U36952 ( .A(n41946), .B(n41316), .Y(n22814) );
  XOR2XL U36953 ( .A(n41941), .B(n36759), .Y(n21554) );
  XOR2XL U36954 ( .A(n41943), .B(n36757), .Y(n21544) );
  XNOR2XL U36955 ( .A(n51337), .B(n42701), .Y(n31794) );
  XNOR2XL U36956 ( .A(n51334), .B(n42701), .Y(n31854) );
  XNOR2XL U36957 ( .A(n51336), .B(n42701), .Y(n31764) );
  XNOR2XL U36958 ( .A(n51335), .B(n42701), .Y(n31884) );
  XNOR2XL U36959 ( .A(n51330), .B(n42701), .Y(n31824) );
  XNOR2XL U36960 ( .A(n51332), .B(n42701), .Y(n31674) );
  XNOR2XL U36961 ( .A(n51333), .B(n42701), .Y(n31704) );
  XNOR2XL U36962 ( .A(n51331), .B(n42701), .Y(n31734) );
  XNOR2XL U36963 ( .A(n51328), .B(n42702), .Y(n31132) );
  XNOR2XL U36964 ( .A(n51329), .B(n42702), .Y(n31162) );
  XOR2XL U36965 ( .A(n41943), .B(n36893), .Y(n31791) );
  XOR2XL U36966 ( .A(n42202), .B(n36880), .Y(n31795) );
  XOR2XL U36967 ( .A(n42203), .B(n42661), .Y(n31787) );
  XOR2XL U36968 ( .A(n41944), .B(n42608), .Y(n31783) );
  XOR2XL U36969 ( .A(n41942), .B(n41318), .Y(n22886) );
  XOR2XL U36970 ( .A(n41946), .B(n36901), .Y(n31851) );
  XOR2XL U36971 ( .A(n42205), .B(n36889), .Y(n31855) );
  XOR2XL U36972 ( .A(n41947), .B(n42608), .Y(n31843) );
  XOR2XL U36973 ( .A(n42206), .B(n42665), .Y(n31847) );
  XOR2XL U36974 ( .A(n41944), .B(n36901), .Y(n31761) );
  XOR2XL U36975 ( .A(n42203), .B(n36882), .Y(n31765) );
  XOR2XL U36976 ( .A(n41945), .B(n42608), .Y(n31753) );
  XOR2XL U36977 ( .A(n42204), .B(n42667), .Y(n31757) );
  XOR2XL U36978 ( .A(n41945), .B(n36897), .Y(n31881) );
  XOR2XL U36979 ( .A(n42204), .B(n36888), .Y(n31885) );
  XOR2XL U36980 ( .A(n41946), .B(n42608), .Y(n31873) );
  XOR2XL U36981 ( .A(n42205), .B(n42665), .Y(n31877) );
  XOR2XL U36982 ( .A(n41950), .B(n36893), .Y(n31821) );
  XOR2XL U36983 ( .A(n42209), .B(n36881), .Y(n31825) );
  XOR2XL U36984 ( .A(n41951), .B(n42608), .Y(n31813) );
  XOR2XL U36985 ( .A(n42210), .B(n42656), .Y(n31817) );
  XOR2XL U36986 ( .A(n41948), .B(n36901), .Y(n31671) );
  XOR2XL U36987 ( .A(n42207), .B(n36887), .Y(n31675) );
  XOR2XL U36988 ( .A(n42208), .B(n42661), .Y(n31667) );
  XOR2XL U36989 ( .A(n41949), .B(n42608), .Y(n31663) );
  XOR2XL U36990 ( .A(n41949), .B(n36893), .Y(n31731) );
  XOR2XL U36991 ( .A(n41947), .B(n36894), .Y(n31701) );
  XOR2XL U36992 ( .A(n42206), .B(n36879), .Y(n31705) );
  XOR2XL U36993 ( .A(n42208), .B(n36885), .Y(n31735) );
  XOR2XL U36994 ( .A(n41950), .B(n42608), .Y(n31723) );
  XOR2XL U36995 ( .A(n42209), .B(n42661), .Y(n31727) );
  XOR2XL U36996 ( .A(n42207), .B(n42667), .Y(n31697) );
  XOR2XL U36997 ( .A(n41948), .B(n42608), .Y(n31693) );
  XOR2XL U36998 ( .A(n41952), .B(n36899), .Y(n31129) );
  XOR2XL U36999 ( .A(n42211), .B(n36881), .Y(n31133) );
  XOR2XL U37000 ( .A(n41951), .B(n36895), .Y(n31159) );
  XOR2XL U37001 ( .A(n42210), .B(n36880), .Y(n31163) );
  XOR2XL U37002 ( .A(n42211), .B(n42656), .Y(n31155) );
  XOR2XL U37003 ( .A(n41952), .B(n42607), .Y(n31151) );
  XOR2XL U37004 ( .A(n41941), .B(n42518), .Y(n31262) );
  XOR2XL U37005 ( .A(n41940), .B(n42519), .Y(n31472) );
  XOR2XL U37006 ( .A(n41939), .B(n42519), .Y(n31502) );
  XOR2XL U37007 ( .A(n41942), .B(n42518), .Y(n31232) );
  XOR2XL U37008 ( .A(n41944), .B(n42518), .Y(n31202) );
  XOR2XL U37009 ( .A(n41946), .B(n42520), .Y(n31743) );
  XOR2XL U37010 ( .A(n41947), .B(n42520), .Y(n31863) );
  XNOR2XL U37011 ( .A(n51129), .B(n41330), .Y(n22914) );
  XNOR2XL U37012 ( .A(n51132), .B(n36716), .Y(n21512) );
  XNOR2XL U37013 ( .A(n51129), .B(n36717), .Y(n21452) );
  XNOR2XL U37014 ( .A(n51143), .B(n36716), .Y(n19868) );
  XNOR2XL U37015 ( .A(n51145), .B(n36718), .Y(n19878) );
  XNOR2XL U37016 ( .A(n51148), .B(n36720), .Y(n19898) );
  XNOR2XL U37017 ( .A(n51146), .B(n36714), .Y(n19858) );
  XNOR2XL U37018 ( .A(n51128), .B(n41328), .Y(n22904) );
  XNOR2XL U37019 ( .A(n51144), .B(n36718), .Y(n19968) );
  XNOR2XL U37020 ( .A(n51123), .B(n41332), .Y(n22894) );
  XNOR2XL U37021 ( .A(n51126), .B(n41331), .Y(n23024) );
  XNOR2XL U37022 ( .A(n51128), .B(n36722), .Y(n21482) );
  XNOR2XL U37023 ( .A(n51127), .B(n41332), .Y(n22934) );
  XNOR2XL U37024 ( .A(n51122), .B(n41327), .Y(n22822) );
  XNOR2XL U37025 ( .A(n51124), .B(n41329), .Y(n23034) );
  XNOR2XL U37026 ( .A(n51127), .B(n36721), .Y(n21472) );
  XNOR2XL U37027 ( .A(n51121), .B(n41331), .Y(n22812) );
  XNOR2XL U37028 ( .A(n51126), .B(n36720), .Y(n21552) );
  XNOR2XL U37029 ( .A(n51124), .B(n36716), .Y(n21542) );
  XNOR2XL U37030 ( .A(n50701), .B(n36856), .Y(n22915) );
  XNOR2XL U37031 ( .A(n50704), .B(n42459), .Y(n21513) );
  XNOR2XL U37032 ( .A(n50720), .B(n42466), .Y(n19899) );
  XNOR2XL U37033 ( .A(n50701), .B(n42459), .Y(n21453) );
  XNOR2XL U37034 ( .A(n50715), .B(n42466), .Y(n19869) );
  XNOR2XL U37035 ( .A(n50717), .B(n42466), .Y(n19879) );
  XNOR2XL U37036 ( .A(n50718), .B(n42466), .Y(n19859) );
  XNOR2XL U37037 ( .A(n50700), .B(n36857), .Y(n22905) );
  XNOR2XL U37038 ( .A(n50716), .B(n42467), .Y(n19969) );
  XNOR2XL U37039 ( .A(n50695), .B(n36852), .Y(n22895) );
  XNOR2XL U37040 ( .A(n50698), .B(n36854), .Y(n23025) );
  XNOR2XL U37041 ( .A(n50700), .B(n42459), .Y(n21483) );
  XNOR2XL U37042 ( .A(n50699), .B(n36854), .Y(n22935) );
  XNOR2XL U37043 ( .A(n50694), .B(n36854), .Y(n22823) );
  XNOR2XL U37044 ( .A(n50696), .B(n36858), .Y(n23035) );
  XNOR2XL U37045 ( .A(n50699), .B(n42459), .Y(n21473) );
  XNOR2XL U37046 ( .A(n50693), .B(n36851), .Y(n22813) );
  XNOR2XL U37047 ( .A(n50698), .B(n42466), .Y(n21553) );
  XNOR2XL U37048 ( .A(n50696), .B(n42459), .Y(n21543) );
  XNOR2XL U37049 ( .A(n50912), .B(n42615), .Y(n31239) );
  XNOR2XL U37050 ( .A(n50910), .B(n42615), .Y(n31209) );
  XNOR2XL U37051 ( .A(n50284), .B(n42708), .Y(n31521) );
  XNOR2XL U37052 ( .A(n50283), .B(n42670), .Y(n31513) );
  XNOR2XL U37053 ( .A(n50280), .B(n42671), .Y(n31243) );
  XNOR2XL U37054 ( .A(n50281), .B(n42704), .Y(n31251) );
  XNOR2XL U37055 ( .A(n50278), .B(n42676), .Y(n31213) );
  XNOR2XL U37056 ( .A(n50279), .B(n42704), .Y(n31221) );
  XNOR2XL U37057 ( .A(n50908), .B(n42617), .Y(n31750) );
  XNOR2XL U37058 ( .A(n50276), .B(n42670), .Y(n31754) );
  XNOR2XL U37059 ( .A(n50277), .B(n41641), .Y(n31762) );
  XNOR2XL U37060 ( .A(n50907), .B(n41284), .Y(n31870) );
  XNOR2XL U37061 ( .A(n50902), .B(n42620), .Y(n31810) );
  XNOR2XL U37062 ( .A(n50275), .B(n36907), .Y(n31874) );
  XNOR2XL U37063 ( .A(n50276), .B(n41642), .Y(n31882) );
  XNOR2XL U37064 ( .A(n50904), .B(n42617), .Y(n31660) );
  XNOR2XL U37065 ( .A(n50270), .B(n42672), .Y(n31814) );
  XNOR2XL U37066 ( .A(n50271), .B(n42706), .Y(n31822) );
  XNOR2XL U37067 ( .A(n50915), .B(n41292), .Y(n22913) );
  XNOR2XL U37068 ( .A(n50918), .B(n36792), .Y(n21511) );
  XNOR2XL U37069 ( .A(n50915), .B(n36791), .Y(n21451) );
  XNOR2XL U37070 ( .A(n50929), .B(n36790), .Y(n19867) );
  XNOR2XL U37071 ( .A(n50931), .B(n36789), .Y(n19877) );
  XNOR2XL U37072 ( .A(n50934), .B(n36799), .Y(n19897) );
  XNOR2XL U37073 ( .A(n50916), .B(n36792), .Y(n21461) );
  XNOR2XL U37074 ( .A(n50932), .B(n36795), .Y(n19857) );
  XNOR2XL U37075 ( .A(n50914), .B(n41290), .Y(n22903) );
  XNOR2XL U37076 ( .A(n50930), .B(n36789), .Y(n19967) );
  XNOR2XL U37077 ( .A(n50909), .B(n41296), .Y(n22893) );
  XNOR2XL U37078 ( .A(n50912), .B(n41294), .Y(n23023) );
  XNOR2XL U37079 ( .A(n50914), .B(n36796), .Y(n21481) );
  XNOR2XL U37080 ( .A(n50913), .B(n41291), .Y(n22933) );
  XNOR2XL U37081 ( .A(n50908), .B(n41291), .Y(n22821) );
  XNOR2XL U37082 ( .A(n50910), .B(n41293), .Y(n23033) );
  XNOR2XL U37083 ( .A(n50913), .B(n36798), .Y(n21471) );
  XNOR2XL U37084 ( .A(n50907), .B(n41293), .Y(n22811) );
  XNOR2XL U37085 ( .A(n50911), .B(n36789), .Y(n21561) );
  XNOR2XL U37086 ( .A(n50912), .B(n36799), .Y(n21551) );
  XNOR2XL U37087 ( .A(n50910), .B(n36791), .Y(n21541) );
  XNOR2XL U37088 ( .A(n51124), .B(n42552), .Y(n31170) );
  XNOR2XL U37089 ( .A(n51342), .B(n42644), .Y(n31515) );
  XNOR2XL U37090 ( .A(n51339), .B(n42637), .Y(n31245) );
  XNOR2XL U37091 ( .A(n50698), .B(n42588), .Y(n31241) );
  XNOR2XL U37092 ( .A(n50701), .B(n34450), .Y(n31511) );
  XNOR2XL U37093 ( .A(n51337), .B(n42641), .Y(n31215) );
  XNOR2XL U37094 ( .A(n50696), .B(n42588), .Y(n31211) );
  XNOR2XL U37095 ( .A(n51126), .B(n42552), .Y(n31260) );
  XNOR2XL U37096 ( .A(n51127), .B(n42550), .Y(n31470) );
  XNOR2XL U37097 ( .A(n51128), .B(n42550), .Y(n31500) );
  XNOR2XL U37098 ( .A(n51125), .B(n42552), .Y(n31230) );
  XNOR2XL U37099 ( .A(n51123), .B(n42552), .Y(n31200) );
  XNOR2XL U37100 ( .A(n51335), .B(n42642), .Y(n31756) );
  XNOR2XL U37101 ( .A(n50694), .B(n36863), .Y(n31752) );
  XNOR2XL U37102 ( .A(n50693), .B(n42589), .Y(n31872) );
  XNOR2XL U37103 ( .A(n51334), .B(n42638), .Y(n31876) );
  XNOR2XL U37104 ( .A(n50688), .B(n42589), .Y(n31812) );
  XNOR2XL U37105 ( .A(n51329), .B(n42638), .Y(n31816) );
  XNOR2XL U37106 ( .A(n51121), .B(n42550), .Y(n31741) );
  XNOR2XL U37107 ( .A(n51124), .B(n42629), .Y(n31210) );
  XNOR2XL U37108 ( .A(n50486), .B(n36903), .Y(n31244) );
  XNOR2XL U37109 ( .A(n50696), .B(n42508), .Y(n31171) );
  XNOR2XL U37110 ( .A(n50488), .B(n36903), .Y(n31514) );
  XNOR2XL U37111 ( .A(n50484), .B(n41379), .Y(n31214) );
  XNOR2XL U37112 ( .A(n50698), .B(n42505), .Y(n31261) );
  XNOR2XL U37113 ( .A(n50699), .B(n42499), .Y(n31471) );
  XNOR2XL U37114 ( .A(n50483), .B(n36709), .Y(n31763) );
  XNOR2XL U37115 ( .A(n50700), .B(n42505), .Y(n31501) );
  XNOR2XL U37116 ( .A(n50697), .B(n42505), .Y(n31231) );
  XNOR2XL U37117 ( .A(n50695), .B(n42505), .Y(n31201) );
  XNOR2XL U37118 ( .A(n51122), .B(n42627), .Y(n31751) );
  XNOR2XL U37119 ( .A(n50482), .B(n36709), .Y(n31883) );
  XNOR2XL U37120 ( .A(n50482), .B(n36903), .Y(n31755) );
  XNOR2XL U37121 ( .A(n50477), .B(n36709), .Y(n31823) );
  XNOR2XL U37122 ( .A(n50694), .B(n42499), .Y(n31772) );
  XNOR2XL U37123 ( .A(n51121), .B(n42626), .Y(n31871) );
  XNOR2XL U37124 ( .A(n50479), .B(n42717), .Y(n31673) );
  XNOR2XL U37125 ( .A(n50481), .B(n36905), .Y(n31875) );
  XNOR2XL U37126 ( .A(n51116), .B(n42629), .Y(n31811) );
  XNOR2XL U37127 ( .A(n50480), .B(n42717), .Y(n31703) );
  XNOR2XL U37128 ( .A(n50478), .B(n42717), .Y(n31733) );
  XNOR2XL U37129 ( .A(n51118), .B(n42625), .Y(n31661) );
  XNOR2XL U37130 ( .A(n50476), .B(n41319), .Y(n31815) );
  XNOR2XL U37131 ( .A(n50691), .B(n34458), .Y(n31832) );
  XNOR2XL U37132 ( .A(n50693), .B(n42499), .Y(n31742) );
  XNOR2XL U37133 ( .A(n50475), .B(n42720), .Y(n31131) );
  XNOR2XL U37134 ( .A(n50909), .B(net219310), .Y(n31758) );
  XNOR2XL U37135 ( .A(n51123), .B(n41282), .Y(n31759) );
  XNOR2XL U37136 ( .A(n50695), .B(net219434), .Y(n31760) );
  XNOR2XL U37137 ( .A(n50908), .B(net258262), .Y(n31878) );
  XNOR2XL U37138 ( .A(n51122), .B(n41281), .Y(n31879) );
  XNOR2XL U37139 ( .A(n50694), .B(net219434), .Y(n31880) );
  XNOR2XL U37140 ( .A(n50904), .B(net219310), .Y(n31728) );
  XNOR2XL U37141 ( .A(n51118), .B(n41283), .Y(n31729) );
  XNOR2XL U37142 ( .A(n50690), .B(net219434), .Y(n31730) );
  XNOR2XL U37143 ( .A(n50906), .B(net219330), .Y(n31698) );
  XNOR2XL U37144 ( .A(n51120), .B(n41283), .Y(n31699) );
  XNOR2XL U37145 ( .A(n50692), .B(net219450), .Y(n31700) );
  XNOR2XL U37146 ( .A(n50901), .B(net219330), .Y(n31126) );
  XNOR2XL U37147 ( .A(n51115), .B(n41282), .Y(n31127) );
  XNOR2XL U37148 ( .A(n50687), .B(net219444), .Y(n31128) );
  XNOR2XL U37149 ( .A(n50902), .B(net219330), .Y(n31156) );
  XNOR2XL U37150 ( .A(n51116), .B(n41282), .Y(n31157) );
  XNOR2XL U37151 ( .A(n50688), .B(net219434), .Y(n31158) );
  XOR2XL U37152 ( .A(n42195), .B(n42486), .Y(n21525) );
  XOR2XL U37153 ( .A(n42175), .B(n42491), .Y(n19931) );
  XOR2XL U37154 ( .A(n42197), .B(n36817), .Y(n22917) );
  XOR2XL U37155 ( .A(n42179), .B(n42490), .Y(n19891) );
  XOR2XL U37156 ( .A(n42177), .B(n42490), .Y(n19921) );
  XOR2XL U37157 ( .A(n42194), .B(n42486), .Y(n21515) );
  XOR2XL U37158 ( .A(n42178), .B(n42490), .Y(n19901) );
  XOR2XL U37159 ( .A(n42196), .B(n42486), .Y(n21465) );
  XOR2XL U37160 ( .A(n42197), .B(n42486), .Y(n21455) );
  XOR2XL U37161 ( .A(n42183), .B(n42490), .Y(n19871) );
  XOR2XL U37162 ( .A(n42181), .B(n42490), .Y(n19881) );
  XOR2XL U37163 ( .A(n42180), .B(n42490), .Y(n19861) );
  XOR2XL U37164 ( .A(n42182), .B(n42491), .Y(n19971) );
  XOR2XL U37165 ( .A(n42198), .B(n36815), .Y(n22907) );
  XOR2XL U37166 ( .A(n42203), .B(n36815), .Y(n22897) );
  XOR2XL U37167 ( .A(n42200), .B(n36808), .Y(n23027) );
  XOR2XL U37168 ( .A(n42201), .B(n36816), .Y(n22887) );
  XOR2XL U37169 ( .A(n42198), .B(n42486), .Y(n21485) );
  XOR2XL U37170 ( .A(n42199), .B(n36815), .Y(n22937) );
  XOR2XL U37171 ( .A(n42204), .B(n36816), .Y(n22825) );
  XOR2XL U37172 ( .A(n42202), .B(n36817), .Y(n23037) );
  XOR2XL U37173 ( .A(n42199), .B(n42486), .Y(n21475) );
  XOR2XL U37174 ( .A(n42205), .B(n36808), .Y(n22815) );
  XOR2XL U37175 ( .A(n42201), .B(n42483), .Y(n21565) );
  XOR2XL U37176 ( .A(n42200), .B(n42484), .Y(n21555) );
  XOR2XL U37177 ( .A(n42202), .B(n42486), .Y(n21545) );
  XNOR2XL U37178 ( .A(n50910), .B(n42537), .Y(n31169) );
  XNOR2XL U37179 ( .A(n50912), .B(n42537), .Y(n31259) );
  XNOR2XL U37180 ( .A(n50913), .B(n42538), .Y(n31469) );
  XNOR2XL U37181 ( .A(n50914), .B(n42538), .Y(n31499) );
  XNOR2XL U37182 ( .A(n50911), .B(n42537), .Y(n31229) );
  XNOR2XL U37183 ( .A(n50909), .B(n42537), .Y(n31199) );
  XNOR2XL U37184 ( .A(n50908), .B(n42538), .Y(n31770) );
  XNOR2XL U37185 ( .A(n50907), .B(n42538), .Y(n31740) );
  XNOR2XL U37186 ( .A(n51344), .B(n36750), .Y(n21526) );
  XNOR2XL U37187 ( .A(n51342), .B(n41301), .Y(n22918) );
  XNOR2XL U37188 ( .A(n50505), .B(n36773), .Y(n19892) );
  XNOR2XL U37189 ( .A(n50507), .B(n36770), .Y(n19922) );
  XNOR2XL U37190 ( .A(n51345), .B(n36747), .Y(n21516) );
  XNOR2XL U37191 ( .A(n50506), .B(n36771), .Y(n19902) );
  XNOR2XL U37192 ( .A(n50501), .B(n36764), .Y(n19872) );
  XNOR2XL U37193 ( .A(n50503), .B(n36767), .Y(n19882) );
  XNOR2XL U37194 ( .A(n50504), .B(n36765), .Y(n19862) );
  XNOR2XL U37195 ( .A(n51341), .B(n41299), .Y(n22908) );
  XNOR2XL U37196 ( .A(n50502), .B(n36774), .Y(n19972) );
  XNOR2XL U37197 ( .A(n50483), .B(n36786), .Y(n22898) );
  XNOR2XL U37198 ( .A(n51339), .B(n41302), .Y(n23028) );
  XNOR2XL U37199 ( .A(n51341), .B(n36750), .Y(n21486) );
  XNOR2XL U37200 ( .A(n51340), .B(n41299), .Y(n22938) );
  XNOR2XL U37201 ( .A(n50482), .B(n36778), .Y(n22826) );
  XNOR2XL U37202 ( .A(n50484), .B(n36785), .Y(n23038) );
  XNOR2XL U37203 ( .A(n51340), .B(n36747), .Y(n21476) );
  XNOR2XL U37204 ( .A(n51338), .B(n36748), .Y(n21566) );
  XNOR2XL U37205 ( .A(n51339), .B(n36746), .Y(n21556) );
  XNOR2XL U37206 ( .A(n50484), .B(n36768), .Y(n21546) );
  XOR2XL U37207 ( .A(n41937), .B(n36760), .Y(n21464) );
  XNOR2XL U37208 ( .A(n50702), .B(n42459), .Y(n21463) );
  XNOR2XL U37209 ( .A(n51130), .B(n36715), .Y(n21462) );
  XOR2XL U37210 ( .A(n41942), .B(n36754), .Y(n21564) );
  XNOR2XL U37211 ( .A(n50697), .B(n42466), .Y(n21563) );
  XNOR2XL U37212 ( .A(n51125), .B(n36714), .Y(n21562) );
  XNOR2XL U37213 ( .A(n50489), .B(n42578), .Y(n31444) );
  XNOR2XL U37214 ( .A(n50488), .B(n42578), .Y(n31414) );
  XNOR2XL U37215 ( .A(n50484), .B(n42578), .Y(n31174) );
  XNOR2XL U37216 ( .A(n50486), .B(n42583), .Y(n31264) );
  XNOR2XL U37217 ( .A(n50487), .B(n42578), .Y(n31474) );
  XNOR2XL U37218 ( .A(n37252), .B(n42578), .Y(n31504) );
  XNOR2XL U37219 ( .A(n50485), .B(n42581), .Y(n31234) );
  XNOR2XL U37220 ( .A(n50483), .B(n42578), .Y(n31204) );
  XNOR2XL U37221 ( .A(n50482), .B(n42578), .Y(n31775) );
  XNOR2XL U37222 ( .A(n50911), .B(n41296), .Y(n22883) );
  XNOR2XL U37223 ( .A(n51125), .B(n41333), .Y(n22884) );
  XNOR2XL U37224 ( .A(n50697), .B(n36858), .Y(n22885) );
  XOR2XL U37225 ( .A(n42200), .B(n36877), .Y(n31263) );
  XOR2XL U37226 ( .A(n42199), .B(n36801), .Y(n31473) );
  XOR2XL U37227 ( .A(n42198), .B(n41321), .Y(n31503) );
  XOR2XL U37228 ( .A(n42201), .B(n41321), .Y(n31233) );
  XOR2XL U37229 ( .A(n42203), .B(n36877), .Y(n31203) );
  XOR2XL U37230 ( .A(n42205), .B(n36801), .Y(n31744) );
  XOR2XL U37231 ( .A(n42206), .B(n41323), .Y(n31864) );
  NAND2XL U37232 ( .A(n48159), .B(n48137), .Y(net210688) );
  NAND2XL U37233 ( .A(net209884), .B(net209927), .Y(n47719) );
  XOR2XL U37234 ( .A(n41947), .B(n41318), .Y(n22865) );
  XOR2XL U37235 ( .A(n41944), .B(n36760), .Y(n21534) );
  XOR2XL U37236 ( .A(n41949), .B(n41317), .Y(n22844) );
  XOR2XL U37237 ( .A(n41948), .B(n41313), .Y(n22804) );
  XOR2XL U37238 ( .A(n41945), .B(n36754), .Y(n21767) );
  XOR2XL U37239 ( .A(n41950), .B(n41317), .Y(n22834) );
  XOR2XL U37240 ( .A(n41948), .B(n36754), .Y(n21747) );
  XOR2XL U37241 ( .A(n41951), .B(n41309), .Y(n22875) );
  XOR2XL U37242 ( .A(n41953), .B(n41310), .Y(n23076) );
  XOR2XL U37243 ( .A(n41950), .B(n36757), .Y(n21707) );
  XOR2XL U37244 ( .A(n41949), .B(n36753), .Y(n21717) );
  XOR2XL U37245 ( .A(n41952), .B(n41318), .Y(n22854) );
  XOR2XL U37246 ( .A(n41954), .B(n41313), .Y(n23066) );
  XOR2XL U37247 ( .A(n41951), .B(n36756), .Y(n21727) );
  XOR2XL U37248 ( .A(n41955), .B(n41314), .Y(n23056) );
  XNOR2XL U37249 ( .A(n51326), .B(n42701), .Y(n31072) );
  XNOR2XL U37250 ( .A(n51327), .B(n42702), .Y(n31102) );
  XNOR2XL U37251 ( .A(n51324), .B(n42695), .Y(n31012) );
  XNOR2XL U37252 ( .A(n51325), .B(n42695), .Y(n31042) );
  XNOR2XL U37253 ( .A(n51322), .B(n42695), .Y(n30952) );
  XNOR2XL U37254 ( .A(n51323), .B(n42695), .Y(n30982) );
  XOR2XL U37255 ( .A(n41953), .B(n36897), .Y(n31099) );
  XOR2XL U37256 ( .A(n42212), .B(n36888), .Y(n31103) );
  XOR2XL U37257 ( .A(n41954), .B(n42611), .Y(n31091) );
  XOR2XL U37258 ( .A(n42213), .B(n42652), .Y(n31095) );
  XOR2XL U37259 ( .A(n41956), .B(n36892), .Y(n31009) );
  XOR2XL U37260 ( .A(n42215), .B(n36888), .Y(n31013) );
  XOR2XL U37261 ( .A(n41957), .B(n36711), .Y(n31001) );
  XOR2XL U37262 ( .A(n42216), .B(n42652), .Y(n31005) );
  XOR2XL U37263 ( .A(n41955), .B(n36891), .Y(n31039) );
  XOR2XL U37264 ( .A(n42214), .B(n36880), .Y(n31043) );
  XOR2XL U37265 ( .A(n42215), .B(n42652), .Y(n31035) );
  XOR2XL U37266 ( .A(n41956), .B(n42608), .Y(n31031) );
  XOR2XL U37267 ( .A(n41958), .B(n36891), .Y(n30949) );
  XOR2XL U37268 ( .A(n42217), .B(n36889), .Y(n30953) );
  XOR2XL U37269 ( .A(n41959), .B(n42606), .Y(n30941) );
  XOR2XL U37270 ( .A(n42218), .B(n42652), .Y(n30945) );
  XOR2XL U37271 ( .A(n41957), .B(n36895), .Y(n30979) );
  XOR2XL U37272 ( .A(n42216), .B(n36886), .Y(n30983) );
  XOR2XL U37273 ( .A(n41958), .B(n36711), .Y(n30971) );
  XOR2XL U37274 ( .A(n42217), .B(n42652), .Y(n30975) );
  XOR2XL U37275 ( .A(n42218), .B(n36879), .Y(n32186) );
  XOR2XL U37276 ( .A(n41959), .B(n36900), .Y(n32182) );
  XOR2XL U37277 ( .A(n42219), .B(n42657), .Y(n32178) );
  XOR2XL U37278 ( .A(n41960), .B(n42605), .Y(n32174) );
  XOR2XL U37279 ( .A(n41950), .B(n42519), .Y(n31653) );
  XOR2XL U37280 ( .A(n41952), .B(n42520), .Y(n31803) );
  XOR2XL U37281 ( .A(n41949), .B(n42520), .Y(n31683) );
  XOR2XL U37282 ( .A(n41953), .B(n42518), .Y(n31141) );
  XOR2XL U37283 ( .A(n41954), .B(n42518), .Y(n31111) );
  XOR2XL U37284 ( .A(n41951), .B(n42520), .Y(n31713) );
  XOR2XL U37285 ( .A(n41956), .B(n42518), .Y(n31051) );
  XOR2XL U37286 ( .A(n41955), .B(n42518), .Y(n31081) );
  XOR2XL U37287 ( .A(n41957), .B(n42518), .Y(n31021) );
  XOR2XL U37288 ( .A(n41958), .B(n42518), .Y(n30991) );
  XNOR2XL U37289 ( .A(n51120), .B(n41332), .Y(n22863) );
  XNOR2XL U37290 ( .A(n51123), .B(n36715), .Y(n21532) );
  XNOR2XL U37291 ( .A(n51120), .B(n36717), .Y(n21695) );
  XNOR2XL U37292 ( .A(n51118), .B(n41330), .Y(n22842) );
  XNOR2XL U37293 ( .A(n51119), .B(n41332), .Y(n22802) );
  XNOR2XL U37294 ( .A(n51122), .B(n36718), .Y(n21765) );
  XNOR2XL U37295 ( .A(n51117), .B(n36913), .Y(n22832) );
  XNOR2XL U37296 ( .A(n51119), .B(n36718), .Y(n21745) );
  XNOR2XL U37297 ( .A(n51116), .B(n41327), .Y(n22873) );
  XNOR2XL U37298 ( .A(n51114), .B(n41328), .Y(n23074) );
  XNOR2XL U37299 ( .A(n51117), .B(n36714), .Y(n21705) );
  XNOR2XL U37300 ( .A(n51118), .B(n36718), .Y(n21715) );
  XNOR2XL U37301 ( .A(n51115), .B(n41333), .Y(n22852) );
  XNOR2XL U37302 ( .A(n51113), .B(n41330), .Y(n23064) );
  XNOR2XL U37303 ( .A(n51116), .B(n36714), .Y(n21725) );
  XNOR2XL U37304 ( .A(n51112), .B(n41331), .Y(n23054) );
  XNOR2XL U37305 ( .A(n51115), .B(n36717), .Y(n21735) );
  XNOR2XL U37306 ( .A(n50692), .B(n36856), .Y(n22864) );
  XNOR2XL U37307 ( .A(n50695), .B(n42459), .Y(n21533) );
  XNOR2XL U37308 ( .A(n50690), .B(n36850), .Y(n22843) );
  XNOR2XL U37309 ( .A(n50691), .B(n36858), .Y(n22803) );
  XNOR2XL U37310 ( .A(n50694), .B(n42462), .Y(n21766) );
  XNOR2XL U37311 ( .A(n50689), .B(n36852), .Y(n22833) );
  XNOR2XL U37312 ( .A(n50691), .B(n42462), .Y(n21746) );
  XNOR2XL U37313 ( .A(n50688), .B(n36859), .Y(n22874) );
  XNOR2XL U37314 ( .A(n50686), .B(n36853), .Y(n23075) );
  XNOR2XL U37315 ( .A(n50689), .B(n42462), .Y(n21706) );
  XNOR2XL U37316 ( .A(n50690), .B(n42462), .Y(n21716) );
  XNOR2XL U37317 ( .A(n50687), .B(n36859), .Y(n22853) );
  XNOR2XL U37318 ( .A(n50685), .B(n36857), .Y(n23065) );
  XNOR2XL U37319 ( .A(n50688), .B(n42462), .Y(n21726) );
  XNOR2XL U37320 ( .A(n50684), .B(n36857), .Y(n23055) );
  XNOR2XL U37321 ( .A(n50272), .B(n42670), .Y(n31664) );
  XNOR2XL U37322 ( .A(n50273), .B(n42711), .Y(n31672) );
  XNOR2XL U37323 ( .A(n50903), .B(n42617), .Y(n31720) );
  XNOR2XL U37324 ( .A(n50905), .B(n42617), .Y(n31690) );
  XNOR2XL U37325 ( .A(n50900), .B(n42616), .Y(n31118) );
  XNOR2XL U37326 ( .A(n50274), .B(n42711), .Y(n31702) );
  XNOR2XL U37327 ( .A(n50271), .B(n42670), .Y(n31724) );
  XNOR2XL U37328 ( .A(n50273), .B(n42670), .Y(n31694) );
  XNOR2XL U37329 ( .A(n50272), .B(n42711), .Y(n31732) );
  XNOR2XL U37330 ( .A(n50901), .B(n42616), .Y(n31148) );
  XNOR2XL U37331 ( .A(n50268), .B(n42670), .Y(n31122) );
  XNOR2XL U37332 ( .A(n50269), .B(n42704), .Y(n31130) );
  XNOR2XL U37333 ( .A(n50270), .B(n42710), .Y(n31160) );
  XNOR2XL U37334 ( .A(n50269), .B(n42676), .Y(n31152) );
  XNOR2XL U37335 ( .A(n50898), .B(n42616), .Y(n31058) );
  XNOR2XL U37336 ( .A(n50266), .B(n42669), .Y(n31062) );
  XNOR2XL U37337 ( .A(n50899), .B(n42615), .Y(n31088) );
  XNOR2XL U37338 ( .A(n50267), .B(n42707), .Y(n31070) );
  XNOR2XL U37339 ( .A(n50267), .B(n42669), .Y(n31092) );
  XNOR2XL U37340 ( .A(n50268), .B(n42710), .Y(n31100) );
  XNOR2XL U37341 ( .A(n50896), .B(n42617), .Y(n30998) );
  XNOR2XL U37342 ( .A(n50897), .B(n42617), .Y(n31028) );
  XNOR2XL U37343 ( .A(n50264), .B(n42676), .Y(n31002) );
  XNOR2XL U37344 ( .A(n50265), .B(n42712), .Y(n31010) );
  XNOR2XL U37345 ( .A(n50266), .B(n42704), .Y(n31040) );
  XNOR2XL U37346 ( .A(n50265), .B(n42670), .Y(n31032) );
  XNOR2XL U37347 ( .A(n50894), .B(n42613), .Y(n30938) );
  XNOR2XL U37348 ( .A(n50896), .B(net219336), .Y(n30976) );
  XNOR2XL U37349 ( .A(n51110), .B(n41281), .Y(n30977) );
  XNOR2XL U37350 ( .A(n50682), .B(net258207), .Y(n30978) );
  XNOR2XL U37351 ( .A(n50906), .B(n41295), .Y(n22862) );
  XNOR2XL U37352 ( .A(n50909), .B(n36793), .Y(n21531) );
  XNOR2XL U37353 ( .A(n50906), .B(n36793), .Y(n21694) );
  XNOR2XL U37354 ( .A(n50904), .B(n41294), .Y(n22841) );
  XNOR2XL U37355 ( .A(n50905), .B(n41296), .Y(n22801) );
  XNOR2XL U37356 ( .A(n50908), .B(n36799), .Y(n21764) );
  XNOR2XL U37357 ( .A(n50903), .B(n41297), .Y(n22831) );
  XNOR2XL U37358 ( .A(n50905), .B(n36793), .Y(n21744) );
  XNOR2XL U37359 ( .A(n50902), .B(n41291), .Y(n22872) );
  XNOR2XL U37360 ( .A(n50900), .B(n41290), .Y(n23073) );
  XNOR2XL U37361 ( .A(n50903), .B(n36795), .Y(n21704) );
  XNOR2XL U37362 ( .A(n50904), .B(n36790), .Y(n21714) );
  XNOR2XL U37363 ( .A(n50901), .B(n41296), .Y(n22851) );
  XNOR2XL U37364 ( .A(n50899), .B(n41292), .Y(n23063) );
  XNOR2XL U37365 ( .A(n50902), .B(n36799), .Y(n21724) );
  XNOR2XL U37366 ( .A(n50898), .B(n41291), .Y(n23053) );
  XNOR2XL U37367 ( .A(n50901), .B(n36789), .Y(n21734) );
  XNOR2XL U37368 ( .A(n51331), .B(n42638), .Y(n31666) );
  XNOR2XL U37369 ( .A(n50690), .B(n36863), .Y(n31662) );
  XNOR2XL U37370 ( .A(n50689), .B(n34450), .Y(n31722) );
  XNOR2XL U37371 ( .A(n51330), .B(n42639), .Y(n31726) );
  XNOR2XL U37372 ( .A(n51332), .B(n36867), .Y(n31696) );
  XNOR2XL U37373 ( .A(n50691), .B(n36863), .Y(n31692) );
  XNOR2XL U37374 ( .A(n51120), .B(n42552), .Y(n31861) );
  XNOR2XL U37375 ( .A(n50686), .B(n42588), .Y(n31120) );
  XNOR2XL U37376 ( .A(n51327), .B(n42641), .Y(n31124) );
  XNOR2XL U37377 ( .A(n51328), .B(n36867), .Y(n31154) );
  XNOR2XL U37378 ( .A(n50687), .B(n42588), .Y(n31150) );
  XNOR2XL U37379 ( .A(n51117), .B(n42550), .Y(n31651) );
  XNOR2XL U37380 ( .A(n51115), .B(n42552), .Y(n31801) );
  XNOR2XL U37381 ( .A(n51118), .B(n42550), .Y(n31681) );
  XNOR2XL U37382 ( .A(n50684), .B(n42588), .Y(n31060) );
  XNOR2XL U37383 ( .A(n51325), .B(n42644), .Y(n31064) );
  XNOR2XL U37384 ( .A(n50685), .B(n42588), .Y(n31090) );
  XNOR2XL U37385 ( .A(n51326), .B(n42637), .Y(n31094) );
  XNOR2XL U37386 ( .A(n51114), .B(n42552), .Y(n31139) );
  XNOR2XL U37387 ( .A(n51113), .B(n42552), .Y(n31109) );
  XNOR2XL U37388 ( .A(n51116), .B(n42550), .Y(n31711) );
  XNOR2XL U37389 ( .A(n50682), .B(n42588), .Y(n31000) );
  XNOR2XL U37390 ( .A(n51323), .B(n36867), .Y(n31004) );
  XNOR2XL U37391 ( .A(n51324), .B(n36867), .Y(n31034) );
  XNOR2XL U37392 ( .A(n50683), .B(n42588), .Y(n31030) );
  XNOR2XL U37393 ( .A(n50679), .B(net219434), .Y(n32151) );
  XNOR2XL U37394 ( .A(n51111), .B(n42552), .Y(n31049) );
  XNOR2XL U37395 ( .A(n51321), .B(n42641), .Y(n30944) );
  XNOR2XL U37396 ( .A(n50677), .B(net219434), .Y(n32091) );
  XNOR2XL U37397 ( .A(n50680), .B(net219442), .Y(n32181) );
  XNOR2XL U37398 ( .A(n50680), .B(n36863), .Y(n30940) );
  XNOR2XL U37399 ( .A(n51112), .B(n42552), .Y(n31079) );
  XNOR2XL U37400 ( .A(n50478), .B(n36903), .Y(n31665) );
  XNOR2XL U37401 ( .A(n50476), .B(n42720), .Y(n31161) );
  XNOR2XL U37402 ( .A(n51117), .B(n42629), .Y(n31721) );
  XNOR2XL U37403 ( .A(n51119), .B(n42628), .Y(n31691) );
  XNOR2XL U37404 ( .A(n51114), .B(n34447), .Y(n31119) );
  XNOR2XL U37405 ( .A(n50477), .B(n41380), .Y(n31725) );
  XNOR2XL U37406 ( .A(n50479), .B(n36903), .Y(n31695) );
  XNOR2XL U37407 ( .A(n51115), .B(n42633), .Y(n31149) );
  XNOR2XL U37408 ( .A(n50474), .B(n42680), .Y(n31123) );
  XNOR2XL U37409 ( .A(n50473), .B(n42720), .Y(n31071) );
  XNOR2XL U37410 ( .A(n50475), .B(n36903), .Y(n31153) );
  XNOR2XL U37411 ( .A(n50474), .B(n42720), .Y(n31101) );
  XNOR2XL U37412 ( .A(n51112), .B(n42632), .Y(n31059) );
  XNOR2XL U37413 ( .A(n50689), .B(n42499), .Y(n31652) );
  XNOR2XL U37414 ( .A(n50687), .B(n34458), .Y(n31802) );
  XNOR2XL U37415 ( .A(n50690), .B(n42499), .Y(n31682) );
  XNOR2XL U37416 ( .A(n50472), .B(n36728), .Y(n31063) );
  XNOR2XL U37417 ( .A(n51113), .B(n42624), .Y(n31089) );
  XNOR2XL U37418 ( .A(n50471), .B(n42720), .Y(n31011) );
  XNOR2XL U37419 ( .A(n50472), .B(n42720), .Y(n31041) );
  XNOR2XL U37420 ( .A(n50473), .B(n41379), .Y(n31093) );
  XNOR2XL U37421 ( .A(n50686), .B(n42505), .Y(n31140) );
  XNOR2XL U37422 ( .A(n51110), .B(n42629), .Y(n30999) );
  XNOR2XL U37423 ( .A(n50685), .B(n42508), .Y(n31110) );
  XNOR2XL U37424 ( .A(n50688), .B(n42499), .Y(n31712) );
  XNOR2XL U37425 ( .A(n51111), .B(n42629), .Y(n31029) );
  XNOR2XL U37426 ( .A(n50470), .B(n36903), .Y(n31003) );
  XNOR2XL U37427 ( .A(n50469), .B(n42724), .Y(n30951) );
  XNOR2XL U37428 ( .A(n50471), .B(n42680), .Y(n31033) );
  XNOR2XL U37429 ( .A(n50470), .B(n42720), .Y(n30981) );
  XNOR2XL U37430 ( .A(n51108), .B(n42628), .Y(n30939) );
  XNOR2XL U37431 ( .A(n50468), .B(n36903), .Y(n30943) );
  XNOR2XL U37432 ( .A(n51106), .B(n34447), .Y(n32142) );
  XNOR2XL U37433 ( .A(n51109), .B(n42633), .Y(n30969) );
  XNOR2XL U37434 ( .A(n50899), .B(net219330), .Y(n31066) );
  XNOR2XL U37435 ( .A(n51113), .B(n41281), .Y(n31067) );
  XNOR2XL U37436 ( .A(n50685), .B(net258207), .Y(n31068) );
  XNOR2XL U37437 ( .A(n50900), .B(n40039), .Y(n31096) );
  XNOR2XL U37438 ( .A(n51114), .B(n41281), .Y(n31097) );
  XNOR2XL U37439 ( .A(n50686), .B(net219434), .Y(n31098) );
  XNOR2XL U37440 ( .A(n50897), .B(net219308), .Y(n31006) );
  XNOR2XL U37441 ( .A(n51111), .B(n41281), .Y(n31007) );
  XNOR2XL U37442 ( .A(n50683), .B(net219434), .Y(n31008) );
  XNOR2XL U37443 ( .A(n50898), .B(n40039), .Y(n31036) );
  XNOR2XL U37444 ( .A(n51112), .B(n41283), .Y(n31037) );
  XNOR2XL U37445 ( .A(n50684), .B(net258207), .Y(n31038) );
  XNOR2XL U37446 ( .A(n50895), .B(net219330), .Y(n30946) );
  XNOR2XL U37447 ( .A(n51109), .B(n41283), .Y(n30947) );
  XNOR2XL U37448 ( .A(n50681), .B(net258207), .Y(n30948) );
  XOR2XL U37449 ( .A(n42206), .B(n36809), .Y(n22866) );
  XOR2XL U37450 ( .A(n42203), .B(n42486), .Y(n21535) );
  XOR2XL U37451 ( .A(n42208), .B(n36808), .Y(n22845) );
  XOR2XL U37452 ( .A(n42207), .B(n36809), .Y(n22805) );
  XOR2XL U37453 ( .A(n42204), .B(n42487), .Y(n21768) );
  XOR2XL U37454 ( .A(n42209), .B(n36807), .Y(n22835) );
  XOR2XL U37455 ( .A(n42210), .B(n36813), .Y(n22876) );
  XOR2XL U37456 ( .A(n42207), .B(n42487), .Y(n21748) );
  XOR2XL U37457 ( .A(n42212), .B(n36811), .Y(n23077) );
  XOR2XL U37458 ( .A(n42209), .B(n42487), .Y(n21708) );
  XOR2XL U37459 ( .A(n42208), .B(n42487), .Y(n21718) );
  XOR2XL U37460 ( .A(n42211), .B(n36811), .Y(n22855) );
  XOR2XL U37461 ( .A(n42213), .B(n36808), .Y(n23067) );
  XOR2XL U37462 ( .A(n42210), .B(n42487), .Y(n21728) );
  XOR2XL U37463 ( .A(n42214), .B(n36814), .Y(n23057) );
  XNOR2XL U37464 ( .A(n50906), .B(n42543), .Y(n31860) );
  XNOR2XL U37465 ( .A(n50903), .B(n42538), .Y(n31650) );
  XNOR2XL U37466 ( .A(n50901), .B(n42541), .Y(n31800) );
  XNOR2XL U37467 ( .A(n50904), .B(n42538), .Y(n31680) );
  XNOR2XL U37468 ( .A(n50900), .B(n42537), .Y(n31138) );
  XNOR2XL U37469 ( .A(n50899), .B(n42537), .Y(n31108) );
  XNOR2XL U37470 ( .A(n50902), .B(n42538), .Y(n31710) );
  XNOR2XL U37471 ( .A(n50897), .B(n42537), .Y(n31048) );
  XNOR2XL U37472 ( .A(n50898), .B(n42537), .Y(n31078) );
  XNOR2XL U37473 ( .A(n51333), .B(n41304), .Y(n22867) );
  XNOR2XL U37474 ( .A(n50483), .B(n36764), .Y(n21536) );
  XNOR2XL U37475 ( .A(n51331), .B(n41303), .Y(n22846) );
  XNOR2XL U37476 ( .A(n50482), .B(n36766), .Y(n21769) );
  XNOR2XL U37477 ( .A(n51330), .B(n41303), .Y(n22836) );
  XNOR2XL U37478 ( .A(n51329), .B(n41305), .Y(n22877) );
  XNOR2XL U37479 ( .A(n51332), .B(n36741), .Y(n21749) );
  XNOR2XL U37480 ( .A(n51327), .B(n41299), .Y(n23078) );
  XNOR2XL U37481 ( .A(n51330), .B(n36750), .Y(n21709) );
  XNOR2XL U37482 ( .A(n51328), .B(n41305), .Y(n22857) );
  XNOR2XL U37483 ( .A(n51326), .B(n41301), .Y(n23068) );
  XNOR2XL U37484 ( .A(n51331), .B(n36746), .Y(n21719) );
  XNOR2XL U37485 ( .A(n51329), .B(n36741), .Y(n21729) );
  XNOR2XL U37486 ( .A(n51325), .B(n41301), .Y(n23058) );
  XNOR2XL U37487 ( .A(n50261), .B(n42708), .Y(n32153) );
  XNOR2XL U37488 ( .A(n50467), .B(n41287), .Y(n32154) );
  XNOR2XL U37489 ( .A(n50259), .B(n42707), .Y(n32093) );
  XNOR2XL U37490 ( .A(n50465), .B(n36709), .Y(n32094) );
  XNOR2XL U37491 ( .A(n50262), .B(n42708), .Y(n32183) );
  XNOR2XL U37492 ( .A(n50468), .B(n41287), .Y(n32184) );
  XNOR2XL U37493 ( .A(n51321), .B(n42697), .Y(n32185) );
  XNOR2XL U37494 ( .A(n50481), .B(n42578), .Y(n31745) );
  XNOR2XL U37495 ( .A(n50480), .B(n42579), .Y(n31865) );
  XNOR2XL U37496 ( .A(n50477), .B(n42578), .Y(n31655) );
  XNOR2XL U37497 ( .A(n50478), .B(n42578), .Y(n31685) );
  XNOR2XL U37498 ( .A(n50475), .B(n42579), .Y(n31805) );
  XNOR2XL U37499 ( .A(n50474), .B(n42579), .Y(n31143) );
  XNOR2XL U37500 ( .A(n50476), .B(n42578), .Y(n31715) );
  XNOR2XL U37501 ( .A(n50473), .B(n42578), .Y(n31113) );
  XNOR2XL U37502 ( .A(n50471), .B(n42578), .Y(n31053) );
  XOR2XL U37503 ( .A(n42209), .B(n36877), .Y(n31654) );
  XOR2XL U37504 ( .A(n42208), .B(n36801), .Y(n31684) );
  XOR2XL U37505 ( .A(n42211), .B(n36877), .Y(n31804) );
  XOR2XL U37506 ( .A(n42212), .B(n41321), .Y(n31142) );
  XOR2XL U37507 ( .A(n42210), .B(n41321), .Y(n31714) );
  XOR2XL U37508 ( .A(n42213), .B(n41323), .Y(n31112) );
  XOR2XL U37509 ( .A(n42215), .B(n41322), .Y(n31052) );
  XOR2XL U37510 ( .A(n42214), .B(n36873), .Y(n31082) );
  XOR2XL U37511 ( .A(n42216), .B(n41323), .Y(n31022) );
  XOR2XL U37512 ( .A(n42217), .B(n36877), .Y(n30992) );
  INVXL U37513 ( .A(n11030), .Y(net209172) );
  AND2XL U37514 ( .A(n11200), .B(n11201), .Y(n11124) );
  XOR2XL U37515 ( .A(n41957), .B(n41311), .Y(n23116) );
  XOR2XL U37516 ( .A(n41958), .B(n41311), .Y(n23106) );
  XOR2XL U37517 ( .A(n41959), .B(n41316), .Y(n23096) );
  XOR2XL U37518 ( .A(n41960), .B(n41316), .Y(n23086) );
  XOR2XL U37519 ( .A(n41952), .B(n36759), .Y(n21737) );
  XOR2XL U37520 ( .A(n41954), .B(n36759), .Y(n21131) );
  XOR2XL U37521 ( .A(n41956), .B(n41312), .Y(n23046) );
  XOR2XL U37522 ( .A(n41953), .B(n36759), .Y(n21141) );
  XOR2XL U37523 ( .A(n41955), .B(n36760), .Y(n21161) );
  XOR2XL U37524 ( .A(n41956), .B(n36753), .Y(n21151) );
  XOR2XL U37525 ( .A(n41958), .B(n36759), .Y(n21191) );
  XOR2XL U37526 ( .A(n41961), .B(n41317), .Y(n22713) );
  XOR2XL U37527 ( .A(n41957), .B(n36761), .Y(n21201) );
  XOR2XL U37528 ( .A(n41959), .B(n36753), .Y(n21181) );
  XOR2XL U37529 ( .A(n41962), .B(n41318), .Y(n22703) );
  XOR2XL U37530 ( .A(n41960), .B(n36753), .Y(n21171) );
  XOR2XL U37531 ( .A(n41965), .B(n41318), .Y(n22743) );
  XNOR2XL U37532 ( .A(n51110), .B(n41332), .Y(n23114) );
  XNOR2XL U37533 ( .A(n51109), .B(n41329), .Y(n23104) );
  XNOR2XL U37534 ( .A(n51108), .B(n41331), .Y(n23094) );
  XNOR2XL U37535 ( .A(n51107), .B(n41330), .Y(n23084) );
  XNOR2XL U37536 ( .A(n50682), .B(n36851), .Y(n23115) );
  XNOR2XL U37537 ( .A(n50681), .B(n36853), .Y(n23105) );
  XNOR2XL U37538 ( .A(n50680), .B(n36850), .Y(n23095) );
  XNOR2XL U37539 ( .A(n50679), .B(n36853), .Y(n23085) );
  XNOR2XL U37540 ( .A(n50896), .B(n41294), .Y(n23113) );
  XNOR2XL U37541 ( .A(n50895), .B(n41293), .Y(n23103) );
  XNOR2XL U37542 ( .A(n50894), .B(n41294), .Y(n23093) );
  XNOR2XL U37543 ( .A(n50893), .B(n41293), .Y(n23083) );
  XOR2XL U37544 ( .A(n41961), .B(n36898), .Y(n32122) );
  XOR2XL U37545 ( .A(n42220), .B(n36889), .Y(n32126) );
  XOR2XL U37546 ( .A(n41962), .B(n42605), .Y(n32114) );
  XOR2XL U37547 ( .A(n42221), .B(n42657), .Y(n32118) );
  XOR2XL U37548 ( .A(n41964), .B(n36892), .Y(n32062) );
  XOR2XL U37549 ( .A(n42223), .B(n36883), .Y(n32066) );
  XOR2XL U37550 ( .A(n41965), .B(n42605), .Y(n32054) );
  XOR2XL U37551 ( .A(n42224), .B(n42657), .Y(n32058) );
  XOR2XL U37552 ( .A(n42222), .B(n36886), .Y(n32006) );
  XOR2XL U37553 ( .A(n41963), .B(n36894), .Y(n32002) );
  XOR2XL U37554 ( .A(n42223), .B(n42657), .Y(n31998) );
  XOR2XL U37555 ( .A(n41964), .B(n42605), .Y(n31994) );
  XOR2XL U37556 ( .A(n41965), .B(n36897), .Y(n31942) );
  XOR2XL U37557 ( .A(n42224), .B(n36885), .Y(n31946) );
  XOR2XL U37558 ( .A(n41966), .B(n42605), .Y(n31934) );
  XOR2XL U37559 ( .A(n42225), .B(n42657), .Y(n31938) );
  XOR2XL U37560 ( .A(n41966), .B(n36892), .Y(n32032) );
  XOR2XL U37561 ( .A(n42225), .B(n36886), .Y(n32036) );
  XOR2XL U37562 ( .A(n41967), .B(n42605), .Y(n32024) );
  XOR2XL U37563 ( .A(n42226), .B(n42657), .Y(n32028) );
  XOR2XL U37564 ( .A(n41968), .B(n36899), .Y(n32212) );
  XOR2XL U37565 ( .A(n42227), .B(n36888), .Y(n32216) );
  XOR2XL U37566 ( .A(n41969), .B(n42605), .Y(n32204) );
  XOR2XL U37567 ( .A(n42228), .B(n42657), .Y(n32208) );
  XOR2XL U37568 ( .A(n42226), .B(n36882), .Y(n32246) );
  XOR2XL U37569 ( .A(n41967), .B(n36891), .Y(n32242) );
  XOR2XL U37570 ( .A(n42227), .B(n42657), .Y(n32238) );
  XOR2XL U37571 ( .A(n41968), .B(n42605), .Y(n32234) );
  XOR2XL U37572 ( .A(n41961), .B(n42521), .Y(n32164) );
  XOR2XL U37573 ( .A(n41962), .B(n42521), .Y(n32134) );
  XOR2XL U37574 ( .A(n41959), .B(n42518), .Y(n30961) );
  XOR2XL U37575 ( .A(n41964), .B(n42521), .Y(n32074) );
  XOR2XL U37576 ( .A(n41963), .B(n42521), .Y(n32104) );
  XOR2XL U37577 ( .A(n41965), .B(n42520), .Y(n31984) );
  XOR2XL U37578 ( .A(n41966), .B(n42521), .Y(n32044) );
  XNOR2XL U37579 ( .A(n51113), .B(n36721), .Y(n21129) );
  XNOR2XL U37580 ( .A(n51111), .B(n41327), .Y(n23044) );
  XNOR2XL U37581 ( .A(n51114), .B(n36722), .Y(n21139) );
  XNOR2XL U37582 ( .A(n51112), .B(n36714), .Y(n21159) );
  XNOR2XL U37583 ( .A(n51111), .B(n36717), .Y(n21149) );
  XNOR2XL U37584 ( .A(n51109), .B(n36715), .Y(n21189) );
  XNOR2XL U37585 ( .A(n51106), .B(n41332), .Y(n22711) );
  XNOR2XL U37586 ( .A(n51110), .B(n36715), .Y(n21199) );
  XNOR2XL U37587 ( .A(n51108), .B(n36720), .Y(n21179) );
  XNOR2XL U37588 ( .A(n51105), .B(n41333), .Y(n22701) );
  XNOR2XL U37589 ( .A(n51107), .B(n36720), .Y(n21169) );
  XNOR2XL U37590 ( .A(n51102), .B(n41327), .Y(n22741) );
  XNOR2XL U37591 ( .A(n50687), .B(n42462), .Y(n21736) );
  XNOR2XL U37592 ( .A(n50685), .B(n42460), .Y(n21130) );
  XNOR2XL U37593 ( .A(n50683), .B(n36860), .Y(n23045) );
  XNOR2XL U37594 ( .A(n50686), .B(n42460), .Y(n21140) );
  XNOR2XL U37595 ( .A(n50684), .B(n42465), .Y(n21160) );
  XNOR2XL U37596 ( .A(n50683), .B(n42460), .Y(n21150) );
  XNOR2XL U37597 ( .A(n50681), .B(n42460), .Y(n21190) );
  XNOR2XL U37598 ( .A(n50678), .B(n36856), .Y(n22712) );
  XNOR2XL U37599 ( .A(n50682), .B(n42465), .Y(n21200) );
  XNOR2XL U37600 ( .A(n50680), .B(n42465), .Y(n21180) );
  XNOR2XL U37601 ( .A(n50677), .B(n36851), .Y(n22702) );
  XNOR2XL U37602 ( .A(n50679), .B(n42460), .Y(n21170) );
  XNOR2XL U37603 ( .A(n50674), .B(n36850), .Y(n22742) );
  XNOR2XL U37604 ( .A(n50262), .B(n42671), .Y(n30942) );
  XNOR2XL U37605 ( .A(n50892), .B(n41284), .Y(n32141) );
  XNOR2XL U37606 ( .A(n50263), .B(n42707), .Y(n30950) );
  XNOR2XL U37607 ( .A(n50895), .B(n42613), .Y(n30968) );
  XNOR2XL U37608 ( .A(n50890), .B(n41284), .Y(n32081) );
  XNOR2XL U37609 ( .A(n50260), .B(n42672), .Y(n32145) );
  XNOR2XL U37610 ( .A(n50264), .B(n42709), .Y(n30980) );
  XNOR2XL U37611 ( .A(n50893), .B(n40039), .Y(n32149) );
  XNOR2XL U37612 ( .A(n50263), .B(n42671), .Y(n30972) );
  XNOR2XL U37613 ( .A(n50893), .B(n42618), .Y(n32171) );
  XNOR2XL U37614 ( .A(n50258), .B(n36907), .Y(n32085) );
  XNOR2XL U37615 ( .A(n50891), .B(net219324), .Y(n32089) );
  XNOR2XL U37616 ( .A(n50894), .B(net219310), .Y(n32179) );
  XNOR2XL U37617 ( .A(n50261), .B(n42672), .Y(n32175) );
  XNOR2XL U37618 ( .A(n50891), .B(n41284), .Y(n32111) );
  XNOR2XL U37619 ( .A(n50888), .B(n41284), .Y(n32051) );
  XNOR2XL U37620 ( .A(n50259), .B(n42672), .Y(n32115) );
  XNOR2XL U37621 ( .A(n50892), .B(net219310), .Y(n32119) );
  XNOR2XL U37622 ( .A(n50889), .B(n42614), .Y(n31991) );
  XNOR2XL U37623 ( .A(n50256), .B(n36907), .Y(n32055) );
  XNOR2XL U37624 ( .A(n50889), .B(net219330), .Y(n32059) );
  XNOR2XL U37625 ( .A(n50890), .B(net219310), .Y(n31999) );
  XNOR2XL U37626 ( .A(n50257), .B(n36907), .Y(n31995) );
  XNOR2XL U37627 ( .A(n50887), .B(n41284), .Y(n31931) );
  XNOR2XL U37628 ( .A(n50886), .B(n41284), .Y(n32021) );
  XNOR2XL U37629 ( .A(n50255), .B(n42674), .Y(n31935) );
  XNOR2XL U37630 ( .A(n50888), .B(net219310), .Y(n31939) );
  XNOR2XL U37631 ( .A(n50899), .B(n36797), .Y(n21128) );
  XNOR2XL U37632 ( .A(n50897), .B(n41291), .Y(n23043) );
  XNOR2XL U37633 ( .A(n50900), .B(n36790), .Y(n21138) );
  XNOR2XL U37634 ( .A(n50898), .B(n36790), .Y(n21158) );
  XNOR2XL U37635 ( .A(n50897), .B(n36789), .Y(n21148) );
  XNOR2XL U37636 ( .A(n50895), .B(n36792), .Y(n21188) );
  XNOR2XL U37637 ( .A(n50892), .B(n41296), .Y(n22710) );
  XNOR2XL U37638 ( .A(n50896), .B(n36791), .Y(n21198) );
  XNOR2XL U37639 ( .A(n50894), .B(n36798), .Y(n21178) );
  XNOR2XL U37640 ( .A(n50891), .B(n41296), .Y(n22700) );
  XNOR2XL U37641 ( .A(n50893), .B(n36792), .Y(n21168) );
  XNOR2XL U37642 ( .A(n50888), .B(n41297), .Y(n22740) );
  XNOR2XL U37643 ( .A(n51319), .B(n42641), .Y(n32147) );
  XNOR2XL U37644 ( .A(n50678), .B(n42589), .Y(n32143) );
  XNOR2XL U37645 ( .A(n50681), .B(n34450), .Y(n30970) );
  XNOR2XL U37646 ( .A(n51322), .B(n36867), .Y(n30974) );
  XNOR2XL U37647 ( .A(n51110), .B(n42552), .Y(n31019) );
  XNOR2XL U37648 ( .A(n51109), .B(n42552), .Y(n30989) );
  XNOR2XL U37649 ( .A(n50678), .B(net219442), .Y(n32121) );
  XNOR2XL U37650 ( .A(n50676), .B(n42589), .Y(n32083) );
  XNOR2XL U37651 ( .A(n51317), .B(n42642), .Y(n32087) );
  XNOR2XL U37652 ( .A(n51320), .B(n42641), .Y(n32177) );
  XNOR2XL U37653 ( .A(n50679), .B(n34450), .Y(n32173) );
  XNOR2XL U37654 ( .A(n50675), .B(net219434), .Y(n32061) );
  XNOR2XL U37655 ( .A(n51107), .B(n42549), .Y(n30929) );
  XNOR2XL U37656 ( .A(n50676), .B(net219434), .Y(n32001) );
  XNOR2XL U37657 ( .A(n50677), .B(n42589), .Y(n32113) );
  XNOR2XL U37658 ( .A(n51318), .B(n42643), .Y(n32117) );
  XNOR2XL U37659 ( .A(n51106), .B(n42552), .Y(n32162) );
  XNOR2XL U37660 ( .A(n51105), .B(n42552), .Y(n32132) );
  XNOR2XL U37661 ( .A(n51108), .B(n42553), .Y(n30959) );
  XNOR2XL U37662 ( .A(n50674), .B(n42589), .Y(n32053) );
  XNOR2XL U37663 ( .A(n51315), .B(n42639), .Y(n32057) );
  XNOR2XL U37664 ( .A(n51316), .B(n42642), .Y(n31997) );
  XNOR2XL U37665 ( .A(n50675), .B(n42589), .Y(n31993) );
  XNOR2XL U37666 ( .A(n50674), .B(net219434), .Y(n31941) );
  XNOR2XL U37667 ( .A(n51103), .B(n42552), .Y(n32072) );
  XNOR2XL U37668 ( .A(n50673), .B(net219434), .Y(n32031) );
  XNOR2XL U37669 ( .A(n51104), .B(n42548), .Y(n32102) );
  XNOR2XL U37670 ( .A(n50673), .B(n42589), .Y(n31933) );
  XNOR2XL U37671 ( .A(n51314), .B(n42644), .Y(n31937) );
  XNOR2XL U37672 ( .A(n50671), .B(net219442), .Y(n32211) );
  XNOR2XL U37673 ( .A(n51102), .B(n42552), .Y(n31982) );
  XNOR2XL U37674 ( .A(n50672), .B(net219442), .Y(n32241) );
  XNOR2XL U37675 ( .A(n51101), .B(n42552), .Y(n32042) );
  XNOR2XL U37676 ( .A(n50672), .B(n42589), .Y(n32023) );
  XNOR2XL U37677 ( .A(n51313), .B(n36867), .Y(n32027) );
  XNOR2XL U37678 ( .A(n50684), .B(n42505), .Y(n31080) );
  XNOR2XL U37679 ( .A(n51104), .B(n42633), .Y(n32082) );
  XNOR2XL U37680 ( .A(n50466), .B(n41379), .Y(n32146) );
  XNOR2XL U37681 ( .A(n51107), .B(n41281), .Y(n32150) );
  XNOR2XL U37682 ( .A(n50469), .B(n41380), .Y(n30973) );
  XNOR2XL U37683 ( .A(n50682), .B(n42499), .Y(n31020) );
  XNOR2XL U37684 ( .A(n51107), .B(n42633), .Y(n32172) );
  XNOR2XL U37685 ( .A(n50464), .B(n41379), .Y(n32086) );
  XNOR2XL U37686 ( .A(n50681), .B(n42499), .Y(n30990) );
  XNOR2XL U37687 ( .A(n51105), .B(n41282), .Y(n32090) );
  XNOR2XL U37688 ( .A(n51108), .B(n41281), .Y(n32180) );
  XNOR2XL U37689 ( .A(n50467), .B(n36728), .Y(n32176) );
  XNOR2XL U37690 ( .A(n50679), .B(n42499), .Y(n30930) );
  XNOR2XL U37691 ( .A(n51105), .B(n42628), .Y(n32112) );
  XNOR2XL U37692 ( .A(n51102), .B(n42630), .Y(n32052) );
  XNOR2XL U37693 ( .A(n50465), .B(n41379), .Y(n32116) );
  XNOR2XL U37694 ( .A(n51106), .B(n41282), .Y(n32120) );
  XNOR2XL U37695 ( .A(n50678), .B(n42508), .Y(n32163) );
  XNOR2XL U37696 ( .A(n51103), .B(n42629), .Y(n31992) );
  XNOR2XL U37697 ( .A(n50462), .B(n36903), .Y(n32056) );
  XNOR2XL U37698 ( .A(n50677), .B(n42506), .Y(n32133) );
  XNOR2XL U37699 ( .A(n50680), .B(n42499), .Y(n30960) );
  XNOR2XL U37700 ( .A(n51103), .B(n41281), .Y(n32060) );
  XNOR2XL U37701 ( .A(n51104), .B(n41283), .Y(n32000) );
  XNOR2XL U37702 ( .A(n50463), .B(n41379), .Y(n31996) );
  XNOR2XL U37703 ( .A(n50675), .B(n36737), .Y(n32073) );
  XNOR2XL U37704 ( .A(n51101), .B(n42624), .Y(n31932) );
  XNOR2XL U37705 ( .A(n50461), .B(n36834), .Y(n31936) );
  XNOR2XL U37706 ( .A(n51100), .B(n42631), .Y(n32022) );
  XNOR2XL U37707 ( .A(n50676), .B(n34458), .Y(n32103) );
  XNOR2XL U37708 ( .A(n51102), .B(n41281), .Y(n31940) );
  XNOR2XL U37709 ( .A(n50674), .B(n34458), .Y(n31983) );
  XNOR2XL U37710 ( .A(n50460), .B(n36834), .Y(n32026) );
  XNOR2XL U37711 ( .A(n50673), .B(n42506), .Y(n32043) );
  XOR2XL U37712 ( .A(n42216), .B(n36813), .Y(n23117) );
  XOR2XL U37713 ( .A(n42217), .B(n36811), .Y(n23107) );
  XOR2XL U37714 ( .A(n42218), .B(n36814), .Y(n23097) );
  XOR2XL U37715 ( .A(n42219), .B(n36815), .Y(n23087) );
  XOR2XL U37716 ( .A(n42211), .B(n42487), .Y(n21738) );
  XOR2XL U37717 ( .A(n42213), .B(n42484), .Y(n21132) );
  XOR2XL U37718 ( .A(n42215), .B(n36809), .Y(n23047) );
  XOR2XL U37719 ( .A(n42212), .B(n42484), .Y(n21142) );
  XOR2XL U37720 ( .A(n42214), .B(n42490), .Y(n21162) );
  XOR2XL U37721 ( .A(n42215), .B(n42484), .Y(n21152) );
  XOR2XL U37722 ( .A(n42217), .B(n42490), .Y(n21192) );
  XOR2XL U37723 ( .A(n42220), .B(n36811), .Y(n22714) );
  XOR2XL U37724 ( .A(n42216), .B(n42490), .Y(n21202) );
  XOR2XL U37725 ( .A(n42218), .B(n42484), .Y(n21182) );
  XOR2XL U37726 ( .A(n42221), .B(n36808), .Y(n22704) );
  XOR2XL U37727 ( .A(n42219), .B(n42484), .Y(n21172) );
  XOR2XL U37728 ( .A(n42224), .B(n36814), .Y(n22744) );
  XNOR2XL U37729 ( .A(n50896), .B(n42537), .Y(n31018) );
  XNOR2XL U37730 ( .A(n50895), .B(n42536), .Y(n30988) );
  XNOR2XL U37731 ( .A(n50893), .B(n42536), .Y(n30928) );
  XNOR2XL U37732 ( .A(n50892), .B(n42543), .Y(n32161) );
  XNOR2XL U37733 ( .A(n50891), .B(n42543), .Y(n32131) );
  XNOR2XL U37734 ( .A(n50894), .B(n42536), .Y(n30958) );
  XNOR2XL U37735 ( .A(n50889), .B(n42543), .Y(n32071) );
  XNOR2XL U37736 ( .A(n50890), .B(n42544), .Y(n32101) );
  XNOR2XL U37737 ( .A(n50888), .B(n42543), .Y(n31981) );
  XNOR2XL U37738 ( .A(n50887), .B(n42544), .Y(n32041) );
  XNOR2XL U37739 ( .A(n51328), .B(n36741), .Y(n21739) );
  XNOR2XL U37740 ( .A(n51323), .B(n41300), .Y(n23118) );
  XNOR2XL U37741 ( .A(n51326), .B(n36747), .Y(n21133) );
  XNOR2XL U37742 ( .A(n51324), .B(n41300), .Y(n23048) );
  XNOR2XL U37743 ( .A(n51327), .B(n36750), .Y(n21143) );
  XNOR2XL U37744 ( .A(n51325), .B(n36749), .Y(n21163) );
  XNOR2XL U37745 ( .A(n51324), .B(n36749), .Y(n21153) );
  XNOR2XL U37746 ( .A(n50468), .B(n36779), .Y(n23098) );
  XNOR2XL U37747 ( .A(n50469), .B(n36764), .Y(n21193) );
  XNOR2XL U37748 ( .A(n50466), .B(n36776), .Y(n22715) );
  XNOR2XL U37749 ( .A(n51318), .B(n41305), .Y(n22705) );
  XNOR2XL U37750 ( .A(n51323), .B(n36747), .Y(n21203) );
  XNOR2XL U37751 ( .A(n50468), .B(n36766), .Y(n21183) );
  XNOR2XL U37752 ( .A(n50467), .B(n36776), .Y(n23088) );
  XNOR2XL U37753 ( .A(n51317), .B(n41305), .Y(n22695) );
  XNOR2XL U37754 ( .A(n50467), .B(n36765), .Y(n21173) );
  XNOR2XL U37755 ( .A(n51315), .B(n41304), .Y(n22745) );
  XNOR2XL U37756 ( .A(n50469), .B(n36777), .Y(n23108) );
  XNOR2XL U37757 ( .A(n50260), .B(n42711), .Y(n32123) );
  XNOR2XL U37758 ( .A(n50466), .B(n36709), .Y(n32124) );
  XNOR2XL U37759 ( .A(n51319), .B(n42697), .Y(n32125) );
  XNOR2XL U37760 ( .A(n50257), .B(n41641), .Y(n32063) );
  XNOR2XL U37761 ( .A(n50463), .B(n36709), .Y(n32064) );
  XNOR2XL U37762 ( .A(n51316), .B(n42697), .Y(n32065) );
  XNOR2XL U37763 ( .A(n50258), .B(n41642), .Y(n32003) );
  XNOR2XL U37764 ( .A(n50464), .B(n36709), .Y(n32004) );
  XNOR2XL U37765 ( .A(n51317), .B(n42697), .Y(n32005) );
  XNOR2XL U37766 ( .A(n50256), .B(n41642), .Y(n31943) );
  XNOR2XL U37767 ( .A(n50462), .B(n36709), .Y(n31944) );
  XNOR2XL U37768 ( .A(n51315), .B(n42697), .Y(n31945) );
  XNOR2XL U37769 ( .A(n50255), .B(n41642), .Y(n32033) );
  XNOR2XL U37770 ( .A(n50461), .B(n36709), .Y(n32034) );
  XNOR2XL U37771 ( .A(n51314), .B(n42697), .Y(n32035) );
  XNOR2XL U37772 ( .A(n50253), .B(n42708), .Y(n32213) );
  XNOR2XL U37773 ( .A(n50459), .B(n41287), .Y(n32214) );
  XNOR2XL U37774 ( .A(n51312), .B(n42697), .Y(n32215) );
  XNOR2XL U37775 ( .A(n50254), .B(n42708), .Y(n32243) );
  XNOR2XL U37776 ( .A(n50460), .B(n41287), .Y(n32244) );
  XNOR2XL U37777 ( .A(n51313), .B(n42697), .Y(n32245) );
  XNOR2XL U37778 ( .A(n50472), .B(n42583), .Y(n31083) );
  XNOR2XL U37779 ( .A(n50470), .B(n42582), .Y(n31023) );
  XNOR2XL U37780 ( .A(n50469), .B(n42583), .Y(n30993) );
  XNOR2XL U37781 ( .A(n50467), .B(n42579), .Y(n30933) );
  XNOR2XL U37782 ( .A(n50466), .B(n42579), .Y(n32166) );
  XNOR2XL U37783 ( .A(n50465), .B(n42579), .Y(n32136) );
  XNOR2XL U37784 ( .A(n50468), .B(n42584), .Y(n30963) );
  XNOR2XL U37785 ( .A(n50463), .B(n42581), .Y(n32076) );
  XNOR2XL U37786 ( .A(n50464), .B(n42579), .Y(n32106) );
  XNOR2XL U37787 ( .A(n50462), .B(n42579), .Y(n31986) );
  XOR2XL U37788 ( .A(n42220), .B(n36873), .Y(n32165) );
  XOR2XL U37789 ( .A(n42221), .B(n41321), .Y(n32135) );
  XOR2XL U37790 ( .A(n42218), .B(n36877), .Y(n30962) );
  XOR2XL U37791 ( .A(n42223), .B(n36877), .Y(n32075) );
  XOR2XL U37792 ( .A(n42222), .B(n36801), .Y(n32105) );
  XOR2XL U37793 ( .A(n42224), .B(n36877), .Y(n31985) );
  XOR2XL U37794 ( .A(n42225), .B(n41322), .Y(n32045) );
  NOR2BXL U37795 ( .AN(n13016), .B(n36944), .Y(n11406) );
  INVXL U37796 ( .A(n12323), .Y(net171491) );
  INVXL U37797 ( .A(n11410), .Y(net151750) );
  INVXL U37798 ( .A(n11423), .Y(net151594) );
  AND2XL U37799 ( .A(n12146), .B(n12147), .Y(n12066) );
  XOR2XL U37800 ( .A(n41963), .B(n36759), .Y(n21443) );
  XOR2XL U37801 ( .A(n41964), .B(n41313), .Y(n22683) );
  XOR2XL U37802 ( .A(n41966), .B(n41318), .Y(n22723) );
  XOR2XL U37803 ( .A(n41967), .B(n41310), .Y(n22753) );
  XOR2XL U37804 ( .A(n41964), .B(n36753), .Y(n21433) );
  XOR2XL U37805 ( .A(n41966), .B(n36756), .Y(n21383) );
  XOR2XL U37806 ( .A(n41969), .B(n41311), .Y(n22783) );
  XOR2XL U37807 ( .A(n41965), .B(n36757), .Y(n21393) );
  XOR2XL U37808 ( .A(n41967), .B(n36760), .Y(n21293) );
  XOR2XL U37809 ( .A(n41968), .B(n41312), .Y(n22733) );
  XOR2XL U37810 ( .A(n41970), .B(n41313), .Y(n22773) );
  XOR2XL U37811 ( .A(n41968), .B(n36755), .Y(n21403) );
  XOR2XL U37812 ( .A(n41971), .B(n41316), .Y(n22763) );
  XOR2XL U37813 ( .A(n41973), .B(n41311), .Y(n22663) );
  XNOR2XL U37814 ( .A(n51310), .B(n42697), .Y(n32275) );
  XNOR2XL U37815 ( .A(n51305), .B(n42695), .Y(n30772) );
  XNOR2XL U37816 ( .A(n51303), .B(n42695), .Y(n30712) );
  XNOR2XL U37817 ( .A(n37242), .B(n42695), .Y(n30802) );
  XNOR2XL U37818 ( .A(n51304), .B(n42695), .Y(n30742) );
  XNOR2XL U37819 ( .A(n51306), .B(n42693), .Y(n32335) );
  XOR2XL U37820 ( .A(n41969), .B(n36892), .Y(n32302) );
  XOR2XL U37821 ( .A(n42228), .B(n36883), .Y(n32306) );
  XOR2XL U37822 ( .A(n41970), .B(n42605), .Y(n32294) );
  XOR2XL U37823 ( .A(n42229), .B(n42657), .Y(n32298) );
  XOR2XL U37824 ( .A(n41970), .B(n36900), .Y(n32272) );
  XOR2XL U37825 ( .A(n41971), .B(n42605), .Y(n32264) );
  XOR2XL U37826 ( .A(n42230), .B(n42657), .Y(n32268) );
  XOR2XL U37827 ( .A(n41975), .B(n42605), .Y(n32324) );
  XOR2XL U37828 ( .A(n42234), .B(n42658), .Y(n32328) );
  XOR2XL U37829 ( .A(n41972), .B(n36900), .Y(n32362) );
  XOR2XL U37830 ( .A(n42231), .B(n36885), .Y(n32366) );
  XOR2XL U37831 ( .A(n41973), .B(n42605), .Y(n32354) );
  XOR2XL U37832 ( .A(n42232), .B(n42658), .Y(n32358) );
  XOR2XL U37833 ( .A(n41976), .B(n36895), .Y(n30769) );
  XOR2XL U37834 ( .A(n42235), .B(n36882), .Y(n30773) );
  XOR2XL U37835 ( .A(n41977), .B(n42606), .Y(n30761) );
  XOR2XL U37836 ( .A(n42236), .B(n42652), .Y(n30765) );
  XOR2XL U37837 ( .A(n42230), .B(n36885), .Y(n31916) );
  XOR2XL U37838 ( .A(n41978), .B(n36891), .Y(n30709) );
  XOR2XL U37839 ( .A(n41971), .B(n36892), .Y(n31912) );
  XOR2XL U37840 ( .A(n42231), .B(n42661), .Y(n31908) );
  XOR2XL U37841 ( .A(n41972), .B(n42608), .Y(n31904) );
  XOR2XL U37842 ( .A(n42237), .B(n36881), .Y(n30713) );
  XOR2XL U37843 ( .A(n41979), .B(n36819), .Y(n30701) );
  XOR2XL U37844 ( .A(n42238), .B(n42655), .Y(n30705) );
  XOR2XL U37845 ( .A(n41973), .B(n36901), .Y(n31972) );
  XOR2XL U37846 ( .A(n42232), .B(n36881), .Y(n31976) );
  XOR2XL U37847 ( .A(n41974), .B(n42605), .Y(n31964) );
  XOR2XL U37848 ( .A(n42233), .B(n42657), .Y(n31968) );
  XOR2XL U37849 ( .A(n41975), .B(n36900), .Y(n30799) );
  XOR2XL U37850 ( .A(n42234), .B(n36882), .Y(n30803) );
  XOR2XL U37851 ( .A(n42235), .B(n42652), .Y(n30795) );
  XOR2XL U37852 ( .A(n41976), .B(n42606), .Y(n30791) );
  XOR2XL U37853 ( .A(n41977), .B(n36899), .Y(n30739) );
  XOR2XL U37854 ( .A(n42236), .B(n36880), .Y(n30743) );
  XOR2XL U37855 ( .A(n41978), .B(n36819), .Y(n30731) );
  XOR2XL U37856 ( .A(n42237), .B(n42655), .Y(n30735) );
  XOR2XL U37857 ( .A(n41974), .B(n36900), .Y(n32332) );
  XOR2XL U37858 ( .A(n42233), .B(n36886), .Y(n32336) );
  XOR2XL U37859 ( .A(n41968), .B(n42520), .Y(n32014) );
  XOR2XL U37860 ( .A(n41967), .B(n42520), .Y(n31924) );
  XOR2XL U37861 ( .A(n41969), .B(n42521), .Y(n32224) );
  XOR2XL U37862 ( .A(n41970), .B(n42521), .Y(n32194) );
  XOR2XL U37863 ( .A(n41972), .B(n42521), .Y(n32254) );
  XOR2XL U37864 ( .A(n41971), .B(n42521), .Y(n32284) );
  XOR2XL U37865 ( .A(n41974), .B(n42521), .Y(n32344) );
  XOR2XL U37866 ( .A(n41973), .B(n42520), .Y(n31894) );
  XOR2XL U37867 ( .A(n41976), .B(n42521), .Y(n32314) );
  XNOR2XL U37868 ( .A(n51104), .B(n36722), .Y(n21441) );
  XNOR2XL U37869 ( .A(n51103), .B(n41332), .Y(n22681) );
  XNOR2XL U37870 ( .A(n51101), .B(n41328), .Y(n22721) );
  XNOR2XL U37871 ( .A(n51100), .B(n41333), .Y(n22751) );
  XNOR2XL U37872 ( .A(n51103), .B(n36720), .Y(n21431) );
  XNOR2XL U37873 ( .A(n51101), .B(n36720), .Y(n21381) );
  XNOR2XL U37874 ( .A(n51098), .B(n41327), .Y(n22781) );
  XNOR2XL U37875 ( .A(n51102), .B(n36721), .Y(n21391) );
  XNOR2XL U37876 ( .A(n51100), .B(n36716), .Y(n21291) );
  XNOR2XL U37877 ( .A(n51099), .B(n41330), .Y(n22731) );
  XNOR2XL U37878 ( .A(n51097), .B(n41331), .Y(n22771) );
  XNOR2XL U37879 ( .A(n51099), .B(n36716), .Y(n21401) );
  XNOR2XL U37880 ( .A(n51096), .B(n41331), .Y(n22761) );
  XNOR2XL U37881 ( .A(n51094), .B(n41329), .Y(n22661) );
  XNOR2XL U37882 ( .A(n51095), .B(n41330), .Y(n22791) );
  XNOR2XL U37883 ( .A(n50676), .B(n42459), .Y(n21442) );
  XNOR2XL U37884 ( .A(n50675), .B(n36856), .Y(n22682) );
  XNOR2XL U37885 ( .A(n50673), .B(n36852), .Y(n22722) );
  XNOR2XL U37886 ( .A(n50672), .B(n36859), .Y(n22752) );
  XNOR2XL U37887 ( .A(n50675), .B(n42459), .Y(n21432) );
  XNOR2XL U37888 ( .A(n50673), .B(n42461), .Y(n21382) );
  XNOR2XL U37889 ( .A(n50670), .B(n36857), .Y(n22782) );
  XNOR2XL U37890 ( .A(n50674), .B(n42461), .Y(n21392) );
  XNOR2XL U37891 ( .A(n50672), .B(n42459), .Y(n21292) );
  XNOR2XL U37892 ( .A(n50671), .B(n36850), .Y(n22732) );
  XNOR2XL U37893 ( .A(n50669), .B(n36856), .Y(n22772) );
  XNOR2XL U37894 ( .A(n50671), .B(n42461), .Y(n21402) );
  XNOR2XL U37895 ( .A(n50668), .B(n36859), .Y(n22762) );
  XNOR2XL U37896 ( .A(n50666), .B(n36851), .Y(n22662) );
  XNOR2XL U37897 ( .A(n50667), .B(n36858), .Y(n22792) );
  XNOR2XL U37898 ( .A(n50247), .B(n42707), .Y(n32333) );
  XNOR2XL U37899 ( .A(n50254), .B(n42674), .Y(n32025) );
  XNOR2XL U37900 ( .A(n50887), .B(n40039), .Y(n32029) );
  XNOR2XL U37901 ( .A(n50884), .B(n42615), .Y(n32201) );
  XNOR2XL U37902 ( .A(n50885), .B(n42620), .Y(n32231) );
  XNOR2XL U37903 ( .A(n50252), .B(n42672), .Y(n32205) );
  XNOR2XL U37904 ( .A(n50885), .B(net219310), .Y(n32209) );
  XNOR2XL U37905 ( .A(n50886), .B(net258262), .Y(n32239) );
  XNOR2XL U37906 ( .A(n50253), .B(n42672), .Y(n32235) );
  XNOR2XL U37907 ( .A(n50883), .B(n42617), .Y(n32291) );
  XNOR2XL U37908 ( .A(n50882), .B(n42615), .Y(n32261) );
  XNOR2XL U37909 ( .A(n50251), .B(n42672), .Y(n32295) );
  XNOR2XL U37910 ( .A(n50884), .B(net219308), .Y(n32299) );
  XNOR2XL U37911 ( .A(n50250), .B(n42672), .Y(n32265) );
  XNOR2XL U37912 ( .A(n50883), .B(net219310), .Y(n32269) );
  XNOR2XL U37913 ( .A(n50878), .B(n42613), .Y(n32321) );
  XNOR2XL U37914 ( .A(n50246), .B(n42672), .Y(n32325) );
  XNOR2XL U37915 ( .A(n50881), .B(net219310), .Y(n32359) );
  XNOR2XL U37916 ( .A(n50876), .B(n42613), .Y(n30758) );
  XNOR2XL U37917 ( .A(n50881), .B(n42620), .Y(n31901) );
  XNOR2XL U37918 ( .A(n50874), .B(n42615), .Y(n30698) );
  XNOR2XL U37919 ( .A(n50879), .B(n42619), .Y(n31961) );
  XNOR2XL U37920 ( .A(n50244), .B(n42671), .Y(n30762) );
  XNOR2XL U37921 ( .A(n50882), .B(n36870), .Y(n31909) );
  XNOR2XL U37922 ( .A(n50245), .B(n42712), .Y(n30770) );
  XNOR2XL U37923 ( .A(n50877), .B(n42613), .Y(n30788) );
  XNOR2XL U37924 ( .A(n50249), .B(n36907), .Y(n31905) );
  XNOR2XL U37925 ( .A(n50242), .B(n42671), .Y(n30702) );
  XNOR2XL U37926 ( .A(n50247), .B(n36907), .Y(n31965) );
  XNOR2XL U37927 ( .A(n50243), .B(n42707), .Y(n30710) );
  XNOR2XL U37928 ( .A(n50880), .B(net219336), .Y(n31969) );
  XNOR2XL U37929 ( .A(n50875), .B(n41647), .Y(n30728) );
  XNOR2XL U37930 ( .A(n50246), .B(n42707), .Y(n30800) );
  XNOR2XL U37931 ( .A(n50880), .B(n41284), .Y(n32351) );
  XNOR2XL U37932 ( .A(n50248), .B(n34444), .Y(n32355) );
  XNOR2XL U37933 ( .A(n50890), .B(n36796), .Y(n21440) );
  XNOR2XL U37934 ( .A(n50889), .B(n41295), .Y(n22680) );
  XNOR2XL U37935 ( .A(n50887), .B(n41291), .Y(n22720) );
  XNOR2XL U37936 ( .A(n50886), .B(n41290), .Y(n22750) );
  XNOR2XL U37937 ( .A(n50889), .B(n36792), .Y(n21430) );
  XNOR2XL U37938 ( .A(n50887), .B(n36790), .Y(n21380) );
  XNOR2XL U37939 ( .A(n50884), .B(n41292), .Y(n22780) );
  XNOR2XL U37940 ( .A(n50888), .B(n36791), .Y(n21390) );
  XNOR2XL U37941 ( .A(n50886), .B(n36796), .Y(n21290) );
  XNOR2XL U37942 ( .A(n50885), .B(n41294), .Y(n22730) );
  XNOR2XL U37943 ( .A(n50883), .B(n41293), .Y(n22770) );
  XNOR2XL U37944 ( .A(n50885), .B(n36796), .Y(n21400) );
  XNOR2XL U37945 ( .A(n50882), .B(n41293), .Y(n22760) );
  XNOR2XL U37946 ( .A(n50883), .B(n36793), .Y(n21340) );
  XNOR2XL U37947 ( .A(n50880), .B(n41293), .Y(n22660) );
  XNOR2XL U37948 ( .A(n50881), .B(n41294), .Y(n22790) );
  XNOR2XL U37949 ( .A(n36930), .B(n42720), .Y(n32334) );
  XNOR2XL U37950 ( .A(n50670), .B(net219442), .Y(n32301) );
  XNOR2XL U37951 ( .A(n50670), .B(n36863), .Y(n32203) );
  XNOR2XL U37952 ( .A(n51311), .B(n42641), .Y(n32207) );
  XNOR2XL U37953 ( .A(n51312), .B(n42641), .Y(n32237) );
  XNOR2XL U37954 ( .A(n50671), .B(n36863), .Y(n32233) );
  XNOR2XL U37955 ( .A(n50669), .B(net219442), .Y(n32271) );
  XNOR2XL U37956 ( .A(n51099), .B(n42548), .Y(n32012) );
  XNOR2XL U37957 ( .A(n51100), .B(n42548), .Y(n31922) );
  XNOR2XL U37958 ( .A(n50669), .B(n36863), .Y(n32293) );
  XNOR2XL U37959 ( .A(n51310), .B(n36867), .Y(n32297) );
  XNOR2XL U37960 ( .A(n50667), .B(net219434), .Y(n32361) );
  XNOR2XL U37961 ( .A(n51098), .B(n42547), .Y(n32222) );
  XNOR2XL U37962 ( .A(n50668), .B(n42591), .Y(n32263) );
  XNOR2XL U37963 ( .A(n51309), .B(n42641), .Y(n32267) );
  XNOR2XL U37964 ( .A(n51097), .B(n42547), .Y(n32192) );
  XNOR2XL U37965 ( .A(n50668), .B(net219434), .Y(n31911) );
  XNOR2XL U37966 ( .A(n50666), .B(net219434), .Y(n31971) );
  XNOR2XL U37967 ( .A(n50664), .B(n36863), .Y(n32323) );
  XNOR2XL U37968 ( .A(n51307), .B(n42641), .Y(n32357) );
  XNOR2XL U37969 ( .A(n51304), .B(n42642), .Y(n30764) );
  XNOR2XL U37970 ( .A(n51095), .B(n42547), .Y(n32252) );
  XNOR2XL U37971 ( .A(n51096), .B(n42547), .Y(n32282) );
  XNOR2XL U37972 ( .A(n51302), .B(n36867), .Y(n30704) );
  XNOR2XL U37973 ( .A(n50662), .B(n42592), .Y(n30760) );
  XNOR2XL U37974 ( .A(n51308), .B(n42639), .Y(n31907) );
  XNOR2XL U37975 ( .A(n51305), .B(n42641), .Y(n30794) );
  XNOR2XL U37976 ( .A(n50667), .B(n42589), .Y(n31903) );
  XNOR2XL U37977 ( .A(n50660), .B(n36863), .Y(n30700) );
  XNOR2XL U37978 ( .A(n50665), .B(n42589), .Y(n31963) );
  XNOR2XL U37979 ( .A(n51306), .B(n42638), .Y(n31967) );
  XNOR2XL U37980 ( .A(n51303), .B(n42642), .Y(n30734) );
  XNOR2XL U37981 ( .A(n37242), .B(n36867), .Y(n32327) );
  XNOR2XL U37982 ( .A(n50666), .B(n36865), .Y(n32353) );
  XNOR2XL U37983 ( .A(n51101), .B(n41281), .Y(n32030) );
  XNOR2XL U37984 ( .A(n51098), .B(n42630), .Y(n32202) );
  XNOR2XL U37985 ( .A(n51099), .B(n42631), .Y(n32232) );
  XNOR2XL U37986 ( .A(n50458), .B(n36728), .Y(n32206) );
  XNOR2XL U37987 ( .A(n51099), .B(n41281), .Y(n32210) );
  XNOR2XL U37988 ( .A(n51100), .B(n41282), .Y(n32240) );
  XNOR2XL U37989 ( .A(n50459), .B(n36903), .Y(n32236) );
  XNOR2XL U37990 ( .A(n51097), .B(n42626), .Y(n32292) );
  XNOR2XL U37991 ( .A(n50671), .B(n42506), .Y(n32013) );
  XNOR2XL U37992 ( .A(n50672), .B(n42499), .Y(n31923) );
  XNOR2XL U37993 ( .A(n51096), .B(n42627), .Y(n32262) );
  XNOR2XL U37994 ( .A(n50457), .B(n36903), .Y(n32296) );
  XNOR2XL U37995 ( .A(n51098), .B(n41283), .Y(n32300) );
  XNOR2XL U37996 ( .A(n50670), .B(n42499), .Y(n32223) );
  XNOR2XL U37997 ( .A(n50456), .B(n41380), .Y(n32266) );
  XNOR2XL U37998 ( .A(n50669), .B(n42499), .Y(n32193) );
  XNOR2XL U37999 ( .A(n51097), .B(n41282), .Y(n32270) );
  XNOR2XL U38000 ( .A(n51092), .B(n42632), .Y(n32322) );
  XNOR2XL U38001 ( .A(n50454), .B(n42723), .Y(n30771) );
  XNOR2XL U38002 ( .A(n36931), .B(n42724), .Y(n30711) );
  XNOR2XL U38003 ( .A(n50455), .B(n42724), .Y(n30801) );
  XNOR2XL U38004 ( .A(n50455), .B(n36905), .Y(n32326) );
  XNOR2XL U38005 ( .A(n51095), .B(n41283), .Y(n32360) );
  XNOR2XL U38006 ( .A(n51090), .B(n42631), .Y(n30759) );
  XNOR2XL U38007 ( .A(n50667), .B(n42504), .Y(n32253) );
  XNOR2XL U38008 ( .A(n50668), .B(n42504), .Y(n32283) );
  XNOR2XL U38009 ( .A(n51095), .B(n42627), .Y(n31902) );
  XNOR2XL U38010 ( .A(n51088), .B(n42628), .Y(n30699) );
  XNOR2XL U38011 ( .A(n51093), .B(n42632), .Y(n31962) );
  XNOR2XL U38012 ( .A(n50453), .B(n42724), .Y(n30741) );
  XNOR2XL U38013 ( .A(n50453), .B(n36905), .Y(n30763) );
  XNOR2XL U38014 ( .A(n51096), .B(n41283), .Y(n31910) );
  XNOR2XL U38015 ( .A(n51091), .B(n34447), .Y(n30789) );
  XNOR2XL U38016 ( .A(n37244), .B(n36905), .Y(n30703) );
  XNOR2XL U38017 ( .A(n37243), .B(n41379), .Y(n31906) );
  XNOR2XL U38018 ( .A(n36930), .B(n36905), .Y(n31966) );
  XNOR2XL U38019 ( .A(n51094), .B(n41282), .Y(n31970) );
  XNOR2XL U38020 ( .A(n51089), .B(n42625), .Y(n30729) );
  XNOR2XL U38021 ( .A(n37019), .B(n41319), .Y(n32356) );
  XNOR2XL U38022 ( .A(n51094), .B(n42632), .Y(n32352) );
  XNOR2XL U38023 ( .A(n50879), .B(net219324), .Y(n32329) );
  XNOR2XL U38024 ( .A(n51093), .B(n41281), .Y(n32330) );
  XNOR2XL U38025 ( .A(n50665), .B(net258207), .Y(n32331) );
  XNOR2XL U38026 ( .A(n50877), .B(n40039), .Y(n30766) );
  XNOR2XL U38027 ( .A(n51091), .B(n41283), .Y(n30767) );
  XNOR2XL U38028 ( .A(n50663), .B(net219468), .Y(n30768) );
  XNOR2XL U38029 ( .A(n50875), .B(n40039), .Y(n30706) );
  XNOR2XL U38030 ( .A(n51089), .B(n41281), .Y(n30707) );
  XNOR2XL U38031 ( .A(n50661), .B(net219468), .Y(n30708) );
  XNOR2XL U38032 ( .A(n50878), .B(net219314), .Y(n30796) );
  XNOR2XL U38033 ( .A(n51092), .B(n41281), .Y(n30797) );
  XNOR2XL U38034 ( .A(n50664), .B(net219468), .Y(n30798) );
  XNOR2XL U38035 ( .A(n50876), .B(net219310), .Y(n30736) );
  XNOR2XL U38036 ( .A(n51090), .B(n41281), .Y(n30737) );
  XNOR2XL U38037 ( .A(n50662), .B(net219468), .Y(n30738) );
  XOR2XL U38038 ( .A(n42222), .B(n42486), .Y(n21444) );
  XOR2XL U38039 ( .A(n42223), .B(n36811), .Y(n22684) );
  XOR2XL U38040 ( .A(n42225), .B(n36810), .Y(n22724) );
  XOR2XL U38041 ( .A(n42226), .B(n36811), .Y(n22754) );
  XOR2XL U38042 ( .A(n42223), .B(n42486), .Y(n21434) );
  XOR2XL U38043 ( .A(n42225), .B(n42485), .Y(n21384) );
  XOR2XL U38044 ( .A(n42224), .B(n42485), .Y(n21394) );
  XOR2XL U38045 ( .A(n42226), .B(n42490), .Y(n21294) );
  XOR2XL U38046 ( .A(n42228), .B(n36809), .Y(n22784) );
  XOR2XL U38047 ( .A(n42227), .B(n36810), .Y(n22734) );
  XOR2XL U38048 ( .A(n42229), .B(n36816), .Y(n22774) );
  XOR2XL U38049 ( .A(n42227), .B(n42485), .Y(n21404) );
  XOR2XL U38050 ( .A(n42230), .B(n36807), .Y(n22764) );
  XOR2XL U38051 ( .A(n42229), .B(n42485), .Y(n21344) );
  XNOR2XL U38052 ( .A(n50885), .B(n42533), .Y(n32011) );
  XNOR2XL U38053 ( .A(n50886), .B(n42533), .Y(n31921) );
  XNOR2XL U38054 ( .A(n50884), .B(n42533), .Y(n32221) );
  XNOR2XL U38055 ( .A(n50883), .B(n42533), .Y(n32191) );
  XNOR2XL U38056 ( .A(n50881), .B(n42532), .Y(n32251) );
  XNOR2XL U38057 ( .A(n50882), .B(n42532), .Y(n32281) );
  XNOR2XL U38058 ( .A(n50458), .B(n42579), .Y(n32226) );
  XNOR2XL U38059 ( .A(n50457), .B(n42579), .Y(n32196) );
  XNOR2XL U38060 ( .A(n37243), .B(n42579), .Y(n32256) );
  XNOR2XL U38061 ( .A(n50456), .B(n42579), .Y(n32286) );
  XNOR2XL U38062 ( .A(n51318), .B(n36741), .Y(n21415) );
  XNOR2XL U38063 ( .A(n51316), .B(n41303), .Y(n22685) );
  XNOR2XL U38064 ( .A(n51314), .B(n41302), .Y(n22725) );
  XNOR2XL U38065 ( .A(n51317), .B(n36744), .Y(n21445) );
  XNOR2XL U38066 ( .A(n50466), .B(n36771), .Y(n21425) );
  XNOR2XL U38067 ( .A(n51313), .B(n41299), .Y(n22755) );
  XNOR2XL U38068 ( .A(n51316), .B(n36742), .Y(n21435) );
  XNOR2XL U38069 ( .A(n51314), .B(n36749), .Y(n21385) );
  XNOR2XL U38070 ( .A(n51311), .B(n41300), .Y(n22785) );
  XNOR2XL U38071 ( .A(n51315), .B(n36750), .Y(n21395) );
  XNOR2XL U38072 ( .A(n51313), .B(n36742), .Y(n21295) );
  XNOR2XL U38073 ( .A(n51312), .B(n41302), .Y(n22735) );
  XNOR2XL U38074 ( .A(n51310), .B(n41300), .Y(n22775) );
  XNOR2XL U38075 ( .A(n51309), .B(n41302), .Y(n22765) );
  XNOR2XL U38076 ( .A(n51312), .B(n36747), .Y(n21405) );
  XNOR2XL U38077 ( .A(n51310), .B(n36742), .Y(n21345) );
  XOR2XL U38078 ( .A(n41970), .B(n36761), .Y(n21343) );
  XNOR2XL U38079 ( .A(n50669), .B(n42461), .Y(n21342) );
  XNOR2XL U38080 ( .A(n51097), .B(n36721), .Y(n21341) );
  XNOR2XL U38081 ( .A(n50252), .B(n42708), .Y(n32303) );
  XNOR2XL U38082 ( .A(n50458), .B(n41287), .Y(n32304) );
  XNOR2XL U38083 ( .A(n51311), .B(n42697), .Y(n32305) );
  XNOR2XL U38084 ( .A(n50251), .B(n42708), .Y(n32273) );
  XNOR2XL U38085 ( .A(n50457), .B(n41287), .Y(n32274) );
  XOR2XL U38086 ( .A(n42229), .B(n36882), .Y(n32276) );
  XNOR2XL U38087 ( .A(n50249), .B(n42708), .Y(n32363) );
  XNOR2XL U38088 ( .A(n37243), .B(n41287), .Y(n32364) );
  XNOR2XL U38089 ( .A(n51308), .B(n36871), .Y(n32365) );
  XNOR2XL U38090 ( .A(n50250), .B(n41642), .Y(n31913) );
  XNOR2XL U38091 ( .A(n50456), .B(n36709), .Y(n31914) );
  XNOR2XL U38092 ( .A(n51309), .B(n42697), .Y(n31915) );
  XNOR2XL U38093 ( .A(n50248), .B(n42707), .Y(n31973) );
  XNOR2XL U38094 ( .A(n37019), .B(n36709), .Y(n31974) );
  XNOR2XL U38095 ( .A(n51307), .B(n42697), .Y(n31975) );
  XNOR2XL U38096 ( .A(n50461), .B(n42579), .Y(n32046) );
  XNOR2XL U38097 ( .A(n50459), .B(n42580), .Y(n32016) );
  XNOR2XL U38098 ( .A(n50460), .B(n42579), .Y(n31926) );
  XOR2XL U38099 ( .A(n42227), .B(n36873), .Y(n32015) );
  XOR2XL U38100 ( .A(n42226), .B(n41323), .Y(n31925) );
  XOR2XL U38101 ( .A(n42228), .B(n36877), .Y(n32225) );
  XOR2XL U38102 ( .A(n42229), .B(n41321), .Y(n32195) );
  XOR2XL U38103 ( .A(n42231), .B(n36801), .Y(n32255) );
  XOR2XL U38104 ( .A(n42230), .B(n36801), .Y(n32285) );
  XOR2XL U38105 ( .A(n42232), .B(n36873), .Y(n31895) );
  XOR2XL U38106 ( .A(n42233), .B(n36877), .Y(n32345) );
  XOR2XL U38107 ( .A(n42235), .B(n41322), .Y(n32315) );
  XOR2XL U38108 ( .A(n42236), .B(n41323), .Y(n30782) );
  NAND2XL U38109 ( .A(n12715), .B(n12717), .Y(n12047) );
  INVXL U38110 ( .A(n12303), .Y(net151848) );
  INVXL U38111 ( .A(net209817), .Y(net171247) );
  INVXL U38112 ( .A(n12726), .Y(net151757) );
  INVXL U38113 ( .A(n12306), .Y(net151738) );
  NOR2BXL U38114 ( .AN(n10607), .B(net151741), .Y(n12050) );
  INVXL U38115 ( .A(net210109), .Y(net171550) );
  INVXL U38116 ( .A(n12795), .Y(n49509) );
  NOR2BXL U38117 ( .AN(n48225), .B(n49501), .Y(n12041) );
  XNOR2XL U38118 ( .A(n50872), .B(net219310), .Y(n30886) );
  XNOR2XL U38119 ( .A(n51086), .B(n41281), .Y(n30887) );
  XNOR2XL U38120 ( .A(n50658), .B(net219468), .Y(n30888) );
  XNOR2XL U38121 ( .A(n50650), .B(net219434), .Y(n30557) );
  XNOR2XL U38122 ( .A(n50647), .B(net219434), .Y(n30285) );
  XNOR2XL U38123 ( .A(n50868), .B(net219330), .Y(n30645) );
  XNOR2XL U38124 ( .A(n51082), .B(n41281), .Y(n30646) );
  XNOR2XL U38125 ( .A(n50654), .B(net219468), .Y(n30647) );
  NAND4XL U38126 ( .A(n12795), .B(n12731), .C(n12064), .D(n12065), .Y(n10176)
         );
  XOR2XL U38127 ( .A(n41972), .B(n41314), .Y(n22793) );
  XOR2XL U38128 ( .A(n41969), .B(n36755), .Y(n21353) );
  XOR2XL U38129 ( .A(n41971), .B(n36757), .Y(n21333) );
  XOR2XL U38130 ( .A(n41974), .B(n41316), .Y(n22643) );
  XOR2XL U38131 ( .A(n41975), .B(n41318), .Y(n22653) );
  XOR2XL U38132 ( .A(n41972), .B(n36761), .Y(n21323) );
  XOR2XL U38133 ( .A(n41977), .B(n41318), .Y(n22592) );
  XOR2XL U38134 ( .A(n41978), .B(n41309), .Y(n22582) );
  XOR2XL U38135 ( .A(n41976), .B(n41317), .Y(n22673) );
  XOR2XL U38136 ( .A(n41975), .B(n36755), .Y(n21313) );
  XOR2XL U38137 ( .A(n41973), .B(n36756), .Y(n21373) );
  XOR2XL U38138 ( .A(n41979), .B(n41318), .Y(n22572) );
  XOR2XL U38139 ( .A(n41981), .B(n41318), .Y(n22632) );
  XOR2XL U38140 ( .A(n41976), .B(n36754), .Y(n21303) );
  XOR2XL U38141 ( .A(n41980), .B(n41310), .Y(n22562) );
  XOR2XL U38142 ( .A(n41978), .B(n36755), .Y(n21636) );
  XOR2XL U38143 ( .A(n41979), .B(n36760), .Y(n21626) );
  XOR2XL U38144 ( .A(n41977), .B(n36760), .Y(n21646) );
  XOR2XL U38145 ( .A(n41982), .B(n41316), .Y(n22612) );
  XOR2XL U38146 ( .A(n41980), .B(n36759), .Y(n21616) );
  XOR2XL U38147 ( .A(n41983), .B(n41316), .Y(n22602) );
  XOR2XL U38148 ( .A(n41983), .B(n36760), .Y(n21666) );
  XOR2XL U38149 ( .A(n41986), .B(n41312), .Y(n22521) );
  XOR2XL U38150 ( .A(n41989), .B(n41311), .Y(n22491) );
  XOR2XL U38151 ( .A(n41984), .B(n36759), .Y(n21656) );
  XOR2XL U38152 ( .A(n41987), .B(n41313), .Y(n22511) );
  XOR2XL U38153 ( .A(n41985), .B(n36759), .Y(n21232) );
  XOR2XL U38154 ( .A(n41987), .B(n36760), .Y(n21222) );
  XOR2XL U38155 ( .A(n41988), .B(n36756), .Y(n21212) );
  XOR2XL U38156 ( .A(n41985), .B(n41311), .Y(n22501) );
  XOR2XL U38157 ( .A(n41990), .B(n41318), .Y(n22531) );
  XOR2XL U38158 ( .A(n41982), .B(n36754), .Y(n21676) );
  XOR2XL U38159 ( .A(n41986), .B(n36761), .Y(n21242) );
  XOR2XL U38160 ( .A(n41981), .B(n36753), .Y(n21686) );
  XOR2XL U38161 ( .A(n41984), .B(n41311), .Y(n22622) );
  XOR2XL U38162 ( .A(n41988), .B(n41317), .Y(n22551) );
  XOR2XL U38163 ( .A(n41991), .B(n41314), .Y(n22481) );
  XNOR2XL U38164 ( .A(n51301), .B(n42695), .Y(n30832) );
  XNOR2XL U38165 ( .A(n51299), .B(n42695), .Y(n30922) );
  XNOR2XL U38166 ( .A(n51302), .B(n42695), .Y(n30862) );
  XNOR2XL U38167 ( .A(n51300), .B(n42695), .Y(n30892) );
  XNOR2XL U38168 ( .A(n51295), .B(n42695), .Y(n30681) );
  XNOR2XL U38169 ( .A(n51296), .B(n42697), .Y(n30651) );
  XNOR2XL U38170 ( .A(n51293), .B(n42697), .Y(n30471) );
  XNOR2XL U38171 ( .A(n51287), .B(n42697), .Y(n30259) );
  XNOR2XL U38172 ( .A(n51294), .B(n42697), .Y(n30501) );
  XNOR2XL U38173 ( .A(n51286), .B(n42697), .Y(n30409) );
  XNOR2XL U38174 ( .A(n51285), .B(n42697), .Y(n30439) );
  XNOR2XL U38175 ( .A(n51284), .B(n42697), .Y(n30349) );
  XNOR2XL U38176 ( .A(n51283), .B(n42697), .Y(n30379) );
  XNOR2XL U38177 ( .A(n51292), .B(n42697), .Y(n30561) );
  XNOR2XL U38178 ( .A(n51291), .B(n42697), .Y(n30591) );
  XNOR2XL U38179 ( .A(n51290), .B(n42697), .Y(n30319) );
  XNOR2XL U38180 ( .A(n51289), .B(n42697), .Y(n30289) );
  XOR2XL U38181 ( .A(n41980), .B(n36895), .Y(n30829) );
  XOR2XL U38182 ( .A(n42239), .B(n36879), .Y(n30833) );
  XOR2XL U38183 ( .A(n41981), .B(n42608), .Y(n30821) );
  XOR2XL U38184 ( .A(n42240), .B(n42657), .Y(n30825) );
  XOR2XL U38185 ( .A(n41982), .B(n36891), .Y(n30919) );
  XOR2XL U38186 ( .A(n42241), .B(n36879), .Y(n30923) );
  XOR2XL U38187 ( .A(n41979), .B(n36901), .Y(n30859) );
  XOR2XL U38188 ( .A(n41983), .B(n42608), .Y(n30911) );
  XOR2XL U38189 ( .A(n42242), .B(n42652), .Y(n30915) );
  XOR2XL U38190 ( .A(n42238), .B(n36883), .Y(n30863) );
  XOR2XL U38191 ( .A(n41980), .B(n42607), .Y(n30851) );
  XOR2XL U38192 ( .A(n42239), .B(n42657), .Y(n30855) );
  XOR2XL U38193 ( .A(n41981), .B(n36895), .Y(n30889) );
  XOR2XL U38194 ( .A(n42240), .B(n36883), .Y(n30893) );
  XOR2XL U38195 ( .A(n42241), .B(n42652), .Y(n30885) );
  XOR2XL U38196 ( .A(n41982), .B(n36711), .Y(n30881) );
  XOR2XL U38197 ( .A(n41984), .B(n36894), .Y(n30618) );
  XOR2XL U38198 ( .A(n41983), .B(n36897), .Y(n30528) );
  XOR2XL U38199 ( .A(n42243), .B(n36879), .Y(n30622) );
  XOR2XL U38200 ( .A(n41985), .B(n36819), .Y(n30610) );
  XOR2XL U38201 ( .A(n42244), .B(n42655), .Y(n30614) );
  XOR2XL U38202 ( .A(n42242), .B(n36883), .Y(n30532) );
  XOR2XL U38203 ( .A(n41984), .B(n36819), .Y(n30520) );
  XOR2XL U38204 ( .A(n42243), .B(n42655), .Y(n30524) );
  XOR2XL U38205 ( .A(n41986), .B(n36899), .Y(n30678) );
  XOR2XL U38206 ( .A(n42245), .B(n36880), .Y(n30682) );
  XOR2XL U38207 ( .A(n41987), .B(n36819), .Y(n30670) );
  XOR2XL U38208 ( .A(n42246), .B(n42655), .Y(n30674) );
  XOR2XL U38209 ( .A(n41985), .B(n36894), .Y(n30648) );
  XOR2XL U38210 ( .A(n42244), .B(n36880), .Y(n30652) );
  XOR2XL U38211 ( .A(n41986), .B(n36819), .Y(n30640) );
  XOR2XL U38212 ( .A(n42245), .B(n42655), .Y(n30644) );
  XOR2XL U38213 ( .A(n41988), .B(n36898), .Y(n30468) );
  XOR2XL U38214 ( .A(n42247), .B(n36887), .Y(n30472) );
  XOR2XL U38215 ( .A(n41989), .B(n36819), .Y(n30460) );
  XOR2XL U38216 ( .A(n42248), .B(n42655), .Y(n30464) );
  XOR2XL U38217 ( .A(n41987), .B(n36898), .Y(n30498) );
  XOR2XL U38218 ( .A(n42246), .B(n36888), .Y(n30502) );
  XOR2XL U38219 ( .A(n42247), .B(n42655), .Y(n30494) );
  XOR2XL U38220 ( .A(n41988), .B(n36819), .Y(n30490) );
  XOR2XL U38221 ( .A(n41995), .B(n36897), .Y(n30406) );
  XOR2XL U38222 ( .A(n42254), .B(n36883), .Y(n30410) );
  XOR2XL U38223 ( .A(n42255), .B(n42655), .Y(n30402) );
  XOR2XL U38224 ( .A(n41996), .B(n36819), .Y(n30398) );
  XOR2XL U38225 ( .A(n41996), .B(n36892), .Y(n30436) );
  XOR2XL U38226 ( .A(n42255), .B(n36883), .Y(n30440) );
  XOR2XL U38227 ( .A(n42256), .B(n42655), .Y(n30432) );
  XOR2XL U38228 ( .A(n41997), .B(n36819), .Y(n30428) );
  XOR2XL U38229 ( .A(n41998), .B(n36899), .Y(n30376) );
  XOR2XL U38230 ( .A(n42257), .B(n36888), .Y(n30380) );
  XOR2XL U38231 ( .A(n41989), .B(n36897), .Y(n30558) );
  XOR2XL U38232 ( .A(n42248), .B(n36882), .Y(n30562) );
  XOR2XL U38233 ( .A(n42249), .B(n42655), .Y(n30554) );
  XOR2XL U38234 ( .A(n41990), .B(n36819), .Y(n30550) );
  XOR2XL U38235 ( .A(n41990), .B(n36895), .Y(n30588) );
  XOR2XL U38236 ( .A(n42249), .B(n36887), .Y(n30592) );
  XOR2XL U38237 ( .A(n42250), .B(n42655), .Y(n30584) );
  XOR2XL U38238 ( .A(n41991), .B(n36819), .Y(n30580) );
  XNOR2XL U38239 ( .A(n50450), .B(n36780), .Y(n22523) );
  XNOR2XL U38240 ( .A(n50447), .B(n36777), .Y(n22493) );
  XNOR2XL U38241 ( .A(n50449), .B(n36777), .Y(n22513) );
  XNOR2XL U38242 ( .A(n50446), .B(n36780), .Y(n22533) );
  XNOR2XL U38243 ( .A(n50448), .B(n36782), .Y(n22553) );
  XNOR2XL U38244 ( .A(n50445), .B(n36782), .Y(n22483) );
  XOR2XL U38245 ( .A(n41977), .B(n42517), .Y(n30781) );
  XOR2XL U38246 ( .A(n41975), .B(n42520), .Y(n31954) );
  XOR2XL U38247 ( .A(n41978), .B(n42517), .Y(n30751) );
  XOR2XL U38248 ( .A(n41980), .B(n42517), .Y(n30691) );
  XOR2XL U38249 ( .A(n41979), .B(n42517), .Y(n30721) );
  XOR2XL U38250 ( .A(n41981), .B(n42517), .Y(n30841) );
  XOR2XL U38251 ( .A(n41982), .B(n42517), .Y(n30811) );
  XOR2XL U38252 ( .A(n41984), .B(n42517), .Y(n30901) );
  XOR2XL U38253 ( .A(n41983), .B(n42517), .Y(n30871) );
  XOR2XL U38254 ( .A(n41986), .B(n42517), .Y(n30600) );
  XOR2XL U38255 ( .A(n41985), .B(n42516), .Y(n30510) );
  XOR2XL U38256 ( .A(n41989), .B(n42516), .Y(n30480) );
  XOR2XL U38257 ( .A(n41992), .B(n42516), .Y(n30570) );
  XOR2XL U38258 ( .A(n41993), .B(n42516), .Y(n30298) );
  XOR2XL U38259 ( .A(n41991), .B(n42516), .Y(n30540) );
  XOR2XL U38260 ( .A(n41990), .B(n42516), .Y(n30450) );
  XOR2XL U38261 ( .A(n41987), .B(n42517), .Y(n30630) );
  XOR2XL U38262 ( .A(n41988), .B(n42517), .Y(n30660) );
  XOR2XL U38263 ( .A(n41994), .B(n42516), .Y(n30268) );
  XNOR2XL U38264 ( .A(n51098), .B(n36714), .Y(n21351) );
  XNOR2XL U38265 ( .A(n51096), .B(n36717), .Y(n21331) );
  XNOR2XL U38266 ( .A(n51093), .B(n41332), .Y(n22641) );
  XNOR2XL U38267 ( .A(n51092), .B(n41327), .Y(n22651) );
  XNOR2XL U38268 ( .A(n51095), .B(n36715), .Y(n21321) );
  XNOR2XL U38269 ( .A(n51090), .B(n41330), .Y(n22590) );
  XNOR2XL U38270 ( .A(n51089), .B(n41328), .Y(n22580) );
  XNOR2XL U38271 ( .A(n51091), .B(n41332), .Y(n22671) );
  XNOR2XL U38272 ( .A(n51092), .B(n36722), .Y(n21311) );
  XNOR2XL U38273 ( .A(n51094), .B(n36720), .Y(n21371) );
  XNOR2XL U38274 ( .A(n51088), .B(n41328), .Y(n22570) );
  XNOR2XL U38275 ( .A(n51086), .B(n41333), .Y(n22630) );
  XNOR2XL U38276 ( .A(n51091), .B(n36714), .Y(n21301) );
  XNOR2XL U38277 ( .A(n51087), .B(n41327), .Y(n22560) );
  XNOR2XL U38278 ( .A(n51089), .B(n36714), .Y(n21634) );
  XNOR2XL U38279 ( .A(n51088), .B(n36715), .Y(n21624) );
  XNOR2XL U38280 ( .A(n51090), .B(n36716), .Y(n21644) );
  XNOR2XL U38281 ( .A(n51085), .B(n41332), .Y(n22610) );
  XNOR2XL U38282 ( .A(n51087), .B(n36721), .Y(n21614) );
  XNOR2XL U38283 ( .A(n51084), .B(n36913), .Y(n22600) );
  XNOR2XL U38284 ( .A(n51084), .B(n36720), .Y(n21664) );
  XNOR2XL U38285 ( .A(n51081), .B(n41330), .Y(n22519) );
  XNOR2XL U38286 ( .A(n51078), .B(n41327), .Y(n22489) );
  XNOR2XL U38287 ( .A(n51083), .B(n36721), .Y(n21654) );
  XNOR2XL U38288 ( .A(n51080), .B(n41331), .Y(n22509) );
  XNOR2XL U38289 ( .A(n51082), .B(n36715), .Y(n21230) );
  XNOR2XL U38290 ( .A(n51080), .B(n36718), .Y(n21220) );
  XNOR2XL U38291 ( .A(n51079), .B(n36722), .Y(n21210) );
  XNOR2XL U38292 ( .A(n51082), .B(n41331), .Y(n22499) );
  XNOR2XL U38293 ( .A(n51077), .B(n41332), .Y(n22529) );
  XNOR2XL U38294 ( .A(n51085), .B(n36720), .Y(n21674) );
  XNOR2XL U38295 ( .A(n51081), .B(n36717), .Y(n21240) );
  XNOR2XL U38296 ( .A(n51086), .B(n36717), .Y(n21684) );
  XNOR2XL U38297 ( .A(n51083), .B(n41329), .Y(n22620) );
  XNOR2XL U38298 ( .A(n51079), .B(n41333), .Y(n22549) );
  XNOR2XL U38299 ( .A(n51077), .B(n36721), .Y(n21260) );
  XNOR2XL U38300 ( .A(n51076), .B(n41330), .Y(n22479) );
  XNOR2XL U38301 ( .A(n50670), .B(n42461), .Y(n21352) );
  XNOR2XL U38302 ( .A(n50668), .B(n42461), .Y(n21332) );
  XNOR2XL U38303 ( .A(n50665), .B(n36852), .Y(n22642) );
  XNOR2XL U38304 ( .A(n50664), .B(n36860), .Y(n22652) );
  XNOR2XL U38305 ( .A(n50667), .B(n42461), .Y(n21322) );
  XNOR2XL U38306 ( .A(n50662), .B(n36857), .Y(n22591) );
  XNOR2XL U38307 ( .A(n50661), .B(n36860), .Y(n22581) );
  XNOR2XL U38308 ( .A(n50663), .B(n36854), .Y(n22672) );
  XNOR2XL U38309 ( .A(n50664), .B(n42461), .Y(n21312) );
  XNOR2XL U38310 ( .A(n50666), .B(n42461), .Y(n21372) );
  XNOR2XL U38311 ( .A(n50660), .B(n36851), .Y(n22571) );
  XNOR2XL U38312 ( .A(n50658), .B(n36858), .Y(n22631) );
  XNOR2XL U38313 ( .A(n50663), .B(n42461), .Y(n21302) );
  XNOR2XL U38314 ( .A(n50659), .B(n36854), .Y(n22561) );
  XNOR2XL U38315 ( .A(n50661), .B(n42466), .Y(n21635) );
  XNOR2XL U38316 ( .A(n50660), .B(n42466), .Y(n21625) );
  XNOR2XL U38317 ( .A(n50662), .B(n42466), .Y(n21645) );
  XNOR2XL U38318 ( .A(n50657), .B(n36859), .Y(n22611) );
  XNOR2XL U38319 ( .A(n50659), .B(n42466), .Y(n21615) );
  XNOR2XL U38320 ( .A(n50656), .B(n36853), .Y(n22601) );
  XNOR2XL U38321 ( .A(n50656), .B(n42466), .Y(n21665) );
  XNOR2XL U38322 ( .A(n50653), .B(n36859), .Y(n22520) );
  XNOR2XL U38323 ( .A(n50650), .B(n36860), .Y(n22490) );
  XNOR2XL U38324 ( .A(n50655), .B(n42466), .Y(n21655) );
  XNOR2XL U38325 ( .A(n50652), .B(n36860), .Y(n22510) );
  XNOR2XL U38326 ( .A(n50654), .B(n42465), .Y(n21231) );
  XNOR2XL U38327 ( .A(n50652), .B(n42466), .Y(n21221) );
  XNOR2XL U38328 ( .A(n50651), .B(n42465), .Y(n21211) );
  XNOR2XL U38329 ( .A(n50654), .B(n36854), .Y(n22500) );
  XNOR2XL U38330 ( .A(n50649), .B(n36852), .Y(n22530) );
  XNOR2XL U38331 ( .A(n50657), .B(n42466), .Y(n21675) );
  XNOR2XL U38332 ( .A(n50653), .B(n42462), .Y(n21241) );
  XNOR2XL U38333 ( .A(n50658), .B(n42462), .Y(n21685) );
  XNOR2XL U38334 ( .A(n50655), .B(n36857), .Y(n22621) );
  XNOR2XL U38335 ( .A(n50651), .B(n36853), .Y(n22550) );
  XNOR2XL U38336 ( .A(n50649), .B(n42459), .Y(n21261) );
  XNOR2XL U38337 ( .A(n50648), .B(n36853), .Y(n22480) );
  XNOR2XL U38338 ( .A(n50245), .B(n42671), .Y(n30792) );
  XNOR2XL U38339 ( .A(n50243), .B(n42671), .Y(n30732) );
  XNOR2XL U38340 ( .A(n50244), .B(n41641), .Y(n30740) );
  XNOR2XL U38341 ( .A(n50872), .B(n42613), .Y(n30818) );
  XNOR2XL U38342 ( .A(n50870), .B(n42613), .Y(n30908) );
  XNOR2XL U38343 ( .A(n50873), .B(n42615), .Y(n30848) );
  XNOR2XL U38344 ( .A(n50240), .B(n42671), .Y(n30822) );
  XNOR2XL U38345 ( .A(n50241), .B(n42707), .Y(n30830) );
  XNOR2XL U38346 ( .A(n50238), .B(n42671), .Y(n30912) );
  XNOR2XL U38347 ( .A(n50239), .B(n42712), .Y(n30920) );
  XNOR2XL U38348 ( .A(n50241), .B(n42671), .Y(n30852) );
  XNOR2XL U38349 ( .A(n50242), .B(n42707), .Y(n30860) );
  XNOR2XL U38350 ( .A(n50871), .B(n42613), .Y(n30878) );
  XNOR2XL U38351 ( .A(n50239), .B(n42671), .Y(n30882) );
  XNOR2XL U38352 ( .A(n50240), .B(n42707), .Y(n30890) );
  XNOR2XL U38353 ( .A(n50237), .B(n42710), .Y(n30619) );
  XNOR2XL U38354 ( .A(n50866), .B(n42613), .Y(n30667) );
  XNOR2XL U38355 ( .A(n50227), .B(n42707), .Y(n30257) );
  XNOR2XL U38356 ( .A(n50226), .B(n42673), .Y(n30249) );
  XNOR2XL U38357 ( .A(n50858), .B(n42616), .Y(n30245) );
  XNOR2XL U38358 ( .A(n50228), .B(n42704), .Y(n30227) );
  XNOR2XL U38359 ( .A(n50227), .B(n42673), .Y(n30219) );
  XNOR2XL U38360 ( .A(n50859), .B(n42616), .Y(n30215) );
  XNOR2XL U38361 ( .A(n50236), .B(n41641), .Y(n30649) );
  XNOR2XL U38362 ( .A(n50235), .B(n42671), .Y(n30641) );
  XNOR2XL U38363 ( .A(n50867), .B(n42613), .Y(n30637) );
  XNOR2XL U38364 ( .A(n50235), .B(n42707), .Y(n30679) );
  XNOR2XL U38365 ( .A(n50234), .B(n42671), .Y(n30671) );
  XNOR2XL U38366 ( .A(n50234), .B(n42706), .Y(n30499) );
  XNOR2XL U38367 ( .A(n50233), .B(n42673), .Y(n30491) );
  XNOR2XL U38368 ( .A(n50865), .B(n42616), .Y(n30487) );
  XNOR2XL U38369 ( .A(n50233), .B(n42710), .Y(n30469) );
  XNOR2XL U38370 ( .A(n50232), .B(n42672), .Y(n30461) );
  XNOR2XL U38371 ( .A(n50864), .B(n42615), .Y(n30457) );
  XNOR2XL U38372 ( .A(n50232), .B(n42710), .Y(n30559) );
  XNOR2XL U38373 ( .A(n50231), .B(n42676), .Y(n30551) );
  XNOR2XL U38374 ( .A(n50863), .B(n42616), .Y(n30547) );
  XNOR2XL U38375 ( .A(n50231), .B(n41641), .Y(n30589) );
  XNOR2XL U38376 ( .A(n50230), .B(n42675), .Y(n30581) );
  XNOR2XL U38377 ( .A(n50862), .B(n42616), .Y(n30577) );
  XNOR2XL U38378 ( .A(n50230), .B(n42711), .Y(n30317) );
  XNOR2XL U38379 ( .A(n50229), .B(n42675), .Y(n30309) );
  XNOR2XL U38380 ( .A(n50861), .B(n42616), .Y(n30305) );
  XNOR2XL U38381 ( .A(n50229), .B(n42706), .Y(n30287) );
  XNOR2XL U38382 ( .A(n50228), .B(n42669), .Y(n30279) );
  XNOR2XL U38383 ( .A(n50860), .B(n42616), .Y(n30275) );
  XNOR2XL U38384 ( .A(n50884), .B(n36795), .Y(n21350) );
  XNOR2XL U38385 ( .A(n50882), .B(n36797), .Y(n21330) );
  XNOR2XL U38386 ( .A(n50879), .B(n41295), .Y(n22640) );
  XNOR2XL U38387 ( .A(n50878), .B(n41297), .Y(n22650) );
  XNOR2XL U38388 ( .A(n50881), .B(n36790), .Y(n21320) );
  XNOR2XL U38389 ( .A(n50876), .B(n41296), .Y(n22589) );
  XNOR2XL U38390 ( .A(n50879), .B(n36791), .Y(n21360) );
  XNOR2XL U38391 ( .A(n50875), .B(n41291), .Y(n22579) );
  XNOR2XL U38392 ( .A(n50877), .B(n41296), .Y(n22670) );
  XNOR2XL U38393 ( .A(n50878), .B(n36791), .Y(n21310) );
  XNOR2XL U38394 ( .A(n50880), .B(n36791), .Y(n21370) );
  XNOR2XL U38395 ( .A(n50874), .B(n41292), .Y(n22569) );
  XNOR2XL U38396 ( .A(n50872), .B(n41290), .Y(n22629) );
  XNOR2XL U38397 ( .A(n50877), .B(n36792), .Y(n21300) );
  XNOR2XL U38398 ( .A(n50873), .B(n41292), .Y(n22559) );
  XNOR2XL U38399 ( .A(n50875), .B(n36797), .Y(n21633) );
  XNOR2XL U38400 ( .A(n50874), .B(n36793), .Y(n21623) );
  XNOR2XL U38401 ( .A(n50876), .B(n36799), .Y(n21643) );
  XNOR2XL U38402 ( .A(n50871), .B(n41295), .Y(n22609) );
  XNOR2XL U38403 ( .A(n50873), .B(n36789), .Y(n21613) );
  XNOR2XL U38404 ( .A(n50870), .B(n41297), .Y(n22599) );
  XNOR2XL U38405 ( .A(n50870), .B(n36789), .Y(n21663) );
  XNOR2XL U38406 ( .A(n50867), .B(n41294), .Y(n22518) );
  XNOR2XL U38407 ( .A(n50864), .B(n41293), .Y(n22488) );
  XNOR2XL U38408 ( .A(n50869), .B(n36795), .Y(n21653) );
  XNOR2XL U38409 ( .A(n50866), .B(n41294), .Y(n22508) );
  XNOR2XL U38410 ( .A(n50868), .B(n36798), .Y(n21229) );
  XNOR2XL U38411 ( .A(n50866), .B(n36792), .Y(n21219) );
  XNOR2XL U38412 ( .A(n50865), .B(n36795), .Y(n21209) );
  XNOR2XL U38413 ( .A(n50868), .B(n41293), .Y(n22498) );
  XNOR2XL U38414 ( .A(n50863), .B(n41296), .Y(n22528) );
  XNOR2XL U38415 ( .A(n50871), .B(n36798), .Y(n21673) );
  XNOR2XL U38416 ( .A(n50867), .B(n36799), .Y(n21239) );
  XNOR2XL U38417 ( .A(n50872), .B(n36797), .Y(n21683) );
  XNOR2XL U38418 ( .A(n50869), .B(n41293), .Y(n22619) );
  XNOR2XL U38419 ( .A(n50865), .B(n41297), .Y(n22548) );
  XNOR2XL U38420 ( .A(n50863), .B(n36793), .Y(n21259) );
  XNOR2XL U38421 ( .A(n50862), .B(n41294), .Y(n22478) );
  XNOR2XL U38422 ( .A(n50663), .B(n42592), .Y(n30790) );
  XNOR2XL U38423 ( .A(n51093), .B(n42547), .Y(n32342) );
  XNOR2XL U38424 ( .A(n50661), .B(n42592), .Y(n30730) );
  XNOR2XL U38425 ( .A(n51094), .B(n42548), .Y(n31892) );
  XNOR2XL U38426 ( .A(n51090), .B(n42549), .Y(n30779) );
  XNOR2XL U38427 ( .A(n51092), .B(n42552), .Y(n31952) );
  XNOR2XL U38428 ( .A(n51089), .B(n36832), .Y(n30749) );
  XNOR2XL U38429 ( .A(n51300), .B(n36867), .Y(n30824) );
  XNOR2XL U38430 ( .A(n51087), .B(n36832), .Y(n30689) );
  XNOR2XL U38431 ( .A(n51298), .B(n42642), .Y(n30914) );
  XNOR2XL U38432 ( .A(n50658), .B(n34450), .Y(n30820) );
  XNOR2XL U38433 ( .A(n51301), .B(n42641), .Y(n30854) );
  XNOR2XL U38434 ( .A(n50656), .B(n42592), .Y(n30910) );
  XNOR2XL U38435 ( .A(n51088), .B(n36832), .Y(n30719) );
  XNOR2XL U38436 ( .A(n50659), .B(n42592), .Y(n30850) );
  XNOR2XL U38437 ( .A(n51299), .B(n42643), .Y(n30884) );
  XNOR2XL U38438 ( .A(n50657), .B(n42592), .Y(n30880) );
  XNOR2XL U38439 ( .A(n51296), .B(n42643), .Y(n30613) );
  XNOR2XL U38440 ( .A(n51085), .B(n42553), .Y(n30809) );
  XNOR2XL U38441 ( .A(n51086), .B(n42549), .Y(n30839) );
  XNOR2XL U38442 ( .A(n51083), .B(n36832), .Y(n30899) );
  XNOR2XL U38443 ( .A(n51294), .B(n42643), .Y(n30673) );
  XNOR2XL U38444 ( .A(n51082), .B(n42552), .Y(n30508) );
  XNOR2XL U38445 ( .A(n51286), .B(n42639), .Y(n30251) );
  XNOR2XL U38446 ( .A(n50644), .B(n42589), .Y(n30247) );
  XNOR2XL U38447 ( .A(n51287), .B(n42639), .Y(n30221) );
  XNOR2XL U38448 ( .A(n50645), .B(n36865), .Y(n30217) );
  XNOR2XL U38449 ( .A(n51295), .B(n42639), .Y(n30643) );
  XNOR2XL U38450 ( .A(n50653), .B(n36863), .Y(n30639) );
  XNOR2XL U38451 ( .A(n51084), .B(n36832), .Y(n30869) );
  XNOR2XL U38452 ( .A(n50652), .B(n42592), .Y(n30669) );
  XNOR2XL U38453 ( .A(n51293), .B(n42639), .Y(n30493) );
  XNOR2XL U38454 ( .A(n50651), .B(n36865), .Y(n30489) );
  XNOR2XL U38455 ( .A(n51292), .B(n42639), .Y(n30463) );
  XNOR2XL U38456 ( .A(n50650), .B(n36863), .Y(n30459) );
  XNOR2XL U38457 ( .A(n51080), .B(n36832), .Y(n30628) );
  XNOR2XL U38458 ( .A(n51079), .B(n36832), .Y(n30658) );
  XNOR2XL U38459 ( .A(n51291), .B(n42639), .Y(n30553) );
  XNOR2XL U38460 ( .A(n50649), .B(n42589), .Y(n30549) );
  XNOR2XL U38461 ( .A(n51290), .B(n42639), .Y(n30583) );
  XNOR2XL U38462 ( .A(n50648), .B(n42587), .Y(n30579) );
  XNOR2XL U38463 ( .A(n51289), .B(n42639), .Y(n30311) );
  XNOR2XL U38464 ( .A(n50647), .B(n42592), .Y(n30307) );
  XNOR2XL U38465 ( .A(n51288), .B(n42639), .Y(n30281) );
  XNOR2XL U38466 ( .A(n50646), .B(n36865), .Y(n30277) );
  XNOR2XL U38467 ( .A(n50454), .B(n36905), .Y(n30793) );
  XNOR2XL U38468 ( .A(n36931), .B(n36905), .Y(n30733) );
  XNOR2XL U38469 ( .A(n50665), .B(n42504), .Y(n32343) );
  XNOR2XL U38470 ( .A(n50666), .B(n34458), .Y(n31893) );
  XNOR2XL U38471 ( .A(n37020), .B(n42723), .Y(n30831) );
  XNOR2XL U38472 ( .A(n37245), .B(n42724), .Y(n30921) );
  XNOR2XL U38473 ( .A(n50662), .B(n42505), .Y(n30780) );
  XNOR2XL U38474 ( .A(n37244), .B(n36875), .Y(n30861) );
  XNOR2XL U38475 ( .A(n50664), .B(n36737), .Y(n31953) );
  XNOR2XL U38476 ( .A(n51086), .B(n42624), .Y(n30819) );
  XNOR2XL U38477 ( .A(n50661), .B(n42505), .Y(n30750) );
  XNOR2XL U38478 ( .A(n50659), .B(n42505), .Y(n30690) );
  XNOR2XL U38479 ( .A(n51084), .B(n42627), .Y(n30909) );
  XNOR2XL U38480 ( .A(n36925), .B(n41380), .Y(n30823) );
  XNOR2XL U38481 ( .A(n51087), .B(n42624), .Y(n30849) );
  XNOR2XL U38482 ( .A(n36925), .B(n42724), .Y(n30891) );
  XNOR2XL U38483 ( .A(n36946), .B(n36905), .Y(n30913) );
  XNOR2XL U38484 ( .A(n37020), .B(n36905), .Y(n30853) );
  XNOR2XL U38485 ( .A(n50660), .B(n42505), .Y(n30720) );
  XNOR2XL U38486 ( .A(n51085), .B(n42631), .Y(n30879) );
  XNOR2XL U38487 ( .A(n50452), .B(n42723), .Y(n30620) );
  XNOR2XL U38488 ( .A(n36946), .B(n42719), .Y(n30530) );
  XNOR2XL U38489 ( .A(n37245), .B(n36905), .Y(n30883) );
  XNOR2XL U38490 ( .A(n50657), .B(n42499), .Y(n30810) );
  XNOR2XL U38491 ( .A(n50658), .B(n42505), .Y(n30840) );
  XNOR2XL U38492 ( .A(n50450), .B(n42723), .Y(n30680) );
  XNOR2XL U38493 ( .A(n50655), .B(n42499), .Y(n30900) );
  XNOR2XL U38494 ( .A(n50451), .B(n42723), .Y(n30650) );
  XNOR2XL U38495 ( .A(n51080), .B(n34447), .Y(n30668) );
  XNOR2XL U38496 ( .A(n50448), .B(n42719), .Y(n30470) );
  XNOR2XL U38497 ( .A(n50654), .B(n42503), .Y(n30509) );
  XNOR2XL U38498 ( .A(n50653), .B(n42503), .Y(n30599) );
  XNOR2XL U38499 ( .A(n50650), .B(n42503), .Y(n30479) );
  XNOR2XL U38500 ( .A(n50647), .B(n42503), .Y(n30569) );
  XNOR2XL U38501 ( .A(n50442), .B(n42719), .Y(n30258) );
  XNOR2XL U38502 ( .A(n50441), .B(n36903), .Y(n30250) );
  XNOR2XL U38503 ( .A(n51072), .B(n42632), .Y(n30246) );
  XNOR2XL U38504 ( .A(n50648), .B(n42503), .Y(n30539) );
  XNOR2XL U38505 ( .A(n50443), .B(n42719), .Y(n30228) );
  XNOR2XL U38506 ( .A(n50442), .B(n36903), .Y(n30220) );
  XNOR2XL U38507 ( .A(n51073), .B(n42627), .Y(n30216) );
  XNOR2XL U38508 ( .A(n50450), .B(n36903), .Y(n30642) );
  XNOR2XL U38509 ( .A(n51081), .B(n42633), .Y(n30638) );
  XNOR2XL U38510 ( .A(n50656), .B(n42499), .Y(n30870) );
  XNOR2XL U38511 ( .A(n50449), .B(n41380), .Y(n30672) );
  XNOR2XL U38512 ( .A(n50449), .B(n42719), .Y(n30500) );
  XNOR2XL U38513 ( .A(n50448), .B(n41380), .Y(n30492) );
  XNOR2XL U38514 ( .A(n51079), .B(n42626), .Y(n30488) );
  XNOR2XL U38515 ( .A(n50649), .B(n42503), .Y(n30449) );
  XNOR2XL U38516 ( .A(n50447), .B(n36905), .Y(n30462) );
  XNOR2XL U38517 ( .A(n51078), .B(n42627), .Y(n30458) );
  XNOR2XL U38518 ( .A(n50652), .B(n42503), .Y(n30629) );
  XNOR2XL U38519 ( .A(n50651), .B(n42503), .Y(n30659) );
  XNOR2XL U38520 ( .A(n50438), .B(n42719), .Y(n30378) );
  XNOR2XL U38521 ( .A(n50447), .B(n42719), .Y(n30560) );
  XNOR2XL U38522 ( .A(n50446), .B(n36903), .Y(n30552) );
  XNOR2XL U38523 ( .A(n51077), .B(n42630), .Y(n30548) );
  XNOR2XL U38524 ( .A(n50446), .B(n42719), .Y(n30590) );
  XNOR2XL U38525 ( .A(n50445), .B(n36903), .Y(n30582) );
  XNOR2XL U38526 ( .A(n51076), .B(n42628), .Y(n30578) );
  XNOR2XL U38527 ( .A(n50445), .B(n42719), .Y(n30318) );
  XNOR2XL U38528 ( .A(n50444), .B(n36834), .Y(n30310) );
  XNOR2XL U38529 ( .A(n51075), .B(n42633), .Y(n30306) );
  XNOR2XL U38530 ( .A(n50444), .B(n42719), .Y(n30288) );
  XNOR2XL U38531 ( .A(n50443), .B(n36903), .Y(n30280) );
  XNOR2XL U38532 ( .A(n51074), .B(n34447), .Y(n30276) );
  XNOR2XL U38533 ( .A(n51091), .B(n42549), .Y(n32312) );
  XNOR2XL U38534 ( .A(n50663), .B(n36731), .Y(n32313) );
  XNOR2XL U38535 ( .A(n50873), .B(n40039), .Y(n30826) );
  XNOR2XL U38536 ( .A(n51087), .B(n41281), .Y(n30827) );
  XNOR2XL U38537 ( .A(n50659), .B(net219468), .Y(n30828) );
  XNOR2XL U38538 ( .A(n50871), .B(n40039), .Y(n30916) );
  XNOR2XL U38539 ( .A(n51085), .B(n41283), .Y(n30917) );
  XNOR2XL U38540 ( .A(n50657), .B(net219468), .Y(n30918) );
  XNOR2XL U38541 ( .A(n50874), .B(net258262), .Y(n30856) );
  XNOR2XL U38542 ( .A(n51088), .B(n41281), .Y(n30857) );
  XNOR2XL U38543 ( .A(n50660), .B(net219468), .Y(n30858) );
  XNOR2XL U38544 ( .A(n50869), .B(net219330), .Y(n30615) );
  XNOR2XL U38545 ( .A(n51083), .B(n41282), .Y(n30616) );
  XNOR2XL U38546 ( .A(n50655), .B(net219468), .Y(n30617) );
  XNOR2XL U38547 ( .A(n50870), .B(n36870), .Y(n30525) );
  XNOR2XL U38548 ( .A(n51084), .B(n41282), .Y(n30526) );
  XNOR2XL U38549 ( .A(n50867), .B(n40039), .Y(n30675) );
  XNOR2XL U38550 ( .A(n51081), .B(n41283), .Y(n30676) );
  XNOR2XL U38551 ( .A(n50653), .B(net219468), .Y(n30677) );
  XNOR2XL U38552 ( .A(n50865), .B(n40039), .Y(n30465) );
  XNOR2XL U38553 ( .A(n51079), .B(n41281), .Y(n30466) );
  XNOR2XL U38554 ( .A(n50651), .B(net219434), .Y(n30467) );
  XNOR2XL U38555 ( .A(n50859), .B(n40039), .Y(n30253) );
  XNOR2XL U38556 ( .A(n51073), .B(n41281), .Y(n30254) );
  XNOR2XL U38557 ( .A(n50645), .B(net219434), .Y(n30255) );
  XNOR2XL U38558 ( .A(n50860), .B(net258262), .Y(n30223) );
  XNOR2XL U38559 ( .A(n51074), .B(n41282), .Y(n30224) );
  XNOR2XL U38560 ( .A(n50646), .B(net219434), .Y(n30225) );
  XNOR2XL U38561 ( .A(n50866), .B(net219330), .Y(n30495) );
  XNOR2XL U38562 ( .A(n51080), .B(n41281), .Y(n30496) );
  XNOR2XL U38563 ( .A(n50652), .B(net219434), .Y(n30497) );
  XNOR2XL U38564 ( .A(n50858), .B(n40039), .Y(n30403) );
  XNOR2XL U38565 ( .A(n51072), .B(n41281), .Y(n30404) );
  XNOR2XL U38566 ( .A(n50644), .B(net219434), .Y(n30405) );
  XNOR2XL U38567 ( .A(n50857), .B(net219314), .Y(n30433) );
  XNOR2XL U38568 ( .A(n51071), .B(n41282), .Y(n30434) );
  XNOR2XL U38569 ( .A(n50643), .B(net219434), .Y(n30435) );
  XNOR2XL U38570 ( .A(n50856), .B(net219310), .Y(n30343) );
  XNOR2XL U38571 ( .A(n51070), .B(n41282), .Y(n30344) );
  XNOR2XL U38572 ( .A(n50642), .B(net219434), .Y(n30345) );
  XNOR2XL U38573 ( .A(n50855), .B(net219310), .Y(n30373) );
  XNOR2XL U38574 ( .A(n51069), .B(n41283), .Y(n30374) );
  XNOR2XL U38575 ( .A(n50641), .B(net219434), .Y(n30375) );
  XNOR2XL U38576 ( .A(n50863), .B(net219330), .Y(n30585) );
  XNOR2XL U38577 ( .A(n51077), .B(n41281), .Y(n30586) );
  XNOR2XL U38578 ( .A(n50649), .B(net219468), .Y(n30587) );
  XNOR2XL U38579 ( .A(n50862), .B(n40039), .Y(n30313) );
  XNOR2XL U38580 ( .A(n51076), .B(n41281), .Y(n30314) );
  XNOR2XL U38581 ( .A(n50648), .B(net219434), .Y(n30315) );
  XOR2XL U38582 ( .A(n42232), .B(n36807), .Y(n22664) );
  XOR2XL U38583 ( .A(n42228), .B(n42485), .Y(n21354) );
  XOR2XL U38584 ( .A(n42231), .B(n36808), .Y(n22794) );
  XOR2XL U38585 ( .A(n42230), .B(n42485), .Y(n21334) );
  XOR2XL U38586 ( .A(n42233), .B(n36809), .Y(n22644) );
  XOR2XL U38587 ( .A(n42234), .B(n36814), .Y(n22654) );
  XOR2XL U38588 ( .A(n42231), .B(n42485), .Y(n21324) );
  XOR2XL U38589 ( .A(n42236), .B(n36810), .Y(n22593) );
  XOR2XL U38590 ( .A(n42237), .B(n36817), .Y(n22583) );
  XOR2XL U38591 ( .A(n42235), .B(n36810), .Y(n22674) );
  XOR2XL U38592 ( .A(n42233), .B(n42485), .Y(n21364) );
  XOR2XL U38593 ( .A(n42234), .B(n42485), .Y(n21314) );
  XOR2XL U38594 ( .A(n42232), .B(n42485), .Y(n21374) );
  XOR2XL U38595 ( .A(n42238), .B(n36817), .Y(n22573) );
  XOR2XL U38596 ( .A(n42240), .B(n36816), .Y(n22633) );
  XOR2XL U38597 ( .A(n42235), .B(n42485), .Y(n21304) );
  XOR2XL U38598 ( .A(n42239), .B(n36811), .Y(n22563) );
  XOR2XL U38599 ( .A(n42237), .B(n42483), .Y(n21637) );
  XOR2XL U38600 ( .A(n42238), .B(n42483), .Y(n21627) );
  XOR2XL U38601 ( .A(n42236), .B(n42488), .Y(n21647) );
  XOR2XL U38602 ( .A(n42241), .B(n36815), .Y(n22613) );
  XOR2XL U38603 ( .A(n42239), .B(n42483), .Y(n21617) );
  XOR2XL U38604 ( .A(n42242), .B(n36814), .Y(n22603) );
  XOR2XL U38605 ( .A(n42242), .B(n42492), .Y(n21667) );
  XOR2XL U38606 ( .A(n42245), .B(n36816), .Y(n22522) );
  XOR2XL U38607 ( .A(n42248), .B(n36813), .Y(n22492) );
  XOR2XL U38608 ( .A(n42243), .B(n42483), .Y(n21657) );
  XOR2XL U38609 ( .A(n42246), .B(n36814), .Y(n22512) );
  XOR2XL U38610 ( .A(n42244), .B(n42490), .Y(n21233) );
  XOR2XL U38611 ( .A(n42246), .B(n42490), .Y(n21223) );
  XOR2XL U38612 ( .A(n42247), .B(n42490), .Y(n21213) );
  XOR2XL U38613 ( .A(n42244), .B(n36810), .Y(n22502) );
  XOR2XL U38614 ( .A(n42249), .B(n36813), .Y(n22532) );
  XOR2XL U38615 ( .A(n42241), .B(n42488), .Y(n21677) );
  XOR2XL U38616 ( .A(n42245), .B(n42490), .Y(n21243) );
  XOR2XL U38617 ( .A(n42240), .B(n42487), .Y(n21687) );
  XOR2XL U38618 ( .A(n42243), .B(n36809), .Y(n22623) );
  XOR2XL U38619 ( .A(n42247), .B(n36809), .Y(n22552) );
  XOR2XL U38620 ( .A(n42250), .B(n36810), .Y(n22482) );
  XNOR2XL U38621 ( .A(n50879), .B(n42533), .Y(n32341) );
  XNOR2XL U38622 ( .A(n50880), .B(n42544), .Y(n31891) );
  XNOR2XL U38623 ( .A(n50877), .B(n42535), .Y(n32311) );
  XNOR2XL U38624 ( .A(n50876), .B(n42536), .Y(n30778) );
  XNOR2XL U38625 ( .A(n50878), .B(n42538), .Y(n31951) );
  XNOR2XL U38626 ( .A(n50875), .B(n42536), .Y(n30748) );
  XNOR2XL U38627 ( .A(n50873), .B(n42536), .Y(n30688) );
  XNOR2XL U38628 ( .A(n50874), .B(n42536), .Y(n30718) );
  XNOR2XL U38629 ( .A(n50871), .B(n42536), .Y(n30808) );
  XNOR2XL U38630 ( .A(n50872), .B(n42536), .Y(n30838) );
  XNOR2XL U38631 ( .A(n50869), .B(n42536), .Y(n30898) );
  XNOR2XL U38632 ( .A(n50870), .B(n42536), .Y(n30868) );
  XNOR2XL U38633 ( .A(n50868), .B(n42541), .Y(n30507) );
  XNOR2XL U38634 ( .A(n50865), .B(n42536), .Y(n30657) );
  XNOR2XL U38635 ( .A(n36930), .B(n42579), .Y(n32346) );
  XNOR2XL U38636 ( .A(n51307), .B(n41303), .Y(n22665) );
  XNOR2XL U38637 ( .A(n51308), .B(n41301), .Y(n22795) );
  XNOR2XL U38638 ( .A(n51311), .B(n36740), .Y(n21355) );
  XNOR2XL U38639 ( .A(n51309), .B(n36744), .Y(n21335) );
  XNOR2XL U38640 ( .A(n51306), .B(n41304), .Y(n22645) );
  XNOR2XL U38641 ( .A(n50455), .B(n36776), .Y(n22655) );
  XNOR2XL U38642 ( .A(n51308), .B(n36744), .Y(n21325) );
  XNOR2XL U38643 ( .A(n50453), .B(n36780), .Y(n22594) );
  XNOR2XL U38644 ( .A(n51303), .B(n41300), .Y(n22584) );
  XNOR2XL U38645 ( .A(n50454), .B(n36780), .Y(n22675) );
  XNOR2XL U38646 ( .A(n51306), .B(n36741), .Y(n21365) );
  XNOR2XL U38647 ( .A(n37242), .B(n36743), .Y(n21315) );
  XNOR2XL U38648 ( .A(n51307), .B(n36749), .Y(n21375) );
  XNOR2XL U38649 ( .A(n51300), .B(n41305), .Y(n22634) );
  XNOR2XL U38650 ( .A(n50454), .B(n36770), .Y(n21305) );
  XNOR2XL U38651 ( .A(n51303), .B(n36740), .Y(n21638) );
  XNOR2XL U38652 ( .A(n51302), .B(n36750), .Y(n21628) );
  XNOR2XL U38653 ( .A(n50453), .B(n36766), .Y(n21648) );
  XNOR2XL U38654 ( .A(n51299), .B(n41299), .Y(n22614) );
  XNOR2XL U38655 ( .A(n51301), .B(n36744), .Y(n21618) );
  XNOR2XL U38656 ( .A(n51298), .B(n41305), .Y(n22604) );
  XNOR2XL U38657 ( .A(n51298), .B(n36749), .Y(n21668) );
  XNOR2XL U38658 ( .A(n51297), .B(n36740), .Y(n21658) );
  XNOR2XL U38659 ( .A(n51296), .B(n36748), .Y(n21234) );
  XNOR2XL U38660 ( .A(n50449), .B(n36771), .Y(n21224) );
  XNOR2XL U38661 ( .A(n50448), .B(n36767), .Y(n21214) );
  XNOR2XL U38662 ( .A(n51299), .B(n36742), .Y(n21678) );
  XNOR2XL U38663 ( .A(n50450), .B(n36766), .Y(n21244) );
  XNOR2XL U38664 ( .A(n51300), .B(n36740), .Y(n21688) );
  XNOR2XL U38665 ( .A(n51297), .B(n41303), .Y(n22624) );
  XOR2XL U38666 ( .A(n41974), .B(n36761), .Y(n21363) );
  XNOR2XL U38667 ( .A(n50665), .B(n42461), .Y(n21362) );
  XNOR2XL U38668 ( .A(n51093), .B(n36714), .Y(n21361) );
  XNOR2XL U38669 ( .A(n37019), .B(n42579), .Y(n31896) );
  XNOR2XL U38670 ( .A(n50454), .B(n42577), .Y(n32316) );
  XNOR2XL U38671 ( .A(n50453), .B(n42575), .Y(n30783) );
  XNOR2XL U38672 ( .A(n50455), .B(n42579), .Y(n31956) );
  XNOR2XL U38673 ( .A(n36931), .B(n42579), .Y(n30753) );
  XNOR2XL U38674 ( .A(n37020), .B(n42579), .Y(n30693) );
  XNOR2XL U38675 ( .A(n37244), .B(n42579), .Y(n30723) );
  XNOR2XL U38676 ( .A(n37245), .B(n42581), .Y(n30813) );
  XNOR2XL U38677 ( .A(n36925), .B(n42579), .Y(n30843) );
  XNOR2XL U38678 ( .A(n50452), .B(n42583), .Y(n30903) );
  XNOR2XL U38679 ( .A(n36946), .B(n42583), .Y(n30873) );
  XNOR2XL U38680 ( .A(n50448), .B(n42584), .Y(n30662) );
  XNOR2XL U38681 ( .A(n51302), .B(n41299), .Y(n22574) );
  XNOR2XL U38682 ( .A(n51301), .B(n41300), .Y(n22564) );
  XNOR2XL U38683 ( .A(n51296), .B(n41301), .Y(n22503) );
  XOR2XL U38684 ( .A(n42234), .B(n41321), .Y(n31955) );
  XOR2XL U38685 ( .A(n42237), .B(n36873), .Y(n30752) );
  XOR2XL U38686 ( .A(n42239), .B(n41322), .Y(n30692) );
  XOR2XL U38687 ( .A(n42238), .B(n36801), .Y(n30722) );
  XOR2XL U38688 ( .A(n42240), .B(n36873), .Y(n30842) );
  XOR2XL U38689 ( .A(n42243), .B(n36873), .Y(n30902) );
  XOR2XL U38690 ( .A(n42241), .B(n41321), .Y(n30812) );
  XOR2XL U38691 ( .A(n42242), .B(n36877), .Y(n30872) );
  XOR2XL U38692 ( .A(n42245), .B(n36877), .Y(n30601) );
  XOR2XL U38693 ( .A(n42244), .B(n41322), .Y(n30511) );
  XOR2XL U38694 ( .A(n42248), .B(n36801), .Y(n30481) );
  XOR2XL U38695 ( .A(n42251), .B(n36877), .Y(n30571) );
  XOR2XL U38696 ( .A(n42252), .B(n36877), .Y(n30299) );
  XOR2XL U38697 ( .A(n42250), .B(n36873), .Y(n30541) );
  XOR2XL U38698 ( .A(n42249), .B(n41323), .Y(n30451) );
  XOR2XL U38699 ( .A(n42246), .B(n41323), .Y(n30631) );
  XOR2XL U38700 ( .A(n42247), .B(n36877), .Y(n30661) );
  XOR2XL U38701 ( .A(n42253), .B(n36801), .Y(n30269) );
  OAI211XL U38702 ( .A0(n36898), .A1(n42909), .B0(n13126), .C0(n50068), .Y(
        n34548) );
  OA22XL U38703 ( .A0(net263292), .A1(n42527), .B0(n42609), .B1(n40078), .Y(
        n13126) );
  INVX1 U38704 ( .A(n13128), .Y(n50068) );
  OAI211XL U38705 ( .A0(n42609), .A1(n42910), .B0(n13102), .C0(n50070), .Y(
        n34540) );
  OA22XL U38706 ( .A0(net218416), .A1(n41317), .B0(n42527), .B1(n40078), .Y(
        n13102) );
  INVX1 U38707 ( .A(n13104), .Y(n50070) );
  OAI211XL U38708 ( .A0(n42663), .A1(n42910), .B0(n13090), .C0(n50071), .Y(
        n34536) );
  OA22XL U38709 ( .A0(net218428), .A1(n36808), .B0(n36877), .B1(net218672),
        .Y(n13090) );
  INVX1 U38710 ( .A(n13092), .Y(n50071) );
  OAI211XL U38711 ( .A0(n36886), .A1(n42909), .B0(n13114), .C0(n50069), .Y(
        n34544) );
  OA22XL U38712 ( .A0(net218426), .A1(n41321), .B0(n42663), .B1(n40078), .Y(
        n13114) );
  INVX1 U38713 ( .A(n13116), .Y(n50069) );
  OAI211XL U38714 ( .A0(n42691), .A1(n42909), .B0(n13117), .C0(n13118), .Y(
        n34545) );
  OA22XL U38715 ( .A0(net263045), .A1(n36828), .B0(n42644), .B1(n40078), .Y(
        n13117) );
  OAI211XL U38716 ( .A0(n42707), .A1(n42909), .B0(n13111), .C0(n13112), .Y(
        n34543) );
  OA22XL U38717 ( .A0(net263083), .A1(n42568), .B0(n36907), .B1(n40078), .Y(
        n13111) );
  OAI211XL U38718 ( .A0(n42163), .A1(n42735), .B0(n16786), .C0(n49763), .Y(
        n35768) );
  OA22XL U38719 ( .A0(net218294), .A1(n41888), .B0(n41887), .B1(net218610),
        .Y(n17230) );
  OAI211XL U38720 ( .A0(n41889), .A1(n42846), .B0(n17158), .C0(n49732), .Y(
        n35892) );
  OAI211XL U38721 ( .A0(n41890), .A1(n42847), .B0(n17134), .C0(n49734), .Y(
        n35884) );
  OAI211XL U38722 ( .A0(n41892), .A1(n42752), .B0(n17086), .C0(n49738), .Y(
        n35868) );
  OAI211XL U38723 ( .A0(n41893), .A1(n42753), .B0(n17062), .C0(n49740), .Y(
        n35860) );
  OAI211XL U38724 ( .A0(n42145), .A1(n42843), .B0(n17218), .C0(n49727), .Y(
        n35912) );
  OAI211XL U38725 ( .A0(n42146), .A1(n42844), .B0(n17194), .C0(n49729), .Y(
        n35904) );
  OAI211XL U38726 ( .A0(n42147), .A1(n42845), .B0(n17170), .C0(n49731), .Y(
        n35896) );
  OAI211XL U38727 ( .A0(n42148), .A1(n42846), .B0(n17146), .C0(n49733), .Y(
        n35888) );
  OAI211XL U38728 ( .A0(n42149), .A1(n42750), .B0(n17122), .C0(n49735), .Y(
        n35880) );
  OAI211XL U38729 ( .A0(n42150), .A1(n42751), .B0(n17098), .C0(n49737), .Y(
        n35872) );
  OAI211XL U38730 ( .A0(n42151), .A1(n42753), .B0(n17074), .C0(n49739), .Y(
        n35864) );
  OAI211XL U38731 ( .A0(n42152), .A1(n42754), .B0(n17050), .C0(n49741), .Y(
        n35856) );
  OAI211XL U38732 ( .A0(n41810), .A1(n42816), .B0(n19078), .C0(n49572), .Y(
        n36532) );
  OAI211XL U38733 ( .A0(n41811), .A1(n42816), .B0(n19054), .C0(n49574), .Y(
        n36524) );
  OAI211XL U38734 ( .A0(n41813), .A1(n42817), .B0(n19006), .C0(n49578), .Y(
        n36508) );
  OAI211XL U38735 ( .A0(n34351), .A1(n42817), .B0(n18982), .C0(n49580), .Y(
        n36500) );
  OAI211XL U38736 ( .A0(n41815), .A1(n42818), .B0(n18934), .C0(n49584), .Y(
        n36484) );
  OAI211XL U38737 ( .A0(n41816), .A1(n42818), .B0(n18910), .C0(n49586), .Y(
        n36476) );
  OAI211XL U38738 ( .A0(n41817), .A1(n42818), .B0(n18886), .C0(n49588), .Y(
        n36468) );
  OAI211XL U38739 ( .A0(n41819), .A1(n42819), .B0(n18838), .C0(n49592), .Y(
        n36452) );
  OAI211XL U38740 ( .A0(n41820), .A1(n42819), .B0(n18814), .C0(n49594), .Y(
        n36444) );
  OAI211XL U38741 ( .A0(n41822), .A1(n42820), .B0(n18766), .C0(n49598), .Y(
        n36428) );
  OAI211XL U38742 ( .A0(n41823), .A1(n42820), .B0(n18742), .C0(n49600), .Y(
        n36420) );
  OAI211XL U38743 ( .A0(n41824), .A1(n42820), .B0(n18718), .C0(n49602), .Y(
        n36412) );
  OAI211XL U38744 ( .A0(n41826), .A1(n42821), .B0(n18670), .C0(n49606), .Y(
        n36396) );
  OAI211XL U38745 ( .A0(n41827), .A1(n42821), .B0(n18646), .C0(n49608), .Y(
        n36388) );
  OAI211XL U38746 ( .A0(n41829), .A1(n42822), .B0(n18598), .C0(n49612), .Y(
        n36372) );
  OAI211XL U38747 ( .A0(n41830), .A1(n42822), .B0(n18574), .C0(n49614), .Y(
        n36364) );
  OAI211XL U38748 ( .A0(n41831), .A1(n42822), .B0(n18550), .C0(n49616), .Y(
        n36356) );
  OAI211XL U38749 ( .A0(n41833), .A1(n42823), .B0(n18502), .C0(n49620), .Y(
        n36340) );
  OAI211XL U38750 ( .A0(n41834), .A1(n42823), .B0(n18478), .C0(n49622), .Y(
        n36332) );
  OAI211XL U38751 ( .A0(n41836), .A1(n42824), .B0(n18430), .C0(n49626), .Y(
        n36316) );
  OAI211XL U38752 ( .A0(n41837), .A1(n42824), .B0(n18406), .C0(n49628), .Y(
        n36308) );
  OAI211XL U38753 ( .A0(n41839), .A1(n42825), .B0(n18358), .C0(n49632), .Y(
        n36292) );
  OAI211XL U38754 ( .A0(n41840), .A1(n42825), .B0(n18334), .C0(n49634), .Y(
        n36284) );
  OAI211XL U38755 ( .A0(n41841), .A1(n42825), .B0(n18310), .C0(n49636), .Y(
        n36276) );
  OAI211XL U38756 ( .A0(n41842), .A1(n42826), .B0(n18286), .C0(n49638), .Y(
        n36268) );
  OAI211XL U38757 ( .A0(n41843), .A1(n42826), .B0(n18262), .C0(n49640), .Y(
        n36260) );
  OAI211XL U38758 ( .A0(n41844), .A1(n42826), .B0(n18238), .C0(n49642), .Y(
        n36252) );
  OAI211XL U38759 ( .A0(n41845), .A1(n42827), .B0(n18214), .C0(n49644), .Y(
        n36244) );
  OAI211XL U38760 ( .A0(n41846), .A1(n42828), .B0(n18190), .C0(n49646), .Y(
        n36236) );
  OAI211XL U38761 ( .A0(n41847), .A1(n42829), .B0(n18166), .C0(n49648), .Y(
        n36228) );
  OAI211XL U38762 ( .A0(n41850), .A1(n42801), .B0(n18094), .C0(n49654), .Y(
        n36204) );
  OAI211XL U38763 ( .A0(n41851), .A1(n42802), .B0(n18070), .C0(n49656), .Y(
        n36196) );
  OAI211XL U38764 ( .A0(n41852), .A1(n42803), .B0(n18046), .C0(n49658), .Y(
        n36188) );
  OAI211XL U38765 ( .A0(n41853), .A1(n42804), .B0(n18022), .C0(n49660), .Y(
        n36180) );
  OAI211XL U38766 ( .A0(n41854), .A1(n42805), .B0(n17998), .C0(n49662), .Y(
        n36172) );
  OAI211XL U38767 ( .A0(n41856), .A1(n42808), .B0(n17950), .C0(n49666), .Y(
        n36156) );
  OAI211XL U38768 ( .A0(n41858), .A1(n42810), .B0(n17902), .C0(n49670), .Y(
        n36140) );
  OAI211XL U38769 ( .A0(n41859), .A1(n42811), .B0(n17878), .C0(n49672), .Y(
        n36132) );
  OAI211XL U38770 ( .A0(n41861), .A1(n42813), .B0(n17830), .C0(n49676), .Y(
        n36116) );
  OAI211XL U38771 ( .A0(n41867), .A1(n42852), .B0(n17686), .C0(n49688), .Y(
        n36068) );
  OAI211XL U38772 ( .A0(n41868), .A1(n42854), .B0(n17662), .C0(n49690), .Y(
        n36060) );
  OAI211XL U38773 ( .A0(n41870), .A1(n42856), .B0(n17614), .C0(n49694), .Y(
        n36044) );
  OAI211XL U38774 ( .A0(n41871), .A1(n42857), .B0(n17590), .C0(n49696), .Y(
        n36036) );
  OAI211XL U38775 ( .A0(n41872), .A1(n42858), .B0(n17566), .C0(n49698), .Y(
        n36028) );
  OAI211XL U38776 ( .A0(n41873), .A1(n42859), .B0(n17542), .C0(n49700), .Y(
        n36020) );
  OAI211XL U38777 ( .A0(n41874), .A1(n42861), .B0(n17518), .C0(n49702), .Y(
        n36012) );
  OAI211XL U38778 ( .A0(n41876), .A1(n42863), .B0(n17470), .C0(n49706), .Y(
        n35996) );
  OA22XL U38779 ( .A0(net218294), .A1(n41887), .B0(n41886), .B1(net218610),
        .Y(n17254) );
  OAI211XL U38780 ( .A0(n41901), .A1(n42762), .B0(n16870), .C0(n49756), .Y(
        n35796) );
  OAI211XL U38781 ( .A0(n41902), .A1(n42764), .B0(n16846), .C0(n49758), .Y(
        n35788) );
  OAI211XL U38782 ( .A0(n41903), .A1(n42765), .B0(n16822), .C0(n49760), .Y(
        n35780) );
  OAI211XL U38783 ( .A0(n41914), .A1(n42745), .B0(n16558), .C0(n49782), .Y(
        n35692) );
  OAI211XL U38784 ( .A0(n41915), .A1(n42746), .B0(n16534), .C0(n49784), .Y(
        n35684) );
  OAI211XL U38785 ( .A0(n41916), .A1(n42748), .B0(n16510), .C0(n49786), .Y(
        n35676) );
  OAI211XL U38786 ( .A0(n41917), .A1(n42749), .B0(n16486), .C0(n49788), .Y(
        n35668) );
  OAI211XL U38787 ( .A0(n41918), .A1(n42750), .B0(n16462), .C0(n49790), .Y(
        n35660) );
  OAI211XL U38788 ( .A0(n41919), .A1(n42783), .B0(n16438), .C0(n49792), .Y(
        n35652) );
  OAI211XL U38789 ( .A0(n41920), .A1(n42784), .B0(n16414), .C0(n49794), .Y(
        n35644) );
  OAI211XL U38790 ( .A0(n41924), .A1(n42789), .B0(n16318), .C0(n49802), .Y(
        n35612) );
  OAI211XL U38791 ( .A0(n41925), .A1(n42790), .B0(n16294), .C0(n49804), .Y(
        n35604) );
  OAI211XL U38792 ( .A0(n41926), .A1(n42791), .B0(n16270), .C0(n49806), .Y(
        n35596) );
  OAI211XL U38793 ( .A0(n41927), .A1(n42792), .B0(n16246), .C0(n49808), .Y(
        n35588) );
  OAI211XL U38794 ( .A0(n41928), .A1(n42794), .B0(n16222), .C0(n49810), .Y(
        n35580) );
  OAI211XL U38795 ( .A0(n41929), .A1(n42795), .B0(n16198), .C0(n49812), .Y(
        n35572) );
  OAI211XL U38796 ( .A0(n41930), .A1(n42796), .B0(n16174), .C0(n49814), .Y(
        n35564) );
  OAI211XL U38797 ( .A0(n41931), .A1(n42797), .B0(n16150), .C0(n49816), .Y(
        n35556) );
  OAI211XL U38798 ( .A0(n41932), .A1(n42798), .B0(n16126), .C0(n49818), .Y(
        n35548) );
  OAI211XL U38799 ( .A0(n41933), .A1(n42767), .B0(n16102), .C0(n49820), .Y(
        n35540) );
  OAI211XL U38800 ( .A0(n41935), .A1(n42769), .B0(n16054), .C0(n49824), .Y(
        n35524) );
  OAI211XL U38801 ( .A0(n41936), .A1(n42770), .B0(n16030), .C0(n49826), .Y(
        n35516) );
  OAI211XL U38802 ( .A0(n41937), .A1(n42772), .B0(n16006), .C0(n49828), .Y(
        n35508) );
  OAI211XL U38803 ( .A0(n41938), .A1(n42773), .B0(n15982), .C0(n49830), .Y(
        n35500) );
  OAI211XL U38804 ( .A0(n41939), .A1(n42774), .B0(n15958), .C0(n49832), .Y(
        n35492) );
  OAI211XL U38805 ( .A0(n41940), .A1(n42775), .B0(n15934), .C0(n49834), .Y(
        n35484) );
  OAI211XL U38806 ( .A0(n41941), .A1(n42776), .B0(n15910), .C0(n49836), .Y(
        n35476) );
  OAI211XL U38807 ( .A0(n41943), .A1(n42779), .B0(n15862), .C0(n49840), .Y(
        n35460) );
  OAI211XL U38808 ( .A0(n41944), .A1(n42780), .B0(n15838), .C0(n49842), .Y(
        n35452) );
  OAI211XL U38809 ( .A0(n41946), .A1(n42782), .B0(n15790), .C0(n49846), .Y(
        n35436) );
  OAI211XL U38810 ( .A0(n41947), .A1(n42944), .B0(n15766), .C0(n49848), .Y(
        n35428) );
  OAI211XL U38811 ( .A0(n41948), .A1(n42945), .B0(n15742), .C0(n49850), .Y(
        n35420) );
  OAI211XL U38812 ( .A0(n41949), .A1(n42946), .B0(n15718), .C0(n49852), .Y(
        n35412) );
  OAI211XL U38813 ( .A0(n41950), .A1(n42947), .B0(n15694), .C0(n49854), .Y(
        n35404) );
  OAI211XL U38814 ( .A0(n41951), .A1(n42948), .B0(n15670), .C0(n49856), .Y(
        n35396) );
  OAI211XL U38815 ( .A0(n41952), .A1(n42950), .B0(n15646), .C0(n49858), .Y(
        n35388) );
  OAI211XL U38816 ( .A0(n41953), .A1(n42951), .B0(n15622), .C0(n49860), .Y(
        n35380) );
  OAI211XL U38817 ( .A0(n41955), .A1(n42953), .B0(n15574), .C0(n49864), .Y(
        n35364) );
  OAI211XL U38818 ( .A0(n41956), .A1(n42954), .B0(n15550), .C0(n49866), .Y(
        n35356) );
  OAI211XL U38819 ( .A0(n41957), .A1(n42955), .B0(n15526), .C0(n49868), .Y(
        n35348) );
  OAI211XL U38820 ( .A0(n41958), .A1(n42957), .B0(n15502), .C0(n49870), .Y(
        n35340) );
  INVX1 U38821 ( .A(n15480), .Y(n49872) );
  INVX1 U38822 ( .A(n15456), .Y(n49874) );
  INVX1 U38823 ( .A(n15432), .Y(n49876) );
  INVX1 U38824 ( .A(n15408), .Y(n49878) );
  INVX1 U38825 ( .A(n15384), .Y(n49880) );
  INVX1 U38826 ( .A(n15360), .Y(n49882) );
  INVX1 U38827 ( .A(n15336), .Y(n49884) );
  INVX1 U38828 ( .A(n15312), .Y(n49886) );
  INVX1 U38829 ( .A(n15288), .Y(n49888) );
  INVX1 U38830 ( .A(n15264), .Y(n49890) );
  INVX1 U38831 ( .A(n15240), .Y(n49892) );
  INVX1 U38832 ( .A(n15216), .Y(n49894) );
  INVX1 U38833 ( .A(n15192), .Y(n49896) );
  INVX1 U38834 ( .A(n15168), .Y(n49898) );
  INVX1 U38835 ( .A(n14520), .Y(n49952) );
  INVX1 U38836 ( .A(n14496), .Y(n49954) );
  INVX1 U38837 ( .A(n14472), .Y(n49956) );
  INVX1 U38838 ( .A(n14448), .Y(n49958) );
  INVX1 U38839 ( .A(n14424), .Y(n49960) );
  INVX1 U38840 ( .A(n14376), .Y(n49964) );
  INVX1 U38841 ( .A(n14352), .Y(n49966) );
  INVX1 U38842 ( .A(n14328), .Y(n49968) );
  INVX1 U38843 ( .A(n14304), .Y(n49970) );
  INVX1 U38844 ( .A(n14280), .Y(n49972) );
  INVX1 U38845 ( .A(n14256), .Y(n49974) );
  INVX1 U38846 ( .A(n14232), .Y(n49976) );
  INVX1 U38847 ( .A(n14208), .Y(n49978) );
  INVX1 U38848 ( .A(n14184), .Y(n49980) );
  INVX1 U38849 ( .A(n14160), .Y(n49982) );
  INVX1 U38850 ( .A(n14136), .Y(n49984) );
  INVX1 U38851 ( .A(n14112), .Y(n49986) );
  INVX1 U38852 ( .A(n14088), .Y(n49988) );
  INVX1 U38853 ( .A(n14016), .Y(n49994) );
  INVX1 U38854 ( .A(n13728), .Y(n50018) );
  INVX1 U38855 ( .A(n13704), .Y(n50020) );
  INVX1 U38856 ( .A(n13680), .Y(n50022) );
  INVX1 U38857 ( .A(n13656), .Y(n50024) );
  INVX1 U38858 ( .A(n13632), .Y(n50026) );
  INVX1 U38859 ( .A(n13608), .Y(n50028) );
  INVX1 U38860 ( .A(n13584), .Y(n50030) );
  INVX1 U38861 ( .A(n13560), .Y(n50032) );
  INVX1 U38862 ( .A(n13536), .Y(n50034) );
  INVX1 U38863 ( .A(n13512), .Y(n50036) );
  INVX1 U38864 ( .A(n13488), .Y(n50038) );
  INVX1 U38865 ( .A(n13464), .Y(n50040) );
  INVX1 U38866 ( .A(n13440), .Y(n50042) );
  INVX1 U38867 ( .A(n13416), .Y(n50044) );
  INVX1 U38868 ( .A(n13392), .Y(n50046) );
  INVX1 U38869 ( .A(n13368), .Y(n50048) );
  INVX1 U38870 ( .A(n13344), .Y(n50050) );
  INVX1 U38871 ( .A(n13320), .Y(n50052) );
  INVX1 U38872 ( .A(n13296), .Y(n50054) );
  INVX1 U38873 ( .A(n13272), .Y(n50056) );
  INVX1 U38874 ( .A(n13248), .Y(n50058) );
  INVX1 U38875 ( .A(n13224), .Y(n50060) );
  INVX1 U38876 ( .A(n13200), .Y(n50062) );
  INVX1 U38877 ( .A(n13176), .Y(n50064) );
  OA22XL U38878 ( .A0(net263292), .A1(n42609), .B0(n36895), .B1(n40079), .Y(
        n13150) );
  INVX1 U38879 ( .A(n13152), .Y(n50066) );
  OAI211XL U38880 ( .A0(n42527), .A1(n42910), .B0(n13076), .C0(n50072), .Y(
        n34532) );
  OA22XL U38881 ( .A0(net218418), .A1(n36753), .B0(n41318), .B1(net218650),
        .Y(n13076) );
  INVX1 U38882 ( .A(n13078), .Y(n50072) );
  OAI211XL U38883 ( .A0(n42067), .A1(n42816), .B0(n19090), .C0(n49571), .Y(
        n36536) );
  OAI211XL U38884 ( .A0(n42068), .A1(n42816), .B0(n19066), .C0(n49573), .Y(
        n36528) );
  OAI211XL U38885 ( .A0(n42069), .A1(n42817), .B0(n19042), .C0(n49575), .Y(
        n36520) );
  OAI211XL U38886 ( .A0(n42070), .A1(n42817), .B0(n19018), .C0(n49577), .Y(
        n36512) );
  OAI211XL U38887 ( .A0(n42071), .A1(n42817), .B0(n18994), .C0(n49579), .Y(
        n36504) );
  OAI211XL U38888 ( .A0(n42072), .A1(n42817), .B0(n18970), .C0(n49581), .Y(
        n36496) );
  OAI211XL U38889 ( .A0(n42073), .A1(n42818), .B0(n18946), .C0(n49583), .Y(
        n36488) );
  OAI211XL U38890 ( .A0(n42074), .A1(n42818), .B0(n18922), .C0(n49585), .Y(
        n36480) );
  OAI211XL U38891 ( .A0(n42075), .A1(n42818), .B0(n18898), .C0(n49587), .Y(
        n36472) );
  OAI211XL U38892 ( .A0(n42076), .A1(n42819), .B0(n18874), .C0(n49589), .Y(
        n36464) );
  OAI211XL U38893 ( .A0(n42077), .A1(n42819), .B0(n18850), .C0(n49591), .Y(
        n36456) );
  OAI211XL U38894 ( .A0(n42078), .A1(n42819), .B0(n18826), .C0(n49593), .Y(
        n36448) );
  OAI211XL U38895 ( .A0(n42079), .A1(n42819), .B0(n18802), .C0(n49595), .Y(
        n36440) );
  OAI211XL U38896 ( .A0(n42080), .A1(n42820), .B0(n18778), .C0(n49597), .Y(
        n36432) );
  OAI211XL U38897 ( .A0(n42081), .A1(n42820), .B0(n18754), .C0(n49599), .Y(
        n36424) );
  OAI211XL U38898 ( .A0(n42082), .A1(n42820), .B0(n18730), .C0(n49601), .Y(
        n36416) );
  OAI211XL U38899 ( .A0(n42083), .A1(n42821), .B0(n18706), .C0(n49603), .Y(
        n36408) );
  OAI211XL U38900 ( .A0(n42084), .A1(n42821), .B0(n18682), .C0(n49605), .Y(
        n36400) );
  OAI211XL U38901 ( .A0(n42085), .A1(n42821), .B0(n18658), .C0(n49607), .Y(
        n36392) );
  OAI211XL U38902 ( .A0(n42086), .A1(n42821), .B0(n18634), .C0(n49609), .Y(
        n36384) );
  OAI211XL U38903 ( .A0(n42087), .A1(n42822), .B0(n18610), .C0(n49611), .Y(
        n36376) );
  OAI211XL U38904 ( .A0(n42088), .A1(n42822), .B0(n18586), .C0(n49613), .Y(
        n36368) );
  OAI211XL U38905 ( .A0(n42089), .A1(n42822), .B0(n18562), .C0(n49615), .Y(
        n36360) );
  OAI211XL U38906 ( .A0(n42090), .A1(n42823), .B0(n18538), .C0(n49617), .Y(
        n36352) );
  OAI211XL U38907 ( .A0(n42091), .A1(n42823), .B0(n18514), .C0(n49619), .Y(
        n36344) );
  OAI211XL U38908 ( .A0(n42092), .A1(n42823), .B0(n18490), .C0(n49621), .Y(
        n36336) );
  OAI211XL U38909 ( .A0(n42093), .A1(n42824), .B0(n18466), .C0(n49623), .Y(
        n36328) );
  OAI211XL U38910 ( .A0(n42094), .A1(n42824), .B0(n18442), .C0(n49625), .Y(
        n36320) );
  OAI211XL U38911 ( .A0(n42095), .A1(n42824), .B0(n18418), .C0(n49627), .Y(
        n36312) );
  OAI211XL U38912 ( .A0(n42096), .A1(n42824), .B0(n18394), .C0(n49629), .Y(
        n36304) );
  OAI211XL U38913 ( .A0(n42097), .A1(n42825), .B0(n18370), .C0(n49631), .Y(
        n36296) );
  OAI211XL U38914 ( .A0(n42098), .A1(n42825), .B0(n18346), .C0(n49633), .Y(
        n36288) );
  OAI211XL U38915 ( .A0(n42099), .A1(n42825), .B0(n18322), .C0(n49635), .Y(
        n36280) );
  OAI211XL U38916 ( .A0(n42100), .A1(n42826), .B0(n18298), .C0(n49637), .Y(
        n36272) );
  OAI211XL U38917 ( .A0(n42101), .A1(n42826), .B0(n18274), .C0(n49639), .Y(
        n36264) );
  OAI211XL U38918 ( .A0(n42102), .A1(n42826), .B0(n18250), .C0(n49641), .Y(
        n36256) );
  OAI211XL U38919 ( .A0(n42103), .A1(n42827), .B0(n18226), .C0(n49643), .Y(
        n36248) );
  OAI211XL U38920 ( .A0(n42104), .A1(n42828), .B0(n18202), .C0(n49645), .Y(
        n36240) );
  OAI211XL U38921 ( .A0(n42105), .A1(n42829), .B0(n18178), .C0(n49647), .Y(
        n36232) );
  OAI211XL U38922 ( .A0(n42108), .A1(n42800), .B0(n18106), .C0(n49653), .Y(
        n36208) );
  OAI211XL U38923 ( .A0(n42109), .A1(n42801), .B0(n18082), .C0(n49655), .Y(
        n36200) );
  OAI211XL U38924 ( .A0(n42110), .A1(n42802), .B0(n18058), .C0(n49657), .Y(
        n36192) );
  OAI211XL U38925 ( .A0(n42111), .A1(n42804), .B0(n18034), .C0(n49659), .Y(
        n36184) );
  OAI211XL U38926 ( .A0(n42112), .A1(n42805), .B0(n18010), .C0(n49661), .Y(
        n36176) );
  OAI211XL U38927 ( .A0(n42113), .A1(n42806), .B0(n17986), .C0(n49663), .Y(
        n36168) );
  OAI211XL U38928 ( .A0(n42115), .A1(n42808), .B0(n17938), .C0(n49667), .Y(
        n36152) );
  OAI211XL U38929 ( .A0(n42116), .A1(n42809), .B0(n17914), .C0(n49669), .Y(
        n36144) );
  OAI211XL U38930 ( .A0(n42117), .A1(n42811), .B0(n17890), .C0(n49671), .Y(
        n36136) );
  OAI211XL U38931 ( .A0(n42118), .A1(n42812), .B0(n17866), .C0(n49673), .Y(
        n36128) );
  OAI211XL U38932 ( .A0(n42119), .A1(n42813), .B0(n17842), .C0(n49675), .Y(
        n36120) );
  OAI211XL U38933 ( .A0(n42120), .A1(n42814), .B0(n17818), .C0(n49677), .Y(
        n36112) );
  OAI211XL U38934 ( .A0(n42121), .A1(n42847), .B0(n17794), .C0(n49679), .Y(
        n36104) );
  OAI211XL U38935 ( .A0(n42122), .A1(n42848), .B0(n17770), .C0(n49681), .Y(
        n36096) );
  OAI211XL U38936 ( .A0(n42123), .A1(n42850), .B0(n17746), .C0(n49683), .Y(
        n36088) );
  OAI211XL U38937 ( .A0(n42124), .A1(n42851), .B0(n17722), .C0(n49685), .Y(
        n36080) );
  OAI211XL U38938 ( .A0(n42125), .A1(n42852), .B0(n17698), .C0(n49687), .Y(
        n36072) );
  OAI211XL U38939 ( .A0(n42126), .A1(n42853), .B0(n17674), .C0(n49689), .Y(
        n36064) );
  OAI211XL U38940 ( .A0(n42127), .A1(n42854), .B0(n17650), .C0(n49691), .Y(
        n36056) );
  OAI211XL U38941 ( .A0(n42128), .A1(n42855), .B0(n17626), .C0(n49693), .Y(
        n36048) );
  OAI211XL U38942 ( .A0(n42129), .A1(n42857), .B0(n17602), .C0(n49695), .Y(
        n36040) );
  OAI211XL U38943 ( .A0(n42130), .A1(n42858), .B0(n17578), .C0(n49697), .Y(
        n36032) );
  OAI211XL U38944 ( .A0(n42131), .A1(n42859), .B0(n17554), .C0(n49699), .Y(
        n36024) );
  OAI211XL U38945 ( .A0(n42132), .A1(n42860), .B0(n17530), .C0(n49701), .Y(
        n36016) );
  OAI211XL U38946 ( .A0(n42133), .A1(n42861), .B0(n17506), .C0(n49703), .Y(
        n36008) );
  OAI211XL U38947 ( .A0(n42134), .A1(n42862), .B0(n17482), .C0(n49705), .Y(
        n36000) );
  OAI211XL U38948 ( .A0(n42135), .A1(n42831), .B0(n17458), .C0(n49707), .Y(
        n35992) );
  OAI211XL U38949 ( .A0(n42136), .A1(n42832), .B0(n17434), .C0(n49709), .Y(
        n35984) );
  OAI211XL U38950 ( .A0(n42137), .A1(n42833), .B0(n17410), .C0(n49711), .Y(
        n35976) );
  OAI211XL U38951 ( .A0(n42138), .A1(n42835), .B0(n17386), .C0(n49713), .Y(
        n35968) );
  OAI211XL U38952 ( .A0(n42139), .A1(n42836), .B0(n17362), .C0(n49715), .Y(
        n35960) );
  OAI211XL U38953 ( .A0(n42140), .A1(n42837), .B0(n17338), .C0(n49717), .Y(
        n35952) );
  OAI211XL U38954 ( .A0(n42142), .A1(n42839), .B0(n17290), .C0(n49721), .Y(
        n35936) );
  OAI211XL U38955 ( .A0(n42143), .A1(n42840), .B0(n17266), .C0(n49723), .Y(
        n35928) );
  OAI211XL U38956 ( .A0(n42144), .A1(n42842), .B0(n17242), .C0(n49725), .Y(
        n35920) );
  OA22XL U38957 ( .A0(net218294), .A1(n42146), .B0(n42145), .B1(net218610),
        .Y(n17242) );
  OAI211XL U38958 ( .A0(n42159), .A1(n42762), .B0(n16882), .C0(n49755), .Y(
        n35800) );
  OAI211XL U38959 ( .A0(n42160), .A1(n42763), .B0(n16858), .C0(n49757), .Y(
        n35792) );
  OAI211XL U38960 ( .A0(n42161), .A1(n42764), .B0(n16834), .C0(n49759), .Y(
        n35784) );
  OAI211XL U38961 ( .A0(n42162), .A1(n42765), .B0(n16810), .C0(n49761), .Y(
        n35776) );
  OAI211XL U38962 ( .A0(n42169), .A1(n42741), .B0(n16642), .C0(n49775), .Y(
        n35720) );
  OAI211XL U38963 ( .A0(n42170), .A1(n42742), .B0(n16618), .C0(n49777), .Y(
        n35712) );
  OAI211XL U38964 ( .A0(n42171), .A1(n42744), .B0(n16594), .C0(n49779), .Y(
        n35704) );
  OAI211XL U38965 ( .A0(n42172), .A1(n42745), .B0(n16570), .C0(n49781), .Y(
        n35696) );
  OAI211XL U38966 ( .A0(n42173), .A1(n42746), .B0(n16546), .C0(n49783), .Y(
        n35688) );
  OAI211XL U38967 ( .A0(n42174), .A1(n42747), .B0(n16522), .C0(n49785), .Y(
        n35680) );
  OAI211XL U38968 ( .A0(n42175), .A1(n42748), .B0(n16498), .C0(n49787), .Y(
        n35672) );
  OAI211XL U38969 ( .A0(n42176), .A1(n42749), .B0(n16474), .C0(n49789), .Y(
        n35664) );
  OAI211XL U38970 ( .A0(n42177), .A1(n42783), .B0(n16450), .C0(n49791), .Y(
        n35656) );
  OAI211XL U38971 ( .A0(n42178), .A1(n42784), .B0(n16426), .C0(n49793), .Y(
        n35648) );
  OAI211XL U38972 ( .A0(n42179), .A1(n42785), .B0(n16402), .C0(n49795), .Y(
        n35640) );
  OAI211XL U38973 ( .A0(n42181), .A1(n42787), .B0(n16354), .C0(n49799), .Y(
        n35624) );
  OAI211XL U38974 ( .A0(n42182), .A1(n42788), .B0(n16330), .C0(n49801), .Y(
        n35616) );
  OAI211XL U38975 ( .A0(n42183), .A1(n42789), .B0(n16306), .C0(n49803), .Y(
        n35608) );
  OAI211XL U38976 ( .A0(n42184), .A1(n42791), .B0(n16282), .C0(n49805), .Y(
        n35600) );
  OAI211XL U38977 ( .A0(n42185), .A1(n42792), .B0(n16258), .C0(n49807), .Y(
        n35592) );
  OAI211XL U38978 ( .A0(n42186), .A1(n42793), .B0(n16234), .C0(n49809), .Y(
        n35584) );
  OAI211XL U38979 ( .A0(n42187), .A1(n42794), .B0(n16210), .C0(n49811), .Y(
        n35576) );
  OAI211XL U38980 ( .A0(n42188), .A1(n42795), .B0(n16186), .C0(n49813), .Y(
        n35568) );
  OAI211XL U38981 ( .A0(n42189), .A1(n42796), .B0(n16162), .C0(n49815), .Y(
        n35560) );
  OAI211XL U38982 ( .A0(n42190), .A1(n42798), .B0(n16138), .C0(n49817), .Y(
        n35552) );
  OAI211XL U38983 ( .A0(n42191), .A1(n42766), .B0(n16114), .C0(n49819), .Y(
        n35544) );
  OAI211XL U38984 ( .A0(n42192), .A1(n42768), .B0(n16090), .C0(n49821), .Y(
        n35536) );
  OAI211XL U38985 ( .A0(n42193), .A1(n42769), .B0(n16066), .C0(n49823), .Y(
        n35528) );
  OAI211XL U38986 ( .A0(n42194), .A1(n42770), .B0(n16042), .C0(n49825), .Y(
        n35520) );
  OAI211XL U38987 ( .A0(n42195), .A1(n42771), .B0(n16018), .C0(n49827), .Y(
        n35512) );
  OAI211XL U38988 ( .A0(n42196), .A1(n42772), .B0(n15994), .C0(n49829), .Y(
        n35504) );
  OAI211XL U38989 ( .A0(n42197), .A1(n42773), .B0(n15970), .C0(n49831), .Y(
        n35496) );
  OAI211XL U38990 ( .A0(n42198), .A1(n42775), .B0(n15946), .C0(n49833), .Y(
        n35488) );
  OAI211XL U38991 ( .A0(n42199), .A1(n42776), .B0(n15922), .C0(n49835), .Y(
        n35480) );
  OAI211XL U38992 ( .A0(n42200), .A1(n42777), .B0(n15898), .C0(n49837), .Y(
        n35472) );
  OAI211XL U38993 ( .A0(n42202), .A1(n42779), .B0(n15850), .C0(n49841), .Y(
        n35456) );
  OAI211XL U38994 ( .A0(n42203), .A1(n42780), .B0(n15826), .C0(n49843), .Y(
        n35448) );
  OAI211XL U38995 ( .A0(n42204), .A1(n42781), .B0(n15802), .C0(n49845), .Y(
        n35440) );
  OAI211XL U38996 ( .A0(n42205), .A1(n42799), .B0(n15778), .C0(n49847), .Y(
        n35432) );
  OAI211XL U38997 ( .A0(n42206), .A1(n42944), .B0(n15754), .C0(n49849), .Y(
        n35424) );
  OAI211XL U38998 ( .A0(n42207), .A1(n42946), .B0(n15730), .C0(n49851), .Y(
        n35416) );
  OAI211XL U38999 ( .A0(n42208), .A1(n42947), .B0(n15706), .C0(n49853), .Y(
        n35408) );
  OAI211XL U39000 ( .A0(n42209), .A1(n42948), .B0(n15682), .C0(n49855), .Y(
        n35400) );
  OAI211XL U39001 ( .A0(n42211), .A1(n42950), .B0(n15634), .C0(n49859), .Y(
        n35384) );
  OAI211XL U39002 ( .A0(n42212), .A1(n42951), .B0(n15610), .C0(n49861), .Y(
        n35376) );
  OAI211XL U39003 ( .A0(n42213), .A1(n42953), .B0(n15586), .C0(n49863), .Y(
        n35368) );
  OAI211XL U39004 ( .A0(n42214), .A1(n42954), .B0(n15562), .C0(n49865), .Y(
        n35360) );
  OAI211XL U39005 ( .A0(n42215), .A1(n42955), .B0(n15538), .C0(n49867), .Y(
        n35352) );
  OAI211XL U39006 ( .A0(n42216), .A1(n42956), .B0(n15514), .C0(n49869), .Y(
        n35344) );
  OAI211XL U39007 ( .A0(n42217), .A1(n42957), .B0(n15490), .C0(n49871), .Y(
        n35336) );
  INVX1 U39008 ( .A(n15468), .Y(n49873) );
  INVX1 U39009 ( .A(n15444), .Y(n49875) );
  INVX1 U39010 ( .A(n15420), .Y(n49877) );
  INVX1 U39011 ( .A(n15396), .Y(n49879) );
  INVX1 U39012 ( .A(n15372), .Y(n49881) );
  INVX1 U39013 ( .A(n15348), .Y(n49883) );
  INVX1 U39014 ( .A(n15324), .Y(n49885) );
  INVX1 U39015 ( .A(n15300), .Y(n49887) );
  INVX1 U39016 ( .A(n15276), .Y(n49889) );
  INVX1 U39017 ( .A(n15252), .Y(n49891) );
  INVX1 U39018 ( .A(n15228), .Y(n49893) );
  INVX1 U39019 ( .A(n15204), .Y(n49895) );
  INVX1 U39020 ( .A(n14532), .Y(n49951) );
  INVX1 U39021 ( .A(n14508), .Y(n49953) );
  INVX1 U39022 ( .A(n14484), .Y(n49955) );
  INVX1 U39023 ( .A(n14460), .Y(n49957) );
  INVX1 U39024 ( .A(n14436), .Y(n49959) );
  INVX1 U39025 ( .A(n14388), .Y(n49963) );
  INVX1 U39026 ( .A(n14364), .Y(n49965) );
  INVX1 U39027 ( .A(n14340), .Y(n49967) );
  INVX1 U39028 ( .A(n14316), .Y(n49969) );
  INVX1 U39029 ( .A(n14292), .Y(n49971) );
  INVX1 U39030 ( .A(n14268), .Y(n49973) );
  INVX1 U39031 ( .A(n14244), .Y(n49975) );
  INVX1 U39032 ( .A(n14220), .Y(n49977) );
  INVX1 U39033 ( .A(n14196), .Y(n49979) );
  INVX1 U39034 ( .A(n14172), .Y(n49981) );
  INVX1 U39035 ( .A(n14148), .Y(n49983) );
  INVX1 U39036 ( .A(n14124), .Y(n49985) );
  INVX1 U39037 ( .A(n14100), .Y(n49987) );
  INVX1 U39038 ( .A(n14076), .Y(n49989) );
  INVX1 U39039 ( .A(n14028), .Y(n49993) );
  INVX1 U39040 ( .A(n13740), .Y(n50017) );
  INVX1 U39041 ( .A(n13716), .Y(n50019) );
  INVX1 U39042 ( .A(n13692), .Y(n50021) );
  INVX1 U39043 ( .A(n13668), .Y(n50023) );
  INVX1 U39044 ( .A(n13644), .Y(n50025) );
  INVX1 U39045 ( .A(n13620), .Y(n50027) );
  INVX1 U39046 ( .A(n13596), .Y(n50029) );
  INVX1 U39047 ( .A(n13572), .Y(n50031) );
  INVX1 U39048 ( .A(n13548), .Y(n50033) );
  INVX1 U39049 ( .A(n13524), .Y(n50035) );
  INVX1 U39050 ( .A(n13500), .Y(n50037) );
  INVX1 U39051 ( .A(n13476), .Y(n50039) );
  INVX1 U39052 ( .A(n13452), .Y(n50041) );
  INVX1 U39053 ( .A(n13428), .Y(n50043) );
  INVX1 U39054 ( .A(n13404), .Y(n50045) );
  INVX1 U39055 ( .A(n13380), .Y(n50047) );
  INVX1 U39056 ( .A(n13356), .Y(n50049) );
  INVX1 U39057 ( .A(n13332), .Y(n50051) );
  INVX1 U39058 ( .A(n13308), .Y(n50053) );
  INVX1 U39059 ( .A(n13284), .Y(n50055) );
  INVX1 U39060 ( .A(n13260), .Y(n50057) );
  INVX1 U39061 ( .A(n13236), .Y(n50059) );
  INVX1 U39062 ( .A(n13212), .Y(n50061) );
  INVX1 U39063 ( .A(n13188), .Y(n50063) );
  INVX1 U39064 ( .A(n13164), .Y(n50065) );
  OA22XL U39065 ( .A0(net263292), .A1(n42663), .B0(n36882), .B1(n40078), .Y(
        n13138) );
  INVX1 U39066 ( .A(n13140), .Y(n50067) );
  OAI211XL U39067 ( .A0(n36877), .A1(n42910), .B0(n13060), .C0(n50073), .Y(
        n34528) );
  OA22XL U39068 ( .A0(net263330), .A1(n42496), .B0(n36809), .B1(net218918),
        .Y(n13060) );
  INVX1 U39069 ( .A(n13062), .Y(n50073) );
  INVX1 U39070 ( .A(n15144), .Y(n49900) );
  INVX1 U39071 ( .A(n15120), .Y(n49902) );
  INVX1 U39072 ( .A(n15096), .Y(n49904) );
  INVX1 U39073 ( .A(n15072), .Y(n49906) );
  INVX1 U39074 ( .A(n15048), .Y(n49908) );
  INVX1 U39075 ( .A(n15024), .Y(n49910) );
  INVX1 U39076 ( .A(n15000), .Y(n49912) );
  INVX1 U39077 ( .A(n14976), .Y(n49914) );
  INVX1 U39078 ( .A(n14952), .Y(n49916) );
  INVX1 U39079 ( .A(n14928), .Y(n49918) );
  INVX1 U39080 ( .A(n14904), .Y(n49920) );
  INVX1 U39081 ( .A(n14880), .Y(n49922) );
  INVX1 U39082 ( .A(n14856), .Y(n49924) );
  INVX1 U39083 ( .A(n14832), .Y(n49926) );
  INVX1 U39084 ( .A(n14808), .Y(n49928) );
  INVX1 U39085 ( .A(n14760), .Y(n49932) );
  INVX1 U39086 ( .A(n14736), .Y(n49934) );
  INVX1 U39087 ( .A(n14712), .Y(n49936) );
  INVX1 U39088 ( .A(n14688), .Y(n49938) );
  INVX1 U39089 ( .A(n14664), .Y(n49940) );
  INVX1 U39090 ( .A(n14640), .Y(n49942) );
  INVX1 U39091 ( .A(n14616), .Y(n49944) );
  INVX1 U39092 ( .A(n14592), .Y(n49946) );
  INVX1 U39093 ( .A(n14568), .Y(n49948) );
  INVX1 U39094 ( .A(n15180), .Y(n49897) );
  INVX1 U39095 ( .A(n15156), .Y(n49899) );
  INVX1 U39096 ( .A(n15132), .Y(n49901) );
  INVX1 U39097 ( .A(n15108), .Y(n49903) );
  INVX1 U39098 ( .A(n15084), .Y(n49905) );
  INVX1 U39099 ( .A(n15060), .Y(n49907) );
  INVX1 U39100 ( .A(n15036), .Y(n49909) );
  INVX1 U39101 ( .A(n15012), .Y(n49911) );
  INVX1 U39102 ( .A(n14988), .Y(n49913) );
  INVX1 U39103 ( .A(n14964), .Y(n49915) );
  INVX1 U39104 ( .A(n14940), .Y(n49917) );
  INVX1 U39105 ( .A(n14916), .Y(n49919) );
  INVX1 U39106 ( .A(n14892), .Y(n49921) );
  INVX1 U39107 ( .A(n14868), .Y(n49923) );
  INVX1 U39108 ( .A(n14844), .Y(n49925) );
  INVX1 U39109 ( .A(n14820), .Y(n49927) );
  INVX1 U39110 ( .A(n14796), .Y(n49929) );
  INVX1 U39111 ( .A(n14748), .Y(n49933) );
  INVX1 U39112 ( .A(n14724), .Y(n49935) );
  INVX1 U39113 ( .A(n14700), .Y(n49937) );
  INVX1 U39114 ( .A(n14676), .Y(n49939) );
  INVX1 U39115 ( .A(n14652), .Y(n49941) );
  INVX1 U39116 ( .A(n14628), .Y(n49943) );
  INVX1 U39117 ( .A(n14604), .Y(n49945) );
  INVX1 U39118 ( .A(n14580), .Y(n49947) );
  OAI211XL U39119 ( .A0(n41281), .A1(n42909), .B0(n13120), .C0(n13121), .Y(
        n34546) );
  OA22XL U39120 ( .A0(net218422), .A1(n42554), .B0(n42631), .B1(n40078), .Y(
        n13120) );
  OAI211XL U39121 ( .A0(net219310), .A1(n42909), .B0(n13123), .C0(n13124), .Y(
        n34547) );
  OA22XL U39122 ( .A0(net261981), .A1(n42544), .B0(n42620), .B1(n40078), .Y(
        n13123) );
  OAI211XL U39123 ( .A0(n41895), .A1(n42755), .B0(n17014), .C0(n49744), .Y(
        n35844) );
  OAI211XL U39124 ( .A0(net219434), .A1(n42909), .B0(n13129), .C0(n13130), .Y(
        n34549) );
  OA22XL U39125 ( .A0(net263292), .A1(n42508), .B0(n42592), .B1(n40078), .Y(
        n13129) );
  OAI211XL U39126 ( .A0(n42725), .A1(n42910), .B0(n13108), .C0(n13109), .Y(
        n34542) );
  OA22XL U39127 ( .A0(net218412), .A1(n42584), .B0(n41380), .B1(n40078), .Y(
        n13108) );
  OAI211XL U39128 ( .A0(n42153), .A1(n42755), .B0(n17026), .C0(n49743), .Y(
        n35848) );
  OAI211XL U39129 ( .A0(n42155), .A1(n42757), .B0(n16978), .C0(n49747), .Y(
        n35832) );
  OAI211XL U39130 ( .A0(n42156), .A1(n42758), .B0(n16954), .C0(n49749), .Y(
        n35824) );
  OAI211XL U39131 ( .A0(n42157), .A1(n42760), .B0(n16930), .C0(n49751), .Y(
        n35816) );
  OAI211XL U39132 ( .A0(n42158), .A1(n42761), .B0(n16906), .C0(n49753), .Y(
        n35808) );
  OAI211XL U39133 ( .A0(n41908), .A1(n42738), .B0(n16702), .C0(n49770), .Y(
        n35740) );
  OAI211XL U39134 ( .A0(n41909), .A1(n42739), .B0(n16678), .C0(n49772), .Y(
        n35732) );
  INVX1 U39135 ( .A(n14400), .Y(n49962) );
  INVX1 U39136 ( .A(n13992), .Y(n49996) );
  INVX1 U39137 ( .A(n13968), .Y(n49998) );
  INVX1 U39138 ( .A(n13944), .Y(n50000) );
  INVX1 U39139 ( .A(n13920), .Y(n50002) );
  INVX1 U39140 ( .A(n13896), .Y(n50004) );
  INVX1 U39141 ( .A(n13872), .Y(n50006) );
  INVX1 U39142 ( .A(n13848), .Y(n50008) );
  INVX1 U39143 ( .A(n13824), .Y(n50010) );
  INVX1 U39144 ( .A(n13800), .Y(n50012) );
  INVX1 U39145 ( .A(n13776), .Y(n50014) );
  INVX1 U39146 ( .A(n13752), .Y(n50016) );
  OAI211XL U39147 ( .A0(n42164), .A1(n42736), .B0(n16762), .C0(n49765), .Y(
        n35760) );
  OAI211XL U39148 ( .A0(n42166), .A1(n42738), .B0(n16714), .C0(n49769), .Y(
        n35744) );
  OAI211XL U39149 ( .A0(n42167), .A1(n42739), .B0(n16690), .C0(n49771), .Y(
        n35736) );
  INVX1 U39150 ( .A(n14412), .Y(n49961) );
  INVX1 U39151 ( .A(n14004), .Y(n49995) );
  INVX1 U39152 ( .A(n13980), .Y(n49997) );
  INVX1 U39153 ( .A(n13956), .Y(n49999) );
  INVX1 U39154 ( .A(n13932), .Y(n50001) );
  INVX1 U39155 ( .A(n13908), .Y(n50003) );
  INVX1 U39156 ( .A(n13884), .Y(n50005) );
  INVX1 U39157 ( .A(n13860), .Y(n50007) );
  INVX1 U39158 ( .A(n13836), .Y(n50009) );
  INVX1 U39159 ( .A(n13812), .Y(n50011) );
  INVX1 U39160 ( .A(n13788), .Y(n50013) );
  INVX1 U39161 ( .A(n13764), .Y(n50015) );
  OAI211XL U39162 ( .A0(n41906), .A1(n42737), .B0(n16750), .C0(n49766), .Y(
        n35756) );
  OAI211XL U39163 ( .A0(n41907), .A1(n42864), .B0(n16726), .C0(n49768), .Y(
        n35748) );
  INVX1 U39164 ( .A(n14064), .Y(n49990) );
  INVX1 U39165 ( .A(n14040), .Y(n49992) );
  OAI211XL U39166 ( .A0(n42165), .A1(n42864), .B0(n16738), .C0(n49767), .Y(
        n35752) );
  INVX1 U39167 ( .A(n14052), .Y(n49991) );
  INVX1 U39168 ( .A(n14784), .Y(n49930) );
  INVX1 U39169 ( .A(n14772), .Y(n49931) );
  INVXL U39170 ( .A(n12274), .Y(net151473) );
  INVXL U39171 ( .A(n10827), .Y(net171453) );
  INVXL U39172 ( .A(n12255), .Y(net151491) );
  INVXL U39173 ( .A(net209778), .Y(net171122) );
  INVXL U39174 ( .A(n10543), .Y(net171304) );
  NAND2BXL U39175 ( .AN(n36830), .B(n42992), .Y(n48713) );
  NAND2BXL U39176 ( .AN(net217206), .B(n41388), .Y(n48714) );
  NAND2XL U39177 ( .A(n10754), .B(n10757), .Y(n11333) );
  NAND2XL U39178 ( .A(n42992), .B(n42570), .Y(n49489) );
  AOI2BB2XL U39179 ( .B0(n50165), .B1(net264960), .A0N(net217178), .A1N(n36907), .Y(n49488) );
  OA22XL U39180 ( .A0(net263330), .A1(n36734), .B0(n36846), .B1(n40140), .Y(
        n13056) );
  NAND2XL U39181 ( .A(n43000), .B(n42677), .Y(n49486) );
  AOI2BB2XL U39182 ( .B0(n50166), .B1(net265207), .A0N(net217178), .A1N(n42707), .Y(n49485) );
  OA22XL U39183 ( .A0(net263083), .A1(n36844), .B0(n42569), .B1(n40050), .Y(
        n13087) );
  NAND2XL U39184 ( .A(n42998), .B(n41251), .Y(n48710) );
  AOI2BB2XL U39185 ( .B0(n51226), .B1(net221720), .A0N(n40281), .A1N(n42701),
        .Y(n48709) );
  OA22XL U39186 ( .A0(net262988), .A1(n41301), .B0(n36829), .B1(n40126), .Y(
        n13093) );
  NAND2XL U39187 ( .A(n42995), .B(n36805), .Y(n48869) );
  AOI2BB2XL U39188 ( .B0(n51012), .B1(net265036), .A0N(n40283), .A1N(n41282),
        .Y(n48868) );
  OA22XL U39189 ( .A0(net263083), .A1(n41329), .B0(n42554), .B1(n40058), .Y(
        n13096) );
  NAND4XL U39190 ( .A(n13068), .B(n48873), .C(n48872), .D(n48871), .Y(n34530)
         );
  NAND2XL U39191 ( .A(n42995), .B(n42555), .Y(n48872) );
  AOI2BB2XL U39192 ( .B0(n51011), .B1(net264960), .A0N(n40283), .A1N(n42629),
        .Y(n48871) );
  OA22XL U39193 ( .A0(net218464), .A1(n36721), .B0(n41328), .B1(net218674),
        .Y(n13068) );
  NAND2XL U39194 ( .A(n42992), .B(n42621), .Y(n49021) );
  AOI2BB2XL U39195 ( .B0(n50798), .B1(net265036), .A0N(n40285), .A1N(net219314), .Y(n49020) );
  OA22XL U39196 ( .A0(net263178), .A1(n41293), .B0(n42544), .B1(n40056), .Y(
        n13099) );
  NAND4XL U39197 ( .A(n13072), .B(net208565), .C(n49024), .D(n49023), .Y(
        n34531) );
  NAND2XL U39198 ( .A(n42996), .B(n42545), .Y(n49024) );
  AOI2BB2XL U39199 ( .B0(n50797), .B1(net264960), .A0N(n40282), .A1N(n42620),
        .Y(n49023) );
  OA22XL U39200 ( .A0(net261924), .A1(n36793), .B0(n41291), .B1(net218832),
        .Y(n13072) );
  NAND2XL U39201 ( .A(n43006), .B(n42593), .Y(n49176) );
  AOI2BB2XL U39202 ( .B0(n50584), .B1(net265207), .A0N(n40287), .A1N(net219468), .Y(n49175) );
  OA22XL U39203 ( .A0(net263178), .A1(n36859), .B0(n42508), .B1(n40078), .Y(
        n13105) );
  NAND2XL U39204 ( .A(n43006), .B(n42509), .Y(n49179) );
  AOI2BB2XL U39205 ( .B0(n50583), .B1(net264960), .A0N(n40289), .A1N(n42592),
        .Y(n49178) );
  OA22XL U39206 ( .A0(net262988), .A1(n42473), .B0(n36856), .B1(n40059), .Y(
        n13079) );
  NAND2XL U39207 ( .A(n43003), .B(n42685), .Y(n49331) );
  AOI2BB2XL U39208 ( .B0(n50381), .B1(net264960), .A0N(n40279), .A1N(n42725),
        .Y(n49330) );
  OA22XL U39209 ( .A0(net263045), .A1(n36783), .B0(n42584), .B1(n40054), .Y(
        n13084) );
  NAND2XL U39210 ( .A(n43003), .B(n42585), .Y(n49334) );
  AOI2BB2XL U39211 ( .B0(n50380), .B1(net221734), .A0N(n40279), .A1N(n36903),
        .Y(n49333) );
  OA22XL U39212 ( .A0(net263330), .A1(n36770), .B0(n36782), .B1(n40060), .Y(
        n13052) );
  INVXL U39213 ( .A(n12906), .Y(net151467) );
  NAND2XL U39214 ( .A(n11360), .B(n10689), .Y(n11357) );
  NAND2XL U39215 ( .A(n50380), .B(n40266), .Y(n49332) );
  NAND2XL U39216 ( .A(net217938), .B(n49442), .Y(n49441) );
  NAND2XL U39217 ( .A(n40221), .B(n49446), .Y(n49445) );
  NAND2XL U39218 ( .A(n40187), .B(n49458), .Y(n49457) );
  NAND2XL U39219 ( .A(net217932), .B(n48750), .Y(n48749) );
  NAND2XL U39220 ( .A(net217960), .B(n48754), .Y(n48753) );
  NAND2XL U39221 ( .A(net217956), .B(n48758), .Y(n48757) );
  NAND2XL U39222 ( .A(net217962), .B(n48762), .Y(n48761) );
  NAND2XL U39223 ( .A(net217938), .B(n48766), .Y(n48765) );
  NAND2XL U39224 ( .A(net217942), .B(n48770), .Y(n48769) );
  NAND2XL U39225 ( .A(net217944), .B(n48774), .Y(n48773) );
  NAND2XL U39226 ( .A(net217964), .B(n48778), .Y(n48777) );
  NAND2XL U39227 ( .A(net217952), .B(n48782), .Y(n48781) );
  NAND2XL U39228 ( .A(net217952), .B(n48786), .Y(n48785) );
  NAND2XL U39229 ( .A(net217936), .B(n49010), .Y(n49009) );
  NAND2XL U39230 ( .A(n40234), .B(n49450), .Y(n49449) );
  NAND2XL U39231 ( .A(n40222), .B(n49454), .Y(n49453) );
  NAND2XL U39232 ( .A(n40234), .B(n49462), .Y(n49461) );
  NAND2XL U39233 ( .A(n40234), .B(n49466), .Y(n49465) );
  NAND2XL U39234 ( .A(n40234), .B(n49470), .Y(n49469) );
  NAND2XL U39235 ( .A(n40244), .B(n49474), .Y(n49473) );
  NAND2XL U39236 ( .A(n40246), .B(n49478), .Y(n49477) );
  NAND2XL U39237 ( .A(n40272), .B(n48568), .Y(n48567) );
  NAND2XL U39238 ( .A(n40272), .B(n41387), .Y(n48571) );
  NAND2XL U39239 ( .A(n40272), .B(n48575), .Y(n48574) );
  NAND2XL U39240 ( .A(n40272), .B(n48579), .Y(n48578) );
  NAND2XL U39241 ( .A(n40272), .B(n48583), .Y(n48582) );
  NAND2XL U39242 ( .A(n40272), .B(n41270), .Y(n48586) );
  NAND2XL U39243 ( .A(n40272), .B(n48590), .Y(n48589) );
  NAND2XL U39244 ( .A(n40272), .B(n48594), .Y(n48593) );
  NAND2XL U39245 ( .A(n40272), .B(n48561), .Y(n48560) );
  INVXL U39246 ( .A(n10233), .Y(net171467) );
  OR2XL U39247 ( .A(n9872), .B(n9982), .Y(n48555) );
  INVXL U39248 ( .A(n12798), .Y(net171201) );
  INVXL U39249 ( .A(n48099), .Y(n12907) );
  AND2XL U39250 ( .A(n12270), .B(n12389), .Y(n11042) );
  AND2XL U39251 ( .A(n12156), .B(n12157), .Y(n12008) );
  AND2XL U39252 ( .A(n12153), .B(n12154), .Y(n12027) );
  NAND4XL U39253 ( .A(n10273), .B(n10272), .C(n10274), .D(n10810), .Y(n22635)
         );
  INVXL U39254 ( .A(net210528), .Y(net212664) );
  NOR3XL U39255 ( .A(n10798), .B(net171480), .C(net151532), .Y(n22473) );
  INVXL U39256 ( .A(n11334), .Y(net151443) );
  NAND3BXL U39257 ( .AN(n10877), .B(n10875), .C(n10879), .Y(n9978) );
  INVXL U39258 ( .A(n11024), .Y(net171460) );
  NAND4XL U39259 ( .A(n37345), .B(n10724), .C(n20096), .D(n10727), .Y(n9919)
         );
  NOR2XL U39260 ( .A(net151726), .B(net151728), .Y(n20096) );
  NAND4XL U39261 ( .A(n10657), .B(n10658), .C(n10659), .D(n21204), .Y(n9881)
         );
  NAND4XL U39262 ( .A(n10734), .B(n10733), .C(n10732), .D(n20178), .Y(n9918)
         );
  NOR2BXL U39263 ( .AN(n10730), .B(n10729), .Y(n20178) );
  NAND4XL U39264 ( .A(n10232), .B(n10233), .C(n10237), .D(n22878), .Y(n9858)
         );
  NOR3XL U39265 ( .A(n10239), .B(n10230), .C(n10231), .Y(n22878) );
  NAND4XL U39266 ( .A(n40390), .B(n10820), .C(n11034), .D(n22796), .Y(n9857)
         );
  NAND4XL U39267 ( .A(n10710), .B(n10709), .C(n10708), .D(n19649), .Y(n9911)
         );
  NAND2XL U39268 ( .A(n12876), .B(n12872), .Y(n10669) );
  XNOR2XL U39269 ( .A(n50836), .B(net219324), .Y(n29531) );
  XNOR2XL U39270 ( .A(n51050), .B(n41281), .Y(n29532) );
  XNOR2XL U39271 ( .A(n50622), .B(net219450), .Y(n29533) );
  NAND4XL U39272 ( .A(n10719), .B(n10715), .C(n12960), .D(n13015), .Y(n9914)
         );
  NAND4XL U39273 ( .A(n11082), .B(n11084), .C(n11085), .D(n11083), .Y(n10247)
         );
  NAND4BXL U39274 ( .AN(n47578), .B(net210512), .C(net210848), .D(n37018), .Y(
        n47841) );
  NAND3XL U39275 ( .A(net210517), .B(n10045), .C(n10044), .Y(n47578) );
  INVXL U39276 ( .A(n10040), .Y(net210848) );
  XOR2XL U39277 ( .A(n41992), .B(n41310), .Y(n22541) );
  XOR2XL U39278 ( .A(n41992), .B(n36753), .Y(n21252) );
  XOR2XL U39279 ( .A(n41989), .B(n36753), .Y(n21272) );
  XOR2XL U39280 ( .A(n41990), .B(n36761), .Y(n21262) );
  XOR2XL U39281 ( .A(n41991), .B(n36761), .Y(n21282) );
  XNOR2XL U39282 ( .A(n51271), .B(n36871), .Y(n29808) );
  XNOR2XL U39283 ( .A(n51263), .B(n42697), .Y(n29507) );
  XNOR2XL U39284 ( .A(n51262), .B(n36871), .Y(n29627) );
  XNOR2XL U39285 ( .A(n51274), .B(n42697), .Y(n29778) );
  XNOR2XL U39286 ( .A(n51273), .B(n42697), .Y(n29748) );
  XNOR2XL U39287 ( .A(n51266), .B(n36871), .Y(n29597) );
  XNOR2XL U39288 ( .A(n51265), .B(n42697), .Y(n29567) );
  XNOR2XL U39289 ( .A(n51264), .B(n36871), .Y(n29537) );
  XNOR2XL U39290 ( .A(n51261), .B(n36871), .Y(n29657) );
  XNOR2XL U39291 ( .A(n51259), .B(n42697), .Y(n29717) );
  NAND4X1 U39292 ( .A(n10755), .B(n10756), .C(n10757), .D(n21689), .Y(n9884)
         );
  NAND4XL U39293 ( .A(n10855), .B(n10854), .C(n10853), .D(n24010), .Y(n10249)
         );
  XOR2XL U39294 ( .A(n42018), .B(n36893), .Y(n29504) );
  XOR2XL U39295 ( .A(n42277), .B(n36881), .Y(n29508) );
  XOR2XL U39296 ( .A(n42278), .B(n42653), .Y(n29500) );
  XOR2XL U39297 ( .A(n42019), .B(n42602), .Y(n29496) );
  XOR2XL U39298 ( .A(n42279), .B(n42653), .Y(n29620) );
  XOR2XL U39299 ( .A(n42020), .B(n42602), .Y(n29616) );
  XOR2XL U39300 ( .A(n42275), .B(n42653), .Y(n29590) );
  XOR2XL U39301 ( .A(n42016), .B(n42602), .Y(n29586) );
  XOR2XL U39302 ( .A(n42016), .B(n36898), .Y(n29564) );
  XOR2XL U39303 ( .A(n42275), .B(n36889), .Y(n29568) );
  XOR2XL U39304 ( .A(n42276), .B(n42653), .Y(n29560) );
  XOR2XL U39305 ( .A(n42017), .B(n42602), .Y(n29556) );
  XOR2XL U39306 ( .A(n42017), .B(n36897), .Y(n29534) );
  XOR2XL U39307 ( .A(n42276), .B(n36880), .Y(n29538) );
  NAND4X1 U39308 ( .A(n39345), .B(n11299), .C(n11519), .D(n21608), .Y(n9880)
         );
  XNOR2XL U39309 ( .A(n50443), .B(n36765), .Y(n22073) );
  XNOR2XL U39310 ( .A(n50444), .B(n36778), .Y(n22543) );
  XOR2XL U39311 ( .A(n41999), .B(n42516), .Y(n30328) );
  XOR2XL U39312 ( .A(n41997), .B(n42516), .Y(n30388) );
  XOR2XL U39313 ( .A(n41998), .B(n42516), .Y(n30418) );
  XOR2XL U39314 ( .A(n42000), .B(n42516), .Y(n30358) );
  XNOR2XL U39315 ( .A(n51075), .B(n41327), .Y(n22539) );
  XNOR2XL U39316 ( .A(n51075), .B(n36716), .Y(n21250) );
  XNOR2XL U39317 ( .A(n51078), .B(n36721), .Y(n21270) );
  XNOR2XL U39318 ( .A(n51076), .B(n36720), .Y(n21280) );
  XNOR2XL U39319 ( .A(n50647), .B(n36860), .Y(n22540) );
  XNOR2XL U39320 ( .A(n50647), .B(n42465), .Y(n21251) );
  XNOR2XL U39321 ( .A(n50650), .B(n42465), .Y(n21271) );
  XNOR2XL U39322 ( .A(n50648), .B(n42465), .Y(n21281) );
  XNOR2XL U39323 ( .A(n50842), .B(n42615), .Y(n29794) );
  XNOR2XL U39324 ( .A(n50834), .B(n42615), .Y(n29493) );
  XNOR2XL U39325 ( .A(n50202), .B(n42711), .Y(n29625) );
  XNOR2XL U39326 ( .A(n50201), .B(n42671), .Y(n29617) );
  XNOR2XL U39327 ( .A(n50833), .B(n42615), .Y(n29613) );
  XNOR2XL U39328 ( .A(n50226), .B(n42705), .Y(n30407) );
  XNOR2XL U39329 ( .A(n50225), .B(n42674), .Y(n30399) );
  XNOR2XL U39330 ( .A(n50857), .B(n42616), .Y(n30395) );
  XNOR2XL U39331 ( .A(n50225), .B(n42710), .Y(n30437) );
  XNOR2XL U39332 ( .A(n50224), .B(n42673), .Y(n30429) );
  XNOR2XL U39333 ( .A(n50856), .B(n42616), .Y(n30425) );
  XNOR2XL U39334 ( .A(n50224), .B(n42711), .Y(n30347) );
  XNOR2XL U39335 ( .A(n50223), .B(n42672), .Y(n30339) );
  XNOR2XL U39336 ( .A(n50855), .B(n42616), .Y(n30335) );
  XNOR2XL U39337 ( .A(n50223), .B(n42711), .Y(n30377) );
  XNOR2XL U39338 ( .A(n50222), .B(n42673), .Y(n30369) );
  XNOR2XL U39339 ( .A(n50854), .B(n42616), .Y(n30365) );
  XNOR2XL U39340 ( .A(n50844), .B(n42615), .Y(n29734) );
  XNOR2XL U39341 ( .A(n50861), .B(n41292), .Y(n22538) );
  XNOR2XL U39342 ( .A(n50861), .B(n36798), .Y(n21249) );
  XNOR2XL U39343 ( .A(n50864), .B(n36789), .Y(n21269) );
  XNOR2XL U39344 ( .A(n50862), .B(n36799), .Y(n21279) );
  XNOR2XL U39345 ( .A(n51270), .B(n42638), .Y(n29800) );
  XNOR2XL U39346 ( .A(n51262), .B(n42639), .Y(n29499) );
  XNOR2XL U39347 ( .A(n51261), .B(n42638), .Y(n29619) );
  XNOR2XL U39348 ( .A(n50619), .B(n42586), .Y(n29615) );
  XNOR2XL U39349 ( .A(n51285), .B(n42639), .Y(n30401) );
  XNOR2XL U39350 ( .A(n50643), .B(n42586), .Y(n30397) );
  XNOR2XL U39351 ( .A(n51284), .B(n42639), .Y(n30431) );
  XNOR2XL U39352 ( .A(n50642), .B(n36863), .Y(n30427) );
  XNOR2XL U39353 ( .A(n51283), .B(n42639), .Y(n30341) );
  XNOR2XL U39354 ( .A(n50641), .B(n42587), .Y(n30337) );
  XNOR2XL U39355 ( .A(n51282), .B(n42639), .Y(n30371) );
  XNOR2XL U39356 ( .A(n50640), .B(n42592), .Y(n30367) );
  XNOR2XL U39357 ( .A(n51272), .B(n42638), .Y(n29740) );
  XNOR2XL U39358 ( .A(n50426), .B(n42717), .Y(n29807) );
  XNOR2XL U39359 ( .A(n51056), .B(n42624), .Y(n29795) );
  XNOR2XL U39360 ( .A(n50418), .B(n42724), .Y(n29506) );
  XNOR2XL U39361 ( .A(n51048), .B(n42626), .Y(n29494) );
  XNOR2XL U39362 ( .A(n50417), .B(n42724), .Y(n29626) );
  XNOR2XL U39363 ( .A(n50416), .B(n36728), .Y(n29618) );
  XNOR2XL U39364 ( .A(n51047), .B(n42625), .Y(n29614) );
  XNOR2XL U39365 ( .A(n50441), .B(n42719), .Y(n30408) );
  XNOR2XL U39366 ( .A(n50440), .B(n41380), .Y(n30400) );
  XNOR2XL U39367 ( .A(n51071), .B(n42630), .Y(n30396) );
  XNOR2XL U39368 ( .A(n50440), .B(n42719), .Y(n30438) );
  XNOR2XL U39369 ( .A(n50439), .B(n36903), .Y(n30430) );
  XNOR2XL U39370 ( .A(n51070), .B(n42633), .Y(n30426) );
  XNOR2XL U39371 ( .A(n50439), .B(n42719), .Y(n30348) );
  XNOR2XL U39372 ( .A(n50438), .B(n36905), .Y(n30340) );
  XNOR2XL U39373 ( .A(n51069), .B(n42627), .Y(n30336) );
  XNOR2XL U39374 ( .A(n50437), .B(n36903), .Y(n30370) );
  XNOR2XL U39375 ( .A(n51068), .B(n42625), .Y(n30366) );
  XNOR2XL U39376 ( .A(n50429), .B(n36875), .Y(n29777) );
  XNOR2XL U39377 ( .A(n50428), .B(n42717), .Y(n29747) );
  XNOR2XL U39378 ( .A(n51058), .B(n42633), .Y(n29735) );
  XNOR2XL U39379 ( .A(n50421), .B(n42717), .Y(n29596) );
  XNOR2XL U39380 ( .A(n50420), .B(n42717), .Y(n29566) );
  XNOR2XL U39381 ( .A(n50640), .B(n42503), .Y(n30327) );
  XNOR2XL U39382 ( .A(n50642), .B(n42503), .Y(n30387) );
  XNOR2XL U39383 ( .A(n50641), .B(n42503), .Y(n30417) );
  XNOR2XL U39384 ( .A(n50639), .B(n42503), .Y(n30357) );
  XNOR2XL U39385 ( .A(n50414), .B(n42717), .Y(n29716) );
  XNOR2XL U39386 ( .A(n51065), .B(n41281), .Y(n30193) );
  XNOR2XL U39387 ( .A(n50637), .B(net219434), .Y(n30194) );
  XNOR2XL U39388 ( .A(n50843), .B(n40039), .Y(n29802) );
  XNOR2XL U39389 ( .A(n50835), .B(n36870), .Y(n29501) );
  XNOR2XL U39390 ( .A(n51049), .B(n41281), .Y(n29502) );
  XNOR2XL U39391 ( .A(n50621), .B(net219442), .Y(n29503) );
  XNOR2XL U39392 ( .A(n50834), .B(net219336), .Y(n29621) );
  XNOR2XL U39393 ( .A(n51048), .B(n41283), .Y(n29622) );
  XNOR2XL U39394 ( .A(n50620), .B(net219450), .Y(n29623) );
  XNOR2XL U39395 ( .A(n50846), .B(net219310), .Y(n29772) );
  XNOR2XL U39396 ( .A(n51060), .B(n41281), .Y(n29773) );
  XNOR2XL U39397 ( .A(n50632), .B(net219450), .Y(n29774) );
  XNOR2XL U39398 ( .A(n50845), .B(net219336), .Y(n29742) );
  XNOR2XL U39399 ( .A(n51059), .B(n41281), .Y(n29743) );
  XNOR2XL U39400 ( .A(n50631), .B(net219450), .Y(n29744) );
  XNOR2XL U39401 ( .A(n50838), .B(n36870), .Y(n29591) );
  XNOR2XL U39402 ( .A(n51052), .B(n41283), .Y(n29592) );
  XNOR2XL U39403 ( .A(n50624), .B(net219468), .Y(n29593) );
  XNOR2XL U39404 ( .A(n50837), .B(net219308), .Y(n29561) );
  XNOR2XL U39405 ( .A(n51051), .B(n41281), .Y(n29562) );
  XNOR2XL U39406 ( .A(n50623), .B(net219442), .Y(n29563) );
  XNOR2XL U39407 ( .A(n50833), .B(net219308), .Y(n29651) );
  XNOR2XL U39408 ( .A(n51047), .B(n41282), .Y(n29652) );
  XNOR2XL U39409 ( .A(n50619), .B(net219450), .Y(n29653) );
  XNOR2XL U39410 ( .A(n50831), .B(net219310), .Y(n29711) );
  XNOR2XL U39411 ( .A(n51045), .B(n41283), .Y(n29712) );
  XNOR2XL U39412 ( .A(n50617), .B(net219450), .Y(n29713) );
  XOR2XL U39413 ( .A(n42251), .B(n36807), .Y(n22542) );
  XOR2XL U39414 ( .A(n42251), .B(n42490), .Y(n21253) );
  XOR2XL U39415 ( .A(n42248), .B(n42490), .Y(n21273) );
  XOR2XL U39416 ( .A(n42249), .B(n42490), .Y(n21263) );
  XOR2XL U39417 ( .A(n42250), .B(n42490), .Y(n21283) );
  XNOR2XL U39418 ( .A(n50443), .B(n36779), .Y(n24417) );
  XNOR2XL U39419 ( .A(n50444), .B(n36772), .Y(n21254) );
  XNOR2XL U39420 ( .A(n50447), .B(n36771), .Y(n21274) );
  XNOR2XL U39421 ( .A(n50446), .B(n36772), .Y(n21264) );
  XNOR2XL U39422 ( .A(n50445), .B(n36770), .Y(n21284) );
  XNOR2XL U39423 ( .A(n51252), .B(n42697), .Y(n26017) );
  XOR2XL U39424 ( .A(n42258), .B(n41323), .Y(n30329) );
  XOR2XL U39425 ( .A(n42256), .B(n36801), .Y(n30389) );
  XOR2XL U39426 ( .A(n42257), .B(n36873), .Y(n30419) );
  XOR2XL U39427 ( .A(n42259), .B(n41323), .Y(n30359) );
  AND4XL U39428 ( .A(n10751), .B(n10752), .C(n10753), .D(n20960), .Y(n10029)
         );
  NOR2XL U39429 ( .A(net171540), .B(n10699), .Y(n20960) );
  INVXL U39430 ( .A(n10525), .Y(net171134) );
  INVXL U39431 ( .A(n10672), .Y(net151431) );
  INVXL U39432 ( .A(n12896), .Y(net151451) );
  INVXL U39433 ( .A(n12892), .Y(net151453) );
  NAND2XL U39434 ( .A(n11326), .B(n11327), .Y(n11323) );
  INVXL U39435 ( .A(n12800), .Y(net171142) );
  AND3XL U39436 ( .A(n46305), .B(n47802), .C(net209284), .Y(n41788) );
  INVXL U39437 ( .A(n12005), .Y(net171126) );
  NAND3XL U39438 ( .A(n10232), .B(n10233), .C(n10234), .Y(n10229) );
  NOR3XL U39439 ( .A(n46293), .B(net210539), .C(net210561), .Y(n47802) );
  NAND2XL U39440 ( .A(net209277), .B(n41761), .Y(n46293) );
  AND4XL U39441 ( .A(n10184), .B(n39304), .C(net171222), .D(n27614), .Y(n9961)
         );
  NAND2XL U39442 ( .A(n47802), .B(net209284), .Y(n47803) );
  AOI31XL U39443 ( .A0(n47981), .A1(n36936), .A2(n47984), .B0(n47823), .Y(
        n47825) );
  NAND4BBXL U39444 ( .AN(n10150), .BN(n10148), .C(n31886), .D(net261020), .Y(
        n9838) );
  NAND4BXL U39445 ( .AN(net210490), .B(net209902), .C(net209903), .D(n45519),
        .Y(n47835) );
  XNOR2XL U39446 ( .A(n51248), .B(n42697), .Y(n25927) );
  XNOR2XL U39447 ( .A(n51249), .B(n42690), .Y(n25867) );
  XNOR2XL U39448 ( .A(n50185), .B(n42707), .Y(n25715) );
  XNOR2XL U39449 ( .A(n50400), .B(n42720), .Y(n25716) );
  XNOR2XL U39450 ( .A(n51245), .B(n42694), .Y(n25717) );
  INVXL U39451 ( .A(n10483), .Y(net171153) );
  NAND4XL U39452 ( .A(n12154), .B(n12153), .C(n12032), .D(n12033), .Y(n10165)
         );
  NAND4XL U39453 ( .A(net151430), .B(n40388), .C(n10504), .D(n10505), .Y(
        n10150) );
  NAND4BXL U39454 ( .AN(net210543), .B(net209301), .C(net209341), .D(n41763),
        .Y(n47800) );
  NOR2BXL U39455 ( .AN(n10843), .B(n10842), .Y(n24091) );
  XOR2XL U39456 ( .A(n42000), .B(n36756), .Y(n22092) );
  XOR2XL U39457 ( .A(n42033), .B(n41314), .Y(n24659) );
  XOR2XL U39458 ( .A(n41999), .B(n36757), .Y(n22081) );
  XOR2XL U39459 ( .A(n42016), .B(n41317), .Y(n24223) );
  XOR2XL U39460 ( .A(n42017), .B(n41316), .Y(n24203) );
  XOR2XL U39461 ( .A(n42020), .B(n41311), .Y(n24213) );
  XOR2XL U39462 ( .A(n42014), .B(n41313), .Y(n24233) );
  XOR2XL U39463 ( .A(n42035), .B(n41314), .Y(n24637) );
  XOR2XL U39464 ( .A(n42027), .B(n36757), .Y(n20926) );
  XOR2XL U39465 ( .A(n42050), .B(n41317), .Y(n23624) );
  XOR2XL U39466 ( .A(n42051), .B(n41310), .Y(n23614) );
  XOR2XL U39467 ( .A(n42049), .B(n41316), .Y(n23634) );
  XOR2XL U39468 ( .A(n42044), .B(n41312), .Y(n23298) );
  XOR2XL U39469 ( .A(n42042), .B(n41317), .Y(n23308) );
  XOR2XL U39470 ( .A(n42048), .B(n41309), .Y(n23319) );
  XOR2XL U39471 ( .A(n42019), .B(n41312), .Y(n24193) );
  XOR2XL U39472 ( .A(n42018), .B(n41309), .Y(n24183) );
  XNOR2XL U39473 ( .A(n51067), .B(n36718), .Y(n22090) );
  XNOR2XL U39474 ( .A(n51034), .B(n41332), .Y(n24657) );
  XNOR2XL U39475 ( .A(n50639), .B(n42470), .Y(n22091) );
  XNOR2XL U39476 ( .A(n51260), .B(n42696), .Y(n29687) );
  XNOR2XL U39477 ( .A(n50606), .B(n36851), .Y(n24658) );
  XOR2XL U39478 ( .A(n42034), .B(n41310), .Y(n24648) );
  XOR2XL U39479 ( .A(n42041), .B(n41311), .Y(n23288) );
  XNOR2XL U39480 ( .A(n50853), .B(n36799), .Y(n22089) );
  XNOR2XL U39481 ( .A(n50820), .B(n41293), .Y(n24656) );
  XOR2XL U39482 ( .A(n42290), .B(n36882), .Y(n25838) );
  XOR2XL U39483 ( .A(n42031), .B(n36893), .Y(n25834) );
  XOR2XL U39484 ( .A(n42291), .B(n42657), .Y(n25830) );
  XOR2XL U39485 ( .A(n42032), .B(n42606), .Y(n25826) );
  XOR2XL U39486 ( .A(n42293), .B(n36885), .Y(n25898) );
  XOR2XL U39487 ( .A(n42034), .B(n36901), .Y(n25894) );
  XOR2XL U39488 ( .A(n42294), .B(n42656), .Y(n25890) );
  XOR2XL U39489 ( .A(n42035), .B(n36711), .Y(n25886) );
  XOR2XL U39490 ( .A(n42291), .B(n36889), .Y(n25868) );
  XOR2XL U39491 ( .A(n42032), .B(n36897), .Y(n25864) );
  XOR2XL U39492 ( .A(n42292), .B(n42652), .Y(n25860) );
  XOR2XL U39493 ( .A(n42033), .B(n42602), .Y(n25856) );
  XOR2XL U39494 ( .A(n42295), .B(n36882), .Y(n25718) );
  XOR2XL U39495 ( .A(n42036), .B(n36897), .Y(n25714) );
  XOR2XL U39496 ( .A(n42296), .B(n42656), .Y(n25710) );
  XOR2XL U39497 ( .A(n42037), .B(n42606), .Y(n25706) );
  XOR2XL U39498 ( .A(n42294), .B(n36879), .Y(n25748) );
  XOR2XL U39499 ( .A(n42035), .B(n36900), .Y(n25744) );
  XOR2XL U39500 ( .A(n42295), .B(n42663), .Y(n25740) );
  XOR2XL U39501 ( .A(n42036), .B(n42606), .Y(n25736) );
  XOR2XL U39502 ( .A(n42297), .B(n36881), .Y(n25778) );
  XOR2XL U39503 ( .A(n42038), .B(n36900), .Y(n25774) );
  XOR2XL U39504 ( .A(n42298), .B(n42656), .Y(n25770) );
  XOR2XL U39505 ( .A(n42039), .B(n42602), .Y(n25766) );
  XOR2XL U39506 ( .A(n42307), .B(n36886), .Y(n26529) );
  XOR2XL U39507 ( .A(n42048), .B(n36898), .Y(n26525) );
  XOR2XL U39508 ( .A(n42308), .B(n42663), .Y(n26521) );
  XOR2XL U39509 ( .A(n42049), .B(n42597), .Y(n26517) );
  XOR2XL U39510 ( .A(n42306), .B(n36883), .Y(n26499) );
  XOR2XL U39511 ( .A(n42047), .B(n36892), .Y(n26495) );
  XOR2XL U39512 ( .A(n42307), .B(n42663), .Y(n26491) );
  XOR2XL U39513 ( .A(n42048), .B(n42611), .Y(n26487) );
  XOR2XL U39514 ( .A(n42296), .B(n36886), .Y(n25808) );
  XOR2XL U39515 ( .A(n42037), .B(n36891), .Y(n25804) );
  XOR2XL U39516 ( .A(n42297), .B(n42656), .Y(n25800) );
  XOR2XL U39517 ( .A(n42038), .B(n36711), .Y(n25796) );
  XOR2XL U39518 ( .A(n42305), .B(n36887), .Y(n26378) );
  XOR2XL U39519 ( .A(n42046), .B(n36897), .Y(n26374) );
  XOR2XL U39520 ( .A(n42306), .B(n42652), .Y(n26370) );
  XOR2XL U39521 ( .A(n42047), .B(n42601), .Y(n26366) );
  XOR2XL U39522 ( .A(n42304), .B(n36880), .Y(n26408) );
  XOR2XL U39523 ( .A(n42305), .B(n42667), .Y(n26400) );
  XOR2XL U39524 ( .A(n42046), .B(n42612), .Y(n26396) );
  XOR2XL U39525 ( .A(n42045), .B(n36891), .Y(n26404) );
  XOR2XL U39526 ( .A(n42312), .B(n36887), .Y(n26559) );
  XOR2XL U39527 ( .A(n42053), .B(n36895), .Y(n26555) );
  XOR2XL U39528 ( .A(n42313), .B(n42663), .Y(n26551) );
  XOR2XL U39529 ( .A(n42054), .B(n42605), .Y(n26547) );
  XOR2XL U39530 ( .A(n42302), .B(n36885), .Y(n26348) );
  XOR2XL U39531 ( .A(n42043), .B(n36898), .Y(n26344) );
  XOR2XL U39532 ( .A(n42303), .B(n42663), .Y(n26340) );
  XOR2XL U39533 ( .A(n42044), .B(n42605), .Y(n26336) );
  XOR2XL U39534 ( .A(n42309), .B(n36880), .Y(n26439) );
  XOR2XL U39535 ( .A(n42050), .B(n36893), .Y(n26435) );
  XOR2XL U39536 ( .A(n42310), .B(n42665), .Y(n26431) );
  XOR2XL U39537 ( .A(n42051), .B(n42605), .Y(n26427) );
  XOR2XL U39538 ( .A(n42310), .B(n36886), .Y(n26619) );
  XOR2XL U39539 ( .A(n42051), .B(n36899), .Y(n26615) );
  XOR2XL U39540 ( .A(n42311), .B(n42661), .Y(n26611) );
  XOR2XL U39541 ( .A(n42052), .B(n42607), .Y(n26607) );
  XOR2XL U39542 ( .A(n42303), .B(n36887), .Y(n26318) );
  XOR2XL U39543 ( .A(n42044), .B(n36898), .Y(n26314) );
  XOR2XL U39544 ( .A(n42304), .B(n42663), .Y(n26310) );
  XOR2XL U39545 ( .A(n42045), .B(n42597), .Y(n26306) );
  XOR2XL U39546 ( .A(n42311), .B(n36882), .Y(n26649) );
  XOR2XL U39547 ( .A(n42052), .B(n36900), .Y(n26645) );
  XOR2XL U39548 ( .A(n42312), .B(n42664), .Y(n26641) );
  XOR2XL U39549 ( .A(n42053), .B(n42607), .Y(n26637) );
  XOR2XL U39550 ( .A(n42308), .B(n36886), .Y(n26469) );
  XOR2XL U39551 ( .A(n42049), .B(n36895), .Y(n26465) );
  XOR2XL U39552 ( .A(n42309), .B(n42663), .Y(n26461) );
  XOR2XL U39553 ( .A(n42050), .B(n42604), .Y(n26457) );
  XNOR2XL U39554 ( .A(n51281), .B(n36746), .Y(n22094) );
  XNOR2XL U39555 ( .A(n51248), .B(n41302), .Y(n24661) );
  XNOR2XL U39556 ( .A(n51245), .B(n41300), .Y(n24629) );
  XNOR2XL U39557 ( .A(n51246), .B(n41299), .Y(n24640) );
  XOR2XL U39558 ( .A(n42019), .B(n42522), .Y(n29516) );
  XOR2XL U39559 ( .A(n42020), .B(n42516), .Y(n29486) );
  XOR2XL U39560 ( .A(n42033), .B(n42524), .Y(n25816) );
  XOR2XL U39561 ( .A(n42031), .B(n42524), .Y(n25996) );
  XOR2XL U39562 ( .A(n42029), .B(n42524), .Y(n25936) );
  XOR2XL U39563 ( .A(n42030), .B(n42524), .Y(n25966) );
  XOR2XL U39564 ( .A(n42034), .B(n42524), .Y(n25846) );
  XOR2XL U39565 ( .A(n42035), .B(n42524), .Y(n25906) );
  XOR2XL U39566 ( .A(n42036), .B(n42524), .Y(n25876) );
  XOR2XL U39567 ( .A(n42038), .B(n42524), .Y(n25696) );
  XOR2XL U39568 ( .A(n42037), .B(n42524), .Y(n25726) );
  XOR2XL U39569 ( .A(n42040), .B(n42524), .Y(n25756) );
  XOR2XL U39570 ( .A(n42039), .B(n42524), .Y(n25786) );
  XOR2XL U39571 ( .A(n42050), .B(n42522), .Y(n26507) );
  XOR2XL U39572 ( .A(n42049), .B(n42522), .Y(n26477) );
  XOR2XL U39573 ( .A(n42047), .B(n42522), .Y(n26386) );
  XOR2XL U39574 ( .A(n42051), .B(n42522), .Y(n26447) );
  XNOR2XL U39575 ( .A(n51068), .B(n36716), .Y(n22079) );
  XNOR2XL U39576 ( .A(n51051), .B(n41330), .Y(n24221) );
  XNOR2XL U39577 ( .A(n51050), .B(n41328), .Y(n24201) );
  XNOR2XL U39578 ( .A(n51047), .B(n41332), .Y(n24211) );
  XNOR2XL U39579 ( .A(n51053), .B(n41327), .Y(n24231) );
  XNOR2XL U39580 ( .A(n51032), .B(n41330), .Y(n24635) );
  XNOR2XL U39581 ( .A(n51039), .B(n36722), .Y(n20914) );
  XNOR2XL U39582 ( .A(n51017), .B(n41333), .Y(n23622) );
  XNOR2XL U39583 ( .A(n51016), .B(n41327), .Y(n23612) );
  XNOR2XL U39584 ( .A(n51018), .B(n41331), .Y(n23632) );
  XNOR2XL U39585 ( .A(n51023), .B(n41327), .Y(n23296) );
  XNOR2XL U39586 ( .A(n51025), .B(n41332), .Y(n23306) );
  XNOR2XL U39587 ( .A(n51019), .B(n41327), .Y(n23317) );
  XNOR2XL U39588 ( .A(n51020), .B(n41330), .Y(n23327) );
  XNOR2XL U39589 ( .A(n51048), .B(n41329), .Y(n24191) );
  XNOR2XL U39590 ( .A(n51049), .B(n41328), .Y(n24181) );
  XNOR2XL U39591 ( .A(n50640), .B(n42459), .Y(n22080) );
  XNOR2XL U39592 ( .A(n50623), .B(n36853), .Y(n24222) );
  XNOR2XL U39593 ( .A(n50622), .B(n36854), .Y(n24202) );
  XNOR2XL U39594 ( .A(n50619), .B(n36860), .Y(n24212) );
  XNOR2XL U39595 ( .A(n50625), .B(n36850), .Y(n24232) );
  XNOR2XL U39596 ( .A(n50604), .B(n36856), .Y(n24636) );
  XNOR2XL U39597 ( .A(n50611), .B(n42459), .Y(n20915) );
  XNOR2XL U39598 ( .A(n50589), .B(n36860), .Y(n23623) );
  XNOR2XL U39599 ( .A(n50588), .B(n36852), .Y(n23613) );
  XNOR2XL U39600 ( .A(n50590), .B(n36856), .Y(n23633) );
  XNOR2XL U39601 ( .A(n50595), .B(n36858), .Y(n23297) );
  XNOR2XL U39602 ( .A(n50597), .B(n36860), .Y(n23307) );
  XNOR2XL U39603 ( .A(n50591), .B(n36859), .Y(n23318) );
  XNOR2XL U39604 ( .A(n50620), .B(n36850), .Y(n24192) );
  XNOR2XL U39605 ( .A(n50621), .B(n36854), .Y(n24182) );
  XNOR2XL U39606 ( .A(n50211), .B(n42711), .Y(n29806) );
  XNOR2XL U39607 ( .A(n50210), .B(n42671), .Y(n29798) );
  XNOR2XL U39608 ( .A(n50203), .B(n42711), .Y(n29505) );
  XNOR2XL U39609 ( .A(n50202), .B(n42671), .Y(n29497) );
  XNOR2XL U39610 ( .A(n50214), .B(n42712), .Y(n29776) );
  XNOR2XL U39611 ( .A(n50213), .B(n42671), .Y(n29768) );
  XNOR2XL U39612 ( .A(n50845), .B(n42615), .Y(n29764) );
  XNOR2XL U39613 ( .A(n50213), .B(n42704), .Y(n29746) );
  XNOR2XL U39614 ( .A(n50212), .B(n42671), .Y(n29738) );
  XNOR2XL U39615 ( .A(n50206), .B(n42706), .Y(n29595) );
  XNOR2XL U39616 ( .A(n50205), .B(n42671), .Y(n29587) );
  XNOR2XL U39617 ( .A(n50837), .B(n42615), .Y(n29583) );
  XNOR2XL U39618 ( .A(n50205), .B(n42711), .Y(n29565) );
  XNOR2XL U39619 ( .A(n50204), .B(n42671), .Y(n29557) );
  XNOR2XL U39620 ( .A(n50836), .B(n42615), .Y(n29553) );
  XNOR2XL U39621 ( .A(n50204), .B(n42706), .Y(n29535) );
  XNOR2XL U39622 ( .A(n50203), .B(n42671), .Y(n29527) );
  XNOR2XL U39623 ( .A(n50835), .B(n42615), .Y(n29523) );
  XNOR2XL U39624 ( .A(n50201), .B(n42704), .Y(n29655) );
  XNOR2XL U39625 ( .A(n50200), .B(n42671), .Y(n29647) );
  XNOR2XL U39626 ( .A(n50832), .B(n42615), .Y(n29643) );
  XNOR2XL U39627 ( .A(n50200), .B(n42704), .Y(n29685) );
  XNOR2XL U39628 ( .A(n50199), .B(n42671), .Y(n29677) );
  XNOR2XL U39629 ( .A(n50831), .B(n42615), .Y(n29673) );
  XNOR2XL U39630 ( .A(n50199), .B(n42705), .Y(n29715) );
  XNOR2XL U39631 ( .A(n50198), .B(n42671), .Y(n29707) );
  XNOR2XL U39632 ( .A(n50830), .B(n42615), .Y(n29703) );
  XNOR2XL U39633 ( .A(n50822), .B(net219308), .Y(n25831) );
  XNOR2XL U39634 ( .A(n50188), .B(n42670), .Y(n25857) );
  XNOR2XL U39635 ( .A(n50820), .B(n42615), .Y(n25853) );
  XNOR2XL U39636 ( .A(n50817), .B(net219310), .Y(n25711) );
  XNOR2XL U39637 ( .A(n50184), .B(n42671), .Y(n25707) );
  XNOR2XL U39638 ( .A(n50816), .B(n42615), .Y(n25703) );
  XNOR2XL U39639 ( .A(n50818), .B(net219310), .Y(n25741) );
  XNOR2XL U39640 ( .A(n50185), .B(n42672), .Y(n25737) );
  XNOR2XL U39641 ( .A(n50817), .B(n42613), .Y(n25733) );
  XNOR2XL U39642 ( .A(n50802), .B(n40039), .Y(n26612) );
  XNOR2XL U39643 ( .A(n50169), .B(n42671), .Y(n26608) );
  XNOR2XL U39644 ( .A(n50801), .B(n42615), .Y(n26604) );
  XNOR2XL U39645 ( .A(n50801), .B(net219336), .Y(n26642) );
  XNOR2XL U39646 ( .A(n50168), .B(n42669), .Y(n26638) );
  XNOR2XL U39647 ( .A(n50800), .B(n42615), .Y(n26634) );
  XNOR2XL U39648 ( .A(n50854), .B(n36793), .Y(n22078) );
  XNOR2XL U39649 ( .A(n50837), .B(n41294), .Y(n24220) );
  XNOR2XL U39650 ( .A(n50836), .B(n41290), .Y(n24200) );
  XNOR2XL U39651 ( .A(n50833), .B(n41295), .Y(n24210) );
  XNOR2XL U39652 ( .A(n50839), .B(n41292), .Y(n24230) );
  XNOR2XL U39653 ( .A(n50827), .B(n36790), .Y(n20902) );
  XNOR2XL U39654 ( .A(n50818), .B(n41294), .Y(n24634) );
  XNOR2XL U39655 ( .A(n50825), .B(n36791), .Y(n20913) );
  XNOR2XL U39656 ( .A(n50803), .B(n41297), .Y(n23621) );
  XNOR2XL U39657 ( .A(n50802), .B(n41291), .Y(n23611) );
  XNOR2XL U39658 ( .A(n50804), .B(n41294), .Y(n23631) );
  XNOR2XL U39659 ( .A(n50809), .B(n41297), .Y(n23295) );
  XNOR2XL U39660 ( .A(n50811), .B(n41295), .Y(n23305) );
  XNOR2XL U39661 ( .A(n50805), .B(n41291), .Y(n23316) );
  XNOR2XL U39662 ( .A(n50806), .B(n41294), .Y(n23326) );
  XNOR2XL U39663 ( .A(n50834), .B(n41291), .Y(n24190) );
  XNOR2XL U39664 ( .A(n50835), .B(n41291), .Y(n24180) );
  XNOR2XL U39665 ( .A(n50628), .B(n42586), .Y(n29796) );
  XNOR2XL U39666 ( .A(n51058), .B(n42552), .Y(n29755) );
  XNOR2XL U39667 ( .A(n51055), .B(n42552), .Y(n29785) );
  XNOR2XL U39668 ( .A(n51056), .B(n42552), .Y(n29815) );
  XNOR2XL U39669 ( .A(n50620), .B(n42586), .Y(n29495) );
  XNOR2XL U39670 ( .A(n51048), .B(n42553), .Y(n29514) );
  XNOR2XL U39671 ( .A(n51047), .B(n42552), .Y(n29484) );
  XNOR2XL U39672 ( .A(n51046), .B(n42553), .Y(n29604) );
  XNOR2XL U39673 ( .A(n51273), .B(n42638), .Y(n29770) );
  XNOR2XL U39674 ( .A(n50631), .B(n42586), .Y(n29766) );
  XNOR2XL U39675 ( .A(n50630), .B(n42586), .Y(n29736) );
  XNOR2XL U39676 ( .A(n51057), .B(n42550), .Y(n29725) );
  XNOR2XL U39677 ( .A(n51265), .B(n42644), .Y(n29589) );
  XNOR2XL U39678 ( .A(n50623), .B(n42586), .Y(n29585) );
  XNOR2XL U39679 ( .A(n51264), .B(n42644), .Y(n29559) );
  XNOR2XL U39680 ( .A(n50622), .B(n42586), .Y(n29555) );
  XNOR2XL U39681 ( .A(n51263), .B(n42638), .Y(n29529) );
  XNOR2XL U39682 ( .A(n50621), .B(n42586), .Y(n29525) );
  XNOR2XL U39683 ( .A(n51260), .B(n36867), .Y(n29649) );
  XNOR2XL U39684 ( .A(n50618), .B(n42586), .Y(n29645) );
  XNOR2XL U39685 ( .A(n51259), .B(n36867), .Y(n29679) );
  XNOR2XL U39686 ( .A(n50617), .B(n42586), .Y(n29675) );
  XNOR2XL U39687 ( .A(n51258), .B(n42638), .Y(n29709) );
  XNOR2XL U39688 ( .A(n50616), .B(n42586), .Y(n29705) );
  XNOR2XL U39689 ( .A(n50608), .B(net219434), .Y(n25833) );
  XNOR2XL U39690 ( .A(n51246), .B(n36867), .Y(n25889) );
  XNOR2XL U39691 ( .A(n50604), .B(n36865), .Y(n25885) );
  XNOR2XL U39692 ( .A(n51049), .B(n42552), .Y(n29544) );
  XNOR2XL U39693 ( .A(n51050), .B(n42552), .Y(n29574) );
  XNOR2XL U39694 ( .A(n50603), .B(net219434), .Y(n25713) );
  XNOR2XL U39695 ( .A(n51244), .B(n36867), .Y(n25709) );
  XNOR2XL U39696 ( .A(n50602), .B(n42586), .Y(n25705) );
  XNOR2XL U39697 ( .A(n51245), .B(n36867), .Y(n25739) );
  XNOR2XL U39698 ( .A(n50603), .B(n42590), .Y(n25735) );
  XNOR2XL U39699 ( .A(n51044), .B(n42552), .Y(n29664) );
  XNOR2XL U39700 ( .A(n51043), .B(n42552), .Y(n29694) );
  XNOR2XL U39701 ( .A(n51045), .B(n42548), .Y(n29634) );
  XNOR2XL U39702 ( .A(n51029), .B(n42551), .Y(n25694) );
  XNOR2XL U39703 ( .A(n51030), .B(n42552), .Y(n25724) );
  XNOR2XL U39704 ( .A(n50586), .B(net219434), .Y(n26554) );
  XNOR2XL U39705 ( .A(n50588), .B(net219434), .Y(n26614) );
  XNOR2XL U39706 ( .A(n51229), .B(n36867), .Y(n26610) );
  XNOR2XL U39707 ( .A(n50587), .B(n36865), .Y(n26606) );
  XNOR2XL U39708 ( .A(n50587), .B(net219434), .Y(n26644) );
  XNOR2XL U39709 ( .A(n50586), .B(n36865), .Y(n26636) );
  XNOR2XL U39710 ( .A(n50425), .B(n36728), .Y(n29799) );
  XNOR2XL U39711 ( .A(n50417), .B(n36728), .Y(n29498) );
  XNOR2XL U39712 ( .A(n50620), .B(n42502), .Y(n29515) );
  XNOR2XL U39713 ( .A(n50619), .B(n42502), .Y(n29485) );
  XNOR2XL U39714 ( .A(n50428), .B(n36728), .Y(n29769) );
  XNOR2XL U39715 ( .A(n51059), .B(n42631), .Y(n29765) );
  XNOR2XL U39716 ( .A(n50427), .B(n36728), .Y(n29739) );
  XNOR2XL U39717 ( .A(n50420), .B(n36728), .Y(n29588) );
  XNOR2XL U39718 ( .A(n51051), .B(n42633), .Y(n29584) );
  XNOR2XL U39719 ( .A(n50419), .B(n36728), .Y(n29558) );
  XNOR2XL U39720 ( .A(n51050), .B(n42628), .Y(n29554) );
  XNOR2XL U39721 ( .A(n50419), .B(n36875), .Y(n29536) );
  XNOR2XL U39722 ( .A(n50418), .B(n36728), .Y(n29528) );
  XNOR2XL U39723 ( .A(n51049), .B(n42633), .Y(n29524) );
  XNOR2XL U39724 ( .A(n50416), .B(n42717), .Y(n29656) );
  XNOR2XL U39725 ( .A(n50415), .B(n36728), .Y(n29648) );
  XNOR2XL U39726 ( .A(n51046), .B(n42632), .Y(n29644) );
  XNOR2XL U39727 ( .A(n50415), .B(n36875), .Y(n29686) );
  XNOR2XL U39728 ( .A(n50414), .B(n36728), .Y(n29678) );
  XNOR2XL U39729 ( .A(n51045), .B(n42633), .Y(n29674) );
  XNOR2XL U39730 ( .A(n50413), .B(n36728), .Y(n29708) );
  XNOR2XL U39731 ( .A(n51044), .B(n42624), .Y(n29704) );
  XNOR2XL U39732 ( .A(n51036), .B(n41282), .Y(n25832) );
  XNOR2XL U39733 ( .A(n51032), .B(n34447), .Y(n25884) );
  XNOR2XL U39734 ( .A(n50403), .B(n36903), .Y(n25858) );
  XNOR2XL U39735 ( .A(n51031), .B(n41283), .Y(n25712) );
  XNOR2XL U39736 ( .A(n50399), .B(n41379), .Y(n25708) );
  XNOR2XL U39737 ( .A(n51030), .B(n42629), .Y(n25704) );
  XNOR2XL U39738 ( .A(n50400), .B(n41319), .Y(n25738) );
  XNOR2XL U39739 ( .A(n51031), .B(n42629), .Y(n25734) );
  XNOR2XL U39740 ( .A(n50601), .B(n36730), .Y(n25695) );
  XNOR2XL U39741 ( .A(n50602), .B(n36731), .Y(n25725) );
  XNOR2XL U39742 ( .A(n50599), .B(n36730), .Y(n25755) );
  XNOR2XL U39743 ( .A(n50600), .B(n36730), .Y(n25785) );
  XNOR2XL U39744 ( .A(n51016), .B(n41282), .Y(n26613) );
  XNOR2XL U39745 ( .A(n50384), .B(n41380), .Y(n26609) );
  XNOR2XL U39746 ( .A(n51015), .B(n42630), .Y(n26605) );
  XNOR2XL U39747 ( .A(n51015), .B(n41281), .Y(n26643) );
  XNOR2XL U39748 ( .A(n50383), .B(n36905), .Y(n26639) );
  XNOR2XL U39749 ( .A(n51014), .B(n42630), .Y(n26635) );
  XNOR2XL U39750 ( .A(n51033), .B(n41330), .Y(n24646) );
  XNOR2XL U39751 ( .A(n51026), .B(n41328), .Y(n23286) );
  NAND3XL U39752 ( .A(n10272), .B(n10273), .C(n10274), .Y(n10222) );
  XNOR2XL U39753 ( .A(n50605), .B(n36850), .Y(n24647) );
  XNOR2XL U39754 ( .A(n50598), .B(n36850), .Y(n23287) );
  XNOR2XL U39755 ( .A(n50832), .B(net219310), .Y(n29681) );
  XNOR2XL U39756 ( .A(n51046), .B(n41281), .Y(n29682) );
  XNOR2XL U39757 ( .A(n50618), .B(net219450), .Y(n29683) );
  XOR2XL U39758 ( .A(n42259), .B(n42493), .Y(n22093) );
  XOR2XL U39759 ( .A(n42292), .B(n36808), .Y(n24660) );
  XOR2XL U39760 ( .A(n42258), .B(n42483), .Y(n22082) );
  XOR2XL U39761 ( .A(n42275), .B(n36813), .Y(n24224) );
  XOR2XL U39762 ( .A(n42276), .B(n36809), .Y(n24204) );
  XOR2XL U39763 ( .A(n42279), .B(n36813), .Y(n24214) );
  XOR2XL U39764 ( .A(n42273), .B(n36810), .Y(n24234) );
  XOR2XL U39765 ( .A(n42285), .B(n42483), .Y(n20906) );
  XOR2XL U39766 ( .A(n42294), .B(n36814), .Y(n24638) );
  XOR2XL U39767 ( .A(n42286), .B(n42483), .Y(n20927) );
  XOR2XL U39768 ( .A(n42309), .B(n36809), .Y(n23625) );
  XOR2XL U39769 ( .A(n42310), .B(n36810), .Y(n23615) );
  XOR2XL U39770 ( .A(n42308), .B(n36814), .Y(n23635) );
  XOR2XL U39771 ( .A(n42303), .B(n36817), .Y(n23299) );
  XOR2XL U39772 ( .A(n42301), .B(n36808), .Y(n23309) );
  XOR2XL U39773 ( .A(n42307), .B(n36813), .Y(n23320) );
  XOR2XL U39774 ( .A(n42278), .B(n36811), .Y(n24194) );
  XOR2XL U39775 ( .A(n42277), .B(n36808), .Y(n24184) );
  XNOR2XL U39776 ( .A(n50815), .B(n42540), .Y(n25693) );
  XNOR2XL U39777 ( .A(n50816), .B(n42539), .Y(n25723) );
  XNOR2XL U39778 ( .A(n50813), .B(n42539), .Y(n25753) );
  XNOR2XL U39779 ( .A(n50819), .B(n41296), .Y(n24645) );
  XNOR2XL U39780 ( .A(n50812), .B(n41291), .Y(n23285) );
  XOR2XL U39781 ( .A(n42293), .B(n36814), .Y(n24649) );
  XOR2XL U39782 ( .A(n42300), .B(n36808), .Y(n23289) );
  XNOR2XL U39783 ( .A(n50427), .B(n36786), .Y(n24275) );
  XNOR2XL U39784 ( .A(n51265), .B(n41301), .Y(n24225) );
  XNOR2XL U39785 ( .A(n50429), .B(n36785), .Y(n24355) );
  XNOR2XL U39786 ( .A(n50428), .B(n36777), .Y(n24345) );
  XNOR2XL U39787 ( .A(n51264), .B(n41304), .Y(n24205) );
  XNOR2XL U39788 ( .A(n50416), .B(n36777), .Y(n24215) );
  XNOR2XL U39789 ( .A(n50415), .B(n36780), .Y(n24335) );
  XNOR2XL U39790 ( .A(n51267), .B(n41302), .Y(n24235) );
  XNOR2XL U39791 ( .A(n50414), .B(n36782), .Y(n24325) );
  XNOR2XL U39792 ( .A(n50414), .B(n36772), .Y(n21892) );
  XNOR2XL U39793 ( .A(n50413), .B(n36783), .Y(n24305) );
  XNOR2XL U39794 ( .A(n50411), .B(n36783), .Y(n24609) );
  XNOR2XL U39795 ( .A(n50413), .B(n36766), .Y(n21872) );
  XNOR2XL U39796 ( .A(n51247), .B(n41303), .Y(n24651) );
  XNOR2XL U39797 ( .A(n51254), .B(n36744), .Y(n20929) );
  XNOR2XL U39798 ( .A(n50386), .B(n36779), .Y(n23626) );
  XNOR2XL U39799 ( .A(n50398), .B(n36778), .Y(n24537) );
  XNOR2XL U39800 ( .A(n50395), .B(n36780), .Y(n23290) );
  XNOR2XL U39801 ( .A(n50385), .B(n36782), .Y(n23616) );
  XNOR2XL U39802 ( .A(n51237), .B(n41303), .Y(n23300) );
  XNOR2XL U39803 ( .A(n51239), .B(n41303), .Y(n23311) );
  XNOR2XL U39804 ( .A(n50388), .B(n36778), .Y(n23321) );
  XNOR2XL U39805 ( .A(n50417), .B(n36784), .Y(n24195) );
  XNOR2XL U39806 ( .A(n50418), .B(n36784), .Y(n24185) );
  XOR2XL U39807 ( .A(n42026), .B(n36757), .Y(n20905) );
  XNOR2XL U39808 ( .A(n50613), .B(n42459), .Y(n20904) );
  XNOR2XL U39809 ( .A(n51041), .B(n36717), .Y(n20903) );
  XNOR2XL U39810 ( .A(n51254), .B(n42697), .Y(n25957) );
  XNOR2XL U39811 ( .A(n51253), .B(n42690), .Y(n25987) );
  XNOR2XL U39812 ( .A(n50190), .B(n42706), .Y(n25835) );
  XNOR2XL U39813 ( .A(n50405), .B(n42717), .Y(n25836) );
  XNOR2XL U39814 ( .A(n51250), .B(n42690), .Y(n25837) );
  XNOR2XL U39815 ( .A(n51247), .B(n42694), .Y(n25897) );
  XNOR2XL U39816 ( .A(n50186), .B(n42707), .Y(n25745) );
  XNOR2XL U39817 ( .A(n50401), .B(n42720), .Y(n25746) );
  XNOR2XL U39818 ( .A(n51246), .B(n42694), .Y(n25747) );
  XNOR2XL U39819 ( .A(n51243), .B(n42694), .Y(n25777) );
  XNOR2XL U39820 ( .A(n51233), .B(n42696), .Y(n26528) );
  XNOR2XL U39821 ( .A(n51234), .B(n42696), .Y(n26498) );
  XNOR2XL U39822 ( .A(n51244), .B(n42696), .Y(n25807) );
  XNOR2XL U39823 ( .A(n51228), .B(n42696), .Y(n26558) );
  XNOR2XL U39824 ( .A(n50170), .B(n42709), .Y(n26616) );
  XNOR2XL U39825 ( .A(n50385), .B(n34435), .Y(n26617) );
  XNOR2XL U39826 ( .A(n51230), .B(n42696), .Y(n26618) );
  XNOR2XL U39827 ( .A(n50169), .B(n42708), .Y(n26646) );
  XNOR2XL U39828 ( .A(n50384), .B(n34435), .Y(n26647) );
  XNOR2XL U39829 ( .A(n51229), .B(n42696), .Y(n26648) );
  XNOR2XL U39830 ( .A(n51232), .B(n42696), .Y(n26468) );
  XNOR2XL U39831 ( .A(n51282), .B(n36742), .Y(n22084) );
  XNOR2XL U39832 ( .A(n50398), .B(n42576), .Y(n25698) );
  XNOR2XL U39833 ( .A(n50399), .B(n42580), .Y(n25728) );
  XNOR2XL U39834 ( .A(n50396), .B(n42580), .Y(n25758) );
  NAND3XL U39835 ( .A(net234760), .B(n37469), .C(net209930), .Y(n47836) );
  XOR2XL U39836 ( .A(n42278), .B(n36873), .Y(n29517) );
  XOR2XL U39837 ( .A(n42279), .B(n36873), .Y(n29487) );
  XOR2XL U39838 ( .A(n42292), .B(n41322), .Y(n25817) );
  XOR2XL U39839 ( .A(n42290), .B(n36801), .Y(n25997) );
  XOR2XL U39840 ( .A(n42288), .B(n41322), .Y(n25937) );
  XOR2XL U39841 ( .A(n42289), .B(n41323), .Y(n25967) );
  XOR2XL U39842 ( .A(n42293), .B(n36877), .Y(n25847) );
  XOR2XL U39843 ( .A(n42294), .B(n36873), .Y(n25907) );
  XOR2XL U39844 ( .A(n42295), .B(n41323), .Y(n25877) );
  XOR2XL U39845 ( .A(n42297), .B(n36801), .Y(n25697) );
  XOR2XL U39846 ( .A(n42296), .B(n41321), .Y(n25727) );
  XOR2XL U39847 ( .A(n42299), .B(n36801), .Y(n25757) );
  XOR2XL U39848 ( .A(n42298), .B(n41321), .Y(n25787) );
  XOR2XL U39849 ( .A(n42309), .B(n36801), .Y(n26508) );
  XOR2XL U39850 ( .A(n42308), .B(n36877), .Y(n26478) );
  XOR2XL U39851 ( .A(n42306), .B(n36873), .Y(n26387) );
  XOR2XL U39852 ( .A(n42310), .B(n36873), .Y(n26448) );
  NOR3XL U39853 ( .A(n47809), .B(net209899), .C(n47808), .Y(n47811) );
  AND4XL U39854 ( .A(n10863), .B(n10872), .C(n10870), .D(n10869), .Y(n23687)
         );
  NOR4XL U39855 ( .A(net171430), .B(net209254), .C(net171433), .D(net171435),
        .Y(n23688) );
  NAND4BXL U39856 ( .AN(n10040), .B(n10045), .C(n37018), .D(n10044), .Y(n47826) );
  NAND4XL U39857 ( .A(net260247), .B(net260251), .C(net260427), .D(n30683),
        .Y(n9954) );
  NAND2XL U39858 ( .A(n11978), .B(n11979), .Y(n11975) );
  INVXL U39859 ( .A(n10810), .Y(net171476) );
  OAI211XL U39860 ( .A0(n9886), .A1(n10011), .B0(n10012), .C0(n40405), .Y(
        n10007) );
  INVXL U39861 ( .A(n10808), .Y(net171478) );
  NAND4XL U39862 ( .A(n10487), .B(n10485), .C(net260431), .D(n30442), .Y(n9837) );
  AND3XL U39863 ( .A(n10481), .B(n40389), .C(n37347), .Y(n30442) );
  NAND4XL U39864 ( .A(n10567), .B(n10566), .C(n12793), .D(n27132), .Y(n9964)
         );
  NOR3XL U39865 ( .A(n10570), .B(net171240), .C(n10572), .Y(n27132) );
  NAND4BXL U39866 ( .AN(n10577), .B(n12085), .C(n12749), .D(n27373), .Y(n9963)
         );
  NOR4XL U39867 ( .A(net151705), .B(net209846), .C(net171233), .D(net171234),
        .Y(n27373) );
  XOR2XL U39868 ( .A(n42052), .B(n36759), .Y(n20442) );
  XOR2XL U39869 ( .A(n42050), .B(n36761), .Y(n20463) );
  XOR2XL U39870 ( .A(n42051), .B(n36760), .Y(n20452) );
  XOR2XL U39871 ( .A(n42054), .B(n36756), .Y(n20504) );
  XOR2XL U39872 ( .A(n42056), .B(n36759), .Y(n20432) );
  XOR2XL U39873 ( .A(n42049), .B(n36755), .Y(n20474) );
  XOR2XL U39874 ( .A(n42055), .B(n36754), .Y(n20484) );
  XOR2XL U39875 ( .A(n42010), .B(n36757), .Y(n21798) );
  XOR2XL U39876 ( .A(n42009), .B(n36759), .Y(n21809) );
  XOR2XL U39877 ( .A(n42011), .B(n36761), .Y(n21787) );
  XOR2XL U39878 ( .A(n42012), .B(n36753), .Y(n21777) );
  XOR2XL U39879 ( .A(n42031), .B(n36756), .Y(n20947) );
  XOR2XL U39880 ( .A(n42032), .B(n36754), .Y(n20937) );
  XOR2XL U39881 ( .A(n42041), .B(n36756), .Y(n20053) );
  XOR2XL U39882 ( .A(n42042), .B(n36755), .Y(n20043) );
  XOR2XL U39883 ( .A(n42053), .B(n41317), .Y(n23674) );
  XOR2XL U39884 ( .A(n42054), .B(n41311), .Y(n23684) );
  XOR2XL U39885 ( .A(n42046), .B(n41316), .Y(n23350) );
  XOR2XL U39886 ( .A(n42045), .B(n41309), .Y(n23360) );
  XOR2XL U39887 ( .A(n42037), .B(n36757), .Y(n20800) );
  XOR2XL U39888 ( .A(n42052), .B(n41314), .Y(n23644) );
  XOR2XL U39889 ( .A(n42025), .B(n36754), .Y(n20957) );
  XOR2XL U39890 ( .A(n42043), .B(n36755), .Y(n20033) );
  XOR2XL U39891 ( .A(n42043), .B(n41312), .Y(n23339) );
  XOR2XL U39892 ( .A(n42047), .B(n41318), .Y(n23329) );
  XOR2XL U39893 ( .A(n42053), .B(n36753), .Y(n20494) );
  XOR2XL U39894 ( .A(n42044), .B(n36760), .Y(n20023) );
  XOR2XL U39895 ( .A(n42046), .B(n36760), .Y(n20073) );
  XOR2XL U39896 ( .A(n42045), .B(n36759), .Y(n20063) );
  XOR2XL U39897 ( .A(n42048), .B(n36755), .Y(n20083) );
  XOR2XL U39898 ( .A(n42047), .B(n36761), .Y(n20093) );
  XOR2XL U39899 ( .A(n42055), .B(n41318), .Y(n23664) );
  XOR2XL U39900 ( .A(n42056), .B(n41311), .Y(n23654) );
  XNOR2XL U39901 ( .A(n51015), .B(n36714), .Y(n20440) );
  XNOR2XL U39902 ( .A(n51017), .B(n36715), .Y(n20461) );
  XNOR2XL U39903 ( .A(n51016), .B(n36714), .Y(n20450) );
  XNOR2XL U39904 ( .A(n51013), .B(n36720), .Y(n20502) );
  XNOR2XL U39905 ( .A(n51011), .B(n36718), .Y(n20430) );
  XNOR2XL U39906 ( .A(n51018), .B(n36722), .Y(n20472) );
  XNOR2XL U39907 ( .A(n51012), .B(n36716), .Y(n20482) );
  XNOR2XL U39908 ( .A(n50587), .B(n42470), .Y(n20441) );
  XNOR2XL U39909 ( .A(n50589), .B(n42470), .Y(n20462) );
  XNOR2XL U39910 ( .A(n50588), .B(n42470), .Y(n20451) );
  XNOR2XL U39911 ( .A(n50585), .B(n42470), .Y(n20503) );
  XNOR2XL U39912 ( .A(n50583), .B(n42470), .Y(n20431) );
  XNOR2XL U39913 ( .A(n50590), .B(n42470), .Y(n20473) );
  XNOR2XL U39914 ( .A(n50584), .B(n42470), .Y(n20483) );
  XNOR2XL U39915 ( .A(n50801), .B(n36792), .Y(n20439) );
  XNOR2XL U39916 ( .A(n50803), .B(n36797), .Y(n20460) );
  XNOR2XL U39917 ( .A(n50802), .B(n36796), .Y(n20449) );
  XNOR2XL U39918 ( .A(n50799), .B(n36797), .Y(n20501) );
  XNOR2XL U39919 ( .A(n50797), .B(n36792), .Y(n20429) );
  XNOR2XL U39920 ( .A(n50804), .B(n36790), .Y(n20471) );
  XNOR2XL U39921 ( .A(n50798), .B(n36799), .Y(n20481) );
  XOR2XL U39922 ( .A(n42314), .B(n36886), .Y(n24705) );
  XOR2XL U39923 ( .A(n42055), .B(n36892), .Y(n24701) );
  XOR2XL U39924 ( .A(n42315), .B(n42661), .Y(n24697) );
  XOR2XL U39925 ( .A(n42056), .B(n42608), .Y(n24693) );
  XOR2XL U39926 ( .A(n42313), .B(n36888), .Y(n26589) );
  XOR2XL U39927 ( .A(n42054), .B(n36900), .Y(n26585) );
  XOR2XL U39928 ( .A(n42314), .B(n42663), .Y(n26581) );
  XOR2XL U39929 ( .A(n42055), .B(n42607), .Y(n26577) );
  XOR2XL U39930 ( .A(n42053), .B(n42522), .Y(n26597) );
  XOR2XL U39931 ( .A(n42054), .B(n42522), .Y(n26627) );
  XOR2XL U39932 ( .A(n42055), .B(n42522), .Y(n26537) );
  XOR2XL U39933 ( .A(n42052), .B(n42522), .Y(n26417) );
  XNOR2XL U39934 ( .A(n51057), .B(n36717), .Y(n21796) );
  XNOR2XL U39935 ( .A(n51058), .B(n36721), .Y(n21807) );
  XNOR2XL U39936 ( .A(n51056), .B(n36722), .Y(n21785) );
  XNOR2XL U39937 ( .A(n51055), .B(n36714), .Y(n21775) );
  XNOR2XL U39938 ( .A(n51036), .B(n36717), .Y(n20945) );
  XNOR2XL U39939 ( .A(n51035), .B(n36722), .Y(n20935) );
  XNOR2XL U39940 ( .A(n51026), .B(n36716), .Y(n20051) );
  XNOR2XL U39941 ( .A(n51025), .B(n36720), .Y(n20041) );
  XNOR2XL U39942 ( .A(n51014), .B(n41329), .Y(n23672) );
  XNOR2XL U39943 ( .A(n51013), .B(n41332), .Y(n23682) );
  XNOR2XL U39944 ( .A(n51021), .B(n41327), .Y(n23348) );
  XNOR2XL U39945 ( .A(n51022), .B(n41330), .Y(n23358) );
  XNOR2XL U39946 ( .A(n51030), .B(n36716), .Y(n20798) );
  XNOR2XL U39947 ( .A(n51015), .B(n41333), .Y(n23642) );
  XNOR2XL U39948 ( .A(n51042), .B(n36721), .Y(n20955) );
  XNOR2XL U39949 ( .A(n51024), .B(n36720), .Y(n20031) );
  XNOR2XL U39950 ( .A(n51024), .B(n41327), .Y(n23337) );
  XNOR2XL U39951 ( .A(n51014), .B(n36715), .Y(n20492) );
  XNOR2XL U39952 ( .A(n51023), .B(n36715), .Y(n20021) );
  XNOR2XL U39953 ( .A(n51021), .B(n36714), .Y(n20071) );
  XNOR2XL U39954 ( .A(n51022), .B(n36716), .Y(n20061) );
  XNOR2XL U39955 ( .A(n51019), .B(n36714), .Y(n20081) );
  XNOR2XL U39956 ( .A(n51020), .B(n36715), .Y(n20091) );
  XNOR2XL U39957 ( .A(n51012), .B(n41328), .Y(n23662) );
  XNOR2XL U39958 ( .A(n51011), .B(n41327), .Y(n23652) );
  XNOR2XL U39959 ( .A(n50629), .B(n42462), .Y(n21797) );
  XNOR2XL U39960 ( .A(n50630), .B(n42462), .Y(n21808) );
  XNOR2XL U39961 ( .A(n50628), .B(n42462), .Y(n21786) );
  XNOR2XL U39962 ( .A(n50627), .B(n42462), .Y(n21776) );
  XNOR2XL U39963 ( .A(n50608), .B(n42459), .Y(n20946) );
  XNOR2XL U39964 ( .A(n50607), .B(n42460), .Y(n20936) );
  XNOR2XL U39965 ( .A(n50598), .B(n42468), .Y(n20052) );
  XNOR2XL U39966 ( .A(n50597), .B(n42467), .Y(n20042) );
  XNOR2XL U39967 ( .A(n50586), .B(n36860), .Y(n23673) );
  XNOR2XL U39968 ( .A(n50585), .B(n36857), .Y(n23683) );
  XNOR2XL U39969 ( .A(n50593), .B(n36851), .Y(n23349) );
  XNOR2XL U39970 ( .A(n50594), .B(n36859), .Y(n23359) );
  XNOR2XL U39971 ( .A(n50602), .B(n42459), .Y(n20799) );
  XNOR2XL U39972 ( .A(n50587), .B(n36850), .Y(n23643) );
  XNOR2XL U39973 ( .A(n50614), .B(n42459), .Y(n20956) );
  XNOR2XL U39974 ( .A(n50596), .B(n42467), .Y(n20032) );
  XNOR2XL U39975 ( .A(n50596), .B(n36851), .Y(n23338) );
  XNOR2XL U39976 ( .A(n50592), .B(n36858), .Y(n23328) );
  XNOR2XL U39977 ( .A(n50586), .B(n42467), .Y(n20493) );
  XNOR2XL U39978 ( .A(n50595), .B(n42467), .Y(n20022) );
  XNOR2XL U39979 ( .A(n50593), .B(n42468), .Y(n20072) );
  XNOR2XL U39980 ( .A(n50594), .B(n42468), .Y(n20062) );
  XNOR2XL U39981 ( .A(n50591), .B(n42468), .Y(n20082) );
  XNOR2XL U39982 ( .A(n50592), .B(n42468), .Y(n20092) );
  XNOR2XL U39983 ( .A(n50584), .B(n36858), .Y(n23663) );
  XNOR2XL U39984 ( .A(n50583), .B(n36852), .Y(n23653) );
  XNOR2XL U39985 ( .A(n50798), .B(net219308), .Y(n24698) );
  XNOR2XL U39986 ( .A(n50165), .B(n42672), .Y(n24694) );
  XNOR2XL U39987 ( .A(n50797), .B(n36868), .Y(n24690) );
  XNOR2XL U39988 ( .A(n50799), .B(net219310), .Y(n26582) );
  XNOR2XL U39989 ( .A(n50166), .B(n42676), .Y(n26578) );
  XNOR2XL U39990 ( .A(n50798), .B(n41647), .Y(n26574) );
  XNOR2XL U39991 ( .A(n50843), .B(n36791), .Y(n21795) );
  XNOR2XL U39992 ( .A(n50844), .B(n36795), .Y(n21806) );
  XNOR2XL U39993 ( .A(n50842), .B(n36796), .Y(n21784) );
  XNOR2XL U39994 ( .A(n50841), .B(n36792), .Y(n21774) );
  XNOR2XL U39995 ( .A(n50822), .B(n36796), .Y(n20944) );
  XNOR2XL U39996 ( .A(n50821), .B(n36799), .Y(n20934) );
  XNOR2XL U39997 ( .A(n50812), .B(n36797), .Y(n20050) );
  XNOR2XL U39998 ( .A(n50811), .B(n36795), .Y(n20040) );
  XNOR2XL U39999 ( .A(n50800), .B(n41293), .Y(n23671) );
  XNOR2XL U40000 ( .A(n50799), .B(n41295), .Y(n23681) );
  XNOR2XL U40001 ( .A(n50807), .B(n41292), .Y(n23347) );
  XNOR2XL U40002 ( .A(n50808), .B(n41294), .Y(n23357) );
  XNOR2XL U40003 ( .A(n50816), .B(n36791), .Y(n20797) );
  XNOR2XL U40004 ( .A(n50801), .B(n41296), .Y(n23641) );
  XNOR2XL U40005 ( .A(n50828), .B(n36798), .Y(n20954) );
  XNOR2XL U40006 ( .A(n50810), .B(n36799), .Y(n20030) );
  XNOR2XL U40007 ( .A(n50810), .B(n41291), .Y(n23336) );
  XNOR2XL U40008 ( .A(n50800), .B(n36790), .Y(n20491) );
  XNOR2XL U40009 ( .A(n50809), .B(n36793), .Y(n20020) );
  XNOR2XL U40010 ( .A(n50807), .B(n36798), .Y(n20070) );
  XNOR2XL U40011 ( .A(n50808), .B(n36790), .Y(n20060) );
  XNOR2XL U40012 ( .A(n50805), .B(n36796), .Y(n20080) );
  XNOR2XL U40013 ( .A(n50806), .B(n36790), .Y(n20090) );
  XNOR2XL U40014 ( .A(n50798), .B(n41290), .Y(n23661) );
  XNOR2XL U40015 ( .A(n50797), .B(n41291), .Y(n23651) );
  XNOR2XL U40016 ( .A(n51014), .B(n42552), .Y(n26595) );
  XNOR2XL U40017 ( .A(n50584), .B(net219468), .Y(n24700) );
  XNOR2XL U40018 ( .A(n51225), .B(n36867), .Y(n24696) );
  XNOR2XL U40019 ( .A(n50583), .B(n42586), .Y(n24692) );
  XNOR2XL U40020 ( .A(n50585), .B(net219434), .Y(n26584) );
  XNOR2XL U40021 ( .A(n51226), .B(n36867), .Y(n26580) );
  XNOR2XL U40022 ( .A(n50584), .B(n36865), .Y(n26576) );
  XNOR2XL U40023 ( .A(n51228), .B(n36867), .Y(n26640) );
  XNOR2XL U40024 ( .A(n51013), .B(n42552), .Y(n26625) );
  XNOR2XL U40025 ( .A(n51012), .B(n42552), .Y(n26535) );
  XNOR2XL U40026 ( .A(n50586), .B(n42505), .Y(n26596) );
  XNOR2XL U40027 ( .A(n51014), .B(n41282), .Y(n26553) );
  XNOR2XL U40028 ( .A(n51012), .B(n41283), .Y(n24699) );
  XNOR2XL U40029 ( .A(n50380), .B(n36905), .Y(n24695) );
  XNOR2XL U40030 ( .A(n51011), .B(n42633), .Y(n24691) );
  XNOR2XL U40031 ( .A(n51013), .B(n41281), .Y(n26583) );
  XNOR2XL U40032 ( .A(n50381), .B(n36905), .Y(n26579) );
  XNOR2XL U40033 ( .A(n51012), .B(n42630), .Y(n26575) );
  XNOR2XL U40034 ( .A(n50585), .B(n42505), .Y(n26626) );
  XOR2XL U40035 ( .A(n42311), .B(n42493), .Y(n20443) );
  XOR2XL U40036 ( .A(n42309), .B(n42493), .Y(n20464) );
  XOR2XL U40037 ( .A(n42310), .B(n42493), .Y(n20453) );
  XOR2XL U40038 ( .A(n42313), .B(n42493), .Y(n20505) );
  XOR2XL U40039 ( .A(n42315), .B(n42493), .Y(n20433) );
  XOR2XL U40040 ( .A(n42308), .B(n42493), .Y(n20475) );
  XOR2XL U40041 ( .A(n42314), .B(n42493), .Y(n20485) );
  XOR2XL U40042 ( .A(n42269), .B(n42487), .Y(n21799) );
  XOR2XL U40043 ( .A(n42268), .B(n42487), .Y(n21810) );
  XOR2XL U40044 ( .A(n42270), .B(n42487), .Y(n21788) );
  XOR2XL U40045 ( .A(n42271), .B(n42487), .Y(n21778) );
  XOR2XL U40046 ( .A(n42290), .B(n42483), .Y(n20948) );
  XOR2XL U40047 ( .A(n42291), .B(n42484), .Y(n20938) );
  XOR2XL U40048 ( .A(n42300), .B(n42492), .Y(n20054) );
  XOR2XL U40049 ( .A(n42301), .B(n42491), .Y(n20044) );
  XOR2XL U40050 ( .A(n42312), .B(n36811), .Y(n23675) );
  XOR2XL U40051 ( .A(n42313), .B(n36813), .Y(n23685) );
  XOR2XL U40052 ( .A(n42305), .B(n36814), .Y(n23351) );
  XOR2XL U40053 ( .A(n42304), .B(n36810), .Y(n23361) );
  XOR2XL U40054 ( .A(n42296), .B(n42486), .Y(n20801) );
  XOR2XL U40055 ( .A(n42311), .B(n36813), .Y(n23645) );
  XOR2XL U40056 ( .A(n42284), .B(n42483), .Y(n20958) );
  XOR2XL U40057 ( .A(n42302), .B(n42491), .Y(n20034) );
  XOR2XL U40058 ( .A(n42302), .B(n36807), .Y(n23340) );
  XOR2XL U40059 ( .A(n42306), .B(n36817), .Y(n23330) );
  XOR2XL U40060 ( .A(n42312), .B(n42491), .Y(n20495) );
  XOR2XL U40061 ( .A(n42303), .B(n42491), .Y(n20024) );
  XOR2XL U40062 ( .A(n42305), .B(n42492), .Y(n20074) );
  XOR2XL U40063 ( .A(n42304), .B(n42492), .Y(n20064) );
  XOR2XL U40064 ( .A(n42307), .B(n42492), .Y(n20084) );
  XOR2XL U40065 ( .A(n42306), .B(n42492), .Y(n20094) );
  XOR2XL U40066 ( .A(n42314), .B(n36809), .Y(n23665) );
  XOR2XL U40067 ( .A(n42315), .B(n36815), .Y(n23655) );
  XNOR2XL U40068 ( .A(n50800), .B(n42540), .Y(n26594) );
  XNOR2XL U40069 ( .A(n50799), .B(n42540), .Y(n26624) );
  XNOR2XL U40070 ( .A(n50427), .B(n36767), .Y(n21811) );
  XNOR2XL U40071 ( .A(n51270), .B(n36746), .Y(n21790) );
  XNOR2XL U40072 ( .A(n51269), .B(n36740), .Y(n21779) );
  XNOR2XL U40073 ( .A(n50418), .B(n36773), .Y(n21913) );
  XNOR2XL U40074 ( .A(n50419), .B(n36766), .Y(n21831) );
  XNOR2XL U40075 ( .A(n50412), .B(n36785), .Y(n24315) );
  XNOR2XL U40076 ( .A(n50421), .B(n36772), .Y(n21851) );
  XNOR2XL U40077 ( .A(n50412), .B(n36773), .Y(n21882) );
  XNOR2XL U40078 ( .A(n51250), .B(n36743), .Y(n20949) );
  XNOR2XL U40079 ( .A(n51249), .B(n36747), .Y(n20939) );
  XNOR2XL U40080 ( .A(n50395), .B(n36765), .Y(n20055) );
  XNOR2XL U40081 ( .A(n51239), .B(n36749), .Y(n20045) );
  XNOR2XL U40082 ( .A(n50387), .B(n36779), .Y(n23636) );
  XNOR2XL U40083 ( .A(n50383), .B(n36784), .Y(n23676) );
  XNOR2XL U40084 ( .A(n50382), .B(n36782), .Y(n23686) );
  XNOR2XL U40085 ( .A(n50396), .B(n36778), .Y(n24507) );
  XNOR2XL U40086 ( .A(n51229), .B(n36750), .Y(n20444) );
  XNOR2XL U40087 ( .A(n50397), .B(n36778), .Y(n24517) );
  XNOR2XL U40088 ( .A(n50390), .B(n36776), .Y(n23352) );
  XNOR2XL U40089 ( .A(n51236), .B(n41302), .Y(n23362) );
  XNOR2XL U40090 ( .A(n50397), .B(n36764), .Y(n20834) );
  XNOR2XL U40091 ( .A(n51230), .B(n36744), .Y(n20455) );
  XNOR2XL U40092 ( .A(n50396), .B(n36766), .Y(n20823) );
  XNOR2XL U40093 ( .A(n50384), .B(n36784), .Y(n23646) );
  XNOR2XL U40094 ( .A(n50411), .B(n36768), .Y(n20959) );
  XNOR2XL U40095 ( .A(n51238), .B(n36748), .Y(n20035) );
  XNOR2XL U40096 ( .A(n51238), .B(n41304), .Y(n23342) );
  XNOR2XL U40097 ( .A(n50389), .B(n36783), .Y(n23331) );
  XNOR2XL U40098 ( .A(n51237), .B(n36741), .Y(n20025) );
  XNOR2XL U40099 ( .A(n51235), .B(n36748), .Y(n20075) );
  XNOR2XL U40100 ( .A(n50380), .B(n36765), .Y(n20434) );
  XNOR2XL U40101 ( .A(n51236), .B(n36747), .Y(n20065) );
  XNOR2XL U40102 ( .A(n50388), .B(n36770), .Y(n20085) );
  XNOR2XL U40103 ( .A(n50389), .B(n36774), .Y(n20095) );
  XNOR2XL U40104 ( .A(n50387), .B(n36774), .Y(n20476) );
  XNOR2XL U40105 ( .A(n50381), .B(n36771), .Y(n20486) );
  XNOR2XL U40106 ( .A(n50381), .B(n36780), .Y(n23666) );
  XNOR2XL U40107 ( .A(n50380), .B(n36777), .Y(n23656) );
  XNOR2XL U40108 ( .A(n50166), .B(n42708), .Y(n24702) );
  XNOR2XL U40109 ( .A(n50381), .B(n41287), .Y(n24703) );
  XNOR2XL U40110 ( .A(n51226), .B(n36871), .Y(n24704) );
  XNOR2XL U40111 ( .A(n50167), .B(n42706), .Y(n26586) );
  XNOR2XL U40112 ( .A(n50382), .B(n34435), .Y(n26587) );
  XNOR2XL U40113 ( .A(n51227), .B(n42696), .Y(n26588) );
  XNOR2XL U40114 ( .A(n50383), .B(n42576), .Y(n26599) );
  XNOR2XL U40115 ( .A(n50382), .B(n42576), .Y(n26629) );
  XOR2XL U40116 ( .A(n42312), .B(n36801), .Y(n26598) );
  XOR2XL U40117 ( .A(n42313), .B(n36873), .Y(n26628) );
  XOR2XL U40118 ( .A(n42314), .B(n36801), .Y(n26538) );
  XOR2XL U40119 ( .A(n42311), .B(n36877), .Y(n26418) );
  NAND3XL U40120 ( .A(n10503), .B(n10502), .C(n10498), .Y(n10148) );
  AND4XL U40121 ( .A(n12794), .B(n12736), .C(n10559), .D(n29117), .Y(n10174)
         );
  NOR2BXL U40122 ( .AN(n10565), .B(n10564), .Y(n29117) );
  AND4XL U40123 ( .A(n10548), .B(n12150), .C(n26891), .D(n10608), .Y(n10173)
         );
  AND2XL U40124 ( .A(n10607), .B(n10606), .Y(n26891) );
  NAND3XL U40125 ( .A(net210435), .B(net171222), .C(n10184), .Y(n47812) );
  INVXL U40126 ( .A(n39304), .Y(net210434) );
  NAND4XL U40127 ( .A(n10554), .B(n10555), .C(n10556), .D(n26650), .Y(n10172)
         );
  AND2XL U40128 ( .A(n37349), .B(n10553), .Y(n26650) );
  XOR2XL U40129 ( .A(n42056), .B(n42522), .Y(n26567) );
  XNOR2XL U40130 ( .A(n51011), .B(n42552), .Y(n26565) );
  XNOR2XL U40131 ( .A(n50583), .B(n42504), .Y(n26566) );
  XNOR2XL U40132 ( .A(n50797), .B(n42540), .Y(n26564) );
  XNOR2XL U40133 ( .A(n50380), .B(n42576), .Y(n26569) );
  XOR2XL U40134 ( .A(n42315), .B(n41322), .Y(n26568) );
  INVX1 U40135 ( .A(n41796), .Y(n50145) );
  NAND2X1 U40136 ( .A(n42316), .B(n50134), .Y(n9737) );
  NAND2X1 U40137 ( .A(n19376), .B(n50132), .Y(n19278) );
  NAND2X1 U40138 ( .A(n50147), .B(n50148), .Y(n9702) );
  XNOR2XL U40139 ( .A(n36844), .B(n33994), .Y(net213353) );
  XNOR2XL U40140 ( .A(n36838), .B(n33818), .Y(n46151) );
  NAND4X2 U40141 ( .A(n46176), .B(n46175), .C(n46174), .D(n46173), .Y(n12723)
         );
  NOR4X2 U40142 ( .A(n26688), .B(n26687), .C(n26686), .D(n26685), .Y(n46173)
         );
  XNOR2XL U40143 ( .A(n36733), .B(n33570), .Y(n46923) );
  NAND4X2 U40144 ( .A(n44439), .B(n44438), .C(n44437), .D(n44436), .Y(n12708)
         );
  NOR4X2 U40145 ( .A(n25155), .B(n25154), .C(n25153), .D(n25152), .Y(n44436)
         );
  XNOR2XL U40146 ( .A(n36735), .B(n33954), .Y(net211489) );
  NAND4X2 U40147 ( .A(n47173), .B(n47172), .C(n47171), .D(n47170), .Y(n11399)
         );
  XNOR2XL U40148 ( .A(n36733), .B(n33698), .Y(n47172) );
  XNOR2XL U40149 ( .A(n36846), .B(n34114), .Y(n46208) );
  NOR2X2 U40150 ( .A(n23809), .B(n23808), .Y(n46197) );
  XNOR2XL U40151 ( .A(n36843), .B(n33714), .Y(n45636) );
  XNOR2XL U40152 ( .A(n36736), .B(n33946), .Y(net211479) );
  NOR2X2 U40153 ( .A(n23819), .B(n23818), .Y(n46181) );
  XNOR2XL U40154 ( .A(n36838), .B(n33914), .Y(n46101) );
  XNOR2XL U40155 ( .A(n36838), .B(n33610), .Y(n45725) );
  XNOR2XL U40156 ( .A(n42508), .B(n34120), .Y(n43884) );
  NAND4X2 U40157 ( .A(n47267), .B(n47266), .C(n47265), .D(n47264), .Y(n13015)
         );
  XNOR2XL U40158 ( .A(n34082), .B(n42569), .Y(n43823) );
  XNOR2XL U40159 ( .A(n34010), .B(n42561), .Y(n44196) );
  NAND4X2 U40160 ( .A(n44286), .B(n44285), .C(n44284), .D(n44283), .Y(n12062)
         );
  XNOR2XL U40161 ( .A(n34128), .B(n42504), .Y(n43915) );
  XNOR2XL U40162 ( .A(n34090), .B(n42569), .Y(n43832) );
  XNOR2XL U40163 ( .A(n42472), .B(n34256), .Y(n47433) );
  XNOR2XL U40164 ( .A(n33978), .B(n42561), .Y(n44220) );
  XNOR2XL U40165 ( .A(n42472), .B(n34232), .Y(n47466) );
  NAND4X2 U40166 ( .A(n45704), .B(n45703), .C(n45702), .D(n45701), .Y(
        net209253) );
  XNOR2XL U40167 ( .A(n36841), .B(n33970), .Y(n45703) );
  XNOR2XL U40168 ( .A(n36850), .B(n34144), .Y(n46280) );
  NAND4X2 U40169 ( .A(n43978), .B(n43977), .C(n43976), .D(n43975), .Y(n48185)
         );
  XNOR2XL U40170 ( .A(n34152), .B(n42504), .Y(n43977) );
  XNOR2XL U40171 ( .A(n42472), .B(n34192), .Y(n47477) );
  XNOR2XL U40172 ( .A(n42508), .B(n34144), .Y(n44008) );
  XNOR2XL U40173 ( .A(n42472), .B(n34216), .Y(n47400) );
  XNOR2XL U40174 ( .A(n36856), .B(n34168), .Y(n46269) );
  XNOR2XL U40175 ( .A(n34224), .B(n42504), .Y(n44702) );
  XNOR2XL U40176 ( .A(n34176), .B(n42504), .Y(n44100) );
  XNOR2XL U40177 ( .A(n34106), .B(n42569), .Y(n43853) );
  NAND4X2 U40178 ( .A(n44763), .B(n44762), .C(n44761), .D(n44760), .Y(n48173)
         );
  XNOR2XL U40179 ( .A(n34208), .B(n42502), .Y(n44762) );
  XNOR2XL U40180 ( .A(n33586), .B(n41630), .Y(n44506) );
  XNOR2XL U40181 ( .A(n42471), .B(n34368), .Y(n47610) );
  XNOR2XL U40182 ( .A(n34160), .B(n42504), .Y(n43946) );
  XNOR2XL U40183 ( .A(n33994), .B(n42561), .Y(n44205) );
  XNOR2XL U40184 ( .A(n33898), .B(n42568), .Y(n43642) );
  XNOR2XL U40185 ( .A(n36854), .B(n34128), .Y(n46219) );
  XNOR2XL U40186 ( .A(n36734), .B(n33714), .Y(n47885) );
  XNOR2XL U40187 ( .A(n36768), .B(n34113), .Y(n47565) );
  XNOR2XL U40188 ( .A(n42472), .B(n34152), .Y(n47519) );
  XOR2XL U40189 ( .A(n34380), .B(n36871), .Y(n44958) );
  XOR2XL U40190 ( .A(n34384), .B(net219434), .Y(n44954) );
  XOR2XL U40191 ( .A(n34369), .B(n42680), .Y(n44953) );
  XOR2XL U40192 ( .A(n34370), .B(n42670), .Y(n44952) );
  XOR2XL U40193 ( .A(n34396), .B(n36827), .Y(n45062) );
  XNOR2XL U40194 ( .A(n36847), .B(n33906), .Y(n46106) );
  XNOR2XL U40195 ( .A(n36840), .B(n34026), .Y(net213363) );
  XNOR2XL U40196 ( .A(n36736), .B(n33938), .Y(net211474) );
  NOR4X2 U40197 ( .A(n20104), .B(n20103), .C(n20102), .D(n20101), .Y(net211476) );
  XOR2XL U40198 ( .A(n34308), .B(n42693), .Y(n45504) );
  XNOR2XL U40199 ( .A(n36852), .B(n34264), .Y(net212475) );
  XOR2XL U40200 ( .A(n34332), .B(n36871), .Y(n45429) );
  XOR2XL U40201 ( .A(n34340), .B(n42700), .Y(n45180) );
  XOR2XL U40202 ( .A(n34244), .B(n36871), .Y(n44838) );
  XOR2XL U40203 ( .A(n34260), .B(n36871), .Y(n44807) );
  XOR2XL U40204 ( .A(n34284), .B(n41385), .Y(n45301) );
  XOR2XL U40205 ( .A(n34300), .B(n42690), .Y(n45390) );
  XOR2XL U40206 ( .A(n34268), .B(n41385), .Y(n44865) );
  XOR2XL U40207 ( .A(n34276), .B(n36871), .Y(n45332) );
  XOR2XL U40208 ( .A(n34392), .B(net219434), .Y(n44918) );
  XNOR2XL U40209 ( .A(n42471), .B(n34144), .Y(n47541) );
  XOR2XL U40210 ( .A(n34382), .B(n36868), .Y(n44912) );
  XOR2XL U40211 ( .A(n34374), .B(net219330), .Y(n44975) );
  XOR2XL U40212 ( .A(n34381), .B(n42628), .Y(n44913) );
  XOR2XL U40213 ( .A(n34365), .B(n42624), .Y(n44968) );
  XOR2XL U40214 ( .A(n36768), .B(n34393), .Y(n47704) );
  NAND4X2 U40215 ( .A(n47262), .B(n47261), .C(n47260), .D(n47259), .Y(n12960)
         );
  XNOR2XL U40216 ( .A(n36734), .B(n33898), .Y(n47261) );
  NOR2X2 U40217 ( .A(n19548), .B(n19547), .Y(n47260) );
  XOR2XL U40218 ( .A(n36717), .B(n34405), .Y(n47676) );
  XNOR2XL U40219 ( .A(n42472), .B(n34184), .Y(n47488) );
  NAND4X2 U40220 ( .A(n47183), .B(n47182), .C(n47181), .D(n47180), .Y(n11398)
         );
  XNOR2XL U40221 ( .A(n42471), .B(n34328), .Y(n47588) );
  XNOR2XL U40222 ( .A(n42472), .B(n34224), .Y(n47389) );
  XNOR2XL U40223 ( .A(n42472), .B(n34240), .Y(n47455) );
  XNOR2XL U40224 ( .A(n36735), .B(n34090), .Y(n47289) );
  XNOR2XL U40225 ( .A(n42472), .B(n34200), .Y(n47422) );
  XNOR2XL U40226 ( .A(n33610), .B(n42559), .Y(n44532) );
  XOR2XL U40227 ( .A(n41290), .B(n34390), .Y(n46583) );
  XNOR2XL U40228 ( .A(n42472), .B(n34272), .Y(n47378) );
  XNOR2XL U40229 ( .A(n42471), .B(n34160), .Y(n47530) );
  XNOR2XL U40230 ( .A(n42472), .B(n34208), .Y(n47411) );
  XOR2XL U40231 ( .A(n34373), .B(n42631), .Y(n44949) );
  XOR2XL U40232 ( .A(n34237), .B(n42629), .Y(n44829) );
  XOR2XL U40233 ( .A(n34253), .B(n42627), .Y(n44798) );
  XOR2XL U40234 ( .A(n34221), .B(n34447), .Y(n44645) );
  XOR2XL U40235 ( .A(n34213), .B(n42631), .Y(n44736) );
  XOR2XL U40236 ( .A(n34245), .B(n42626), .Y(n44767) );
  XOR2XL U40237 ( .A(n34422), .B(n36868), .Y(n45028) );
  XOR2XL U40238 ( .A(n34218), .B(n42560), .Y(n44699) );
  XOR2XL U40239 ( .A(n34178), .B(n42560), .Y(n44128) );
  XOR2XL U40240 ( .A(n34325), .B(n42631), .Y(n45420) );
  XOR2XL U40241 ( .A(n34333), .B(n42626), .Y(n45171) );
  XOR2XL U40242 ( .A(n34329), .B(n41319), .Y(n45175) );
  XOR2XL U40243 ( .A(n34285), .B(n42629), .Y(n45350) );
  XOR2XL U40244 ( .A(n34277), .B(n42629), .Y(n45292) );
  XOR2XL U40245 ( .A(n34313), .B(n41319), .Y(n45444) );
  XOR2XL U40246 ( .A(n34293), .B(n41282), .Y(n45358) );
  XOR2XL U40247 ( .A(n34233), .B(n42684), .Y(n44833) );
  XOR2XL U40248 ( .A(n34245), .B(n41282), .Y(n44837) );
  XOR2XL U40249 ( .A(n34249), .B(n41379), .Y(n44802) );
  XOR2XL U40250 ( .A(n34261), .B(n41283), .Y(n44806) );
  XOR2XL U40251 ( .A(n34237), .B(n41281), .Y(n44684) );
  XOR2XL U40252 ( .A(n34221), .B(n41281), .Y(n44744) );
  XOR2XL U40253 ( .A(n34209), .B(n41379), .Y(n44740) );
  XNOR2XL U40254 ( .A(n36776), .B(n34385), .Y(n46580) );
  XOR2XL U40255 ( .A(n34149), .B(n41282), .Y(n44021) );
  XOR2XL U40256 ( .A(n34181), .B(n41281), .Y(n44051) );
  XOR2XL U40257 ( .A(n34173), .B(n41281), .Y(n43928) );
  XOR2XL U40258 ( .A(n34229), .B(n41281), .Y(n44653) );
  XOR2XL U40259 ( .A(n34165), .B(n41282), .Y(n43959) );
  XOR2XL U40260 ( .A(n34173), .B(n42632), .Y(n44043) );
  XOR2XL U40261 ( .A(n34189), .B(n42628), .Y(n44105) );
  XOR2XL U40262 ( .A(n34169), .B(n36905), .Y(n44047) );
  XOR2XL U40263 ( .A(n34165), .B(n42633), .Y(n43920) );
  XOR2XL U40264 ( .A(n34185), .B(n36903), .Y(n44109) );
  XOR2XL U40265 ( .A(n34229), .B(n34447), .Y(n44676) );
  XOR2XL U40266 ( .A(n34157), .B(n42628), .Y(n43951) );
  XOR2XL U40267 ( .A(n34161), .B(n36905), .Y(n43924) );
  XOR2XL U40268 ( .A(n34225), .B(n36905), .Y(n44680) );
  XOR2XL U40269 ( .A(n34181), .B(n42626), .Y(n44074) );
  XOR2XL U40270 ( .A(n34153), .B(n36903), .Y(n43955) );
  XOR2XL U40271 ( .A(n34125), .B(n42630), .Y(n43858) );
  XOR2XL U40272 ( .A(n34205), .B(n34447), .Y(n44707) );
  XOR2XL U40273 ( .A(n36813), .B(n34419), .Y(n46602) );
  XOR2XL U40274 ( .A(n34426), .B(n42706), .Y(n45029) );
  XOR2XL U40275 ( .A(n34322), .B(n42669), .Y(n45423) );
  XOR2XL U40276 ( .A(n34330), .B(n42672), .Y(n45174) );
  XOR2XL U40277 ( .A(n34338), .B(n42669), .Y(n45203) );
  XOR2XL U40278 ( .A(n34314), .B(n34444), .Y(n45443) );
  XOR2XL U40279 ( .A(n34282), .B(n42672), .Y(n45353) );
  XOR2XL U40280 ( .A(n34274), .B(n42669), .Y(n45295) );
  XOR2XL U40281 ( .A(n34254), .B(n36868), .Y(n44797) );
  XNOR2XL U40282 ( .A(n42471), .B(n34320), .Y(n47302) );
  XOR2XL U40283 ( .A(n34212), .B(n42696), .Y(n44716) );
  XOR2XL U40284 ( .A(n34180), .B(n42696), .Y(n44052) );
  XOR2XL U40285 ( .A(n34252), .B(n42696), .Y(n44776) );
  XOR2XL U40286 ( .A(n33658), .B(n42560), .Y(n44448) );
  XNOR2XL U40287 ( .A(n41329), .B(n34389), .Y(n46578) );
  XOR2XL U40288 ( .A(n34334), .B(n42615), .Y(n45170) );
  XOR2XL U40289 ( .A(n34342), .B(net219330), .Y(n45178) );
  XOR2XL U40290 ( .A(n34342), .B(n36868), .Y(n45199) );
  XOR2XL U40291 ( .A(n34318), .B(n36868), .Y(n45439) );
  XOR2XL U40292 ( .A(n34286), .B(n42615), .Y(n45349) );
  XOR2XL U40293 ( .A(n34278), .B(n36868), .Y(n45291) );
  XOR2XL U40294 ( .A(n34294), .B(n42615), .Y(n45380) );
  XOR2XL U40295 ( .A(n34286), .B(net219330), .Y(n45299) );
  XOR2XL U40296 ( .A(n34302), .B(n42615), .Y(n45494) );
  XOR2XL U40297 ( .A(n34234), .B(n42671), .Y(n44832) );
  XOR2XL U40298 ( .A(n34246), .B(n36870), .Y(n44836) );
  XOR2XL U40299 ( .A(n34250), .B(n42672), .Y(n44801) );
  XOR2XL U40300 ( .A(n34150), .B(net219336), .Y(n44020) );
  XOR2XL U40301 ( .A(n34230), .B(net219330), .Y(n44652) );
  XOR2XL U40302 ( .A(n34174), .B(n41284), .Y(n44042) );
  XOR2XL U40303 ( .A(n34190), .B(n41284), .Y(n44104) );
  XOR2XL U40304 ( .A(n34138), .B(n42671), .Y(n44016) );
  XOR2XL U40305 ( .A(n34170), .B(n42671), .Y(n44046) );
  XOR2XL U40306 ( .A(n34222), .B(n42614), .Y(n44644) );
  XOR2XL U40307 ( .A(n34166), .B(n41284), .Y(n43919) );
  XOR2XL U40308 ( .A(n34186), .B(n36907), .Y(n44108) );
  XOR2XL U40309 ( .A(n34158), .B(n42619), .Y(n43950) );
  XOR2XL U40310 ( .A(n34162), .B(n42671), .Y(n43923) );
  XOR2XL U40311 ( .A(n34218), .B(n42672), .Y(n44648) );
  XOR2XL U40312 ( .A(n34226), .B(n42672), .Y(n44679) );
  XOR2XL U40313 ( .A(n34182), .B(n42620), .Y(n44073) );
  XOR2XL U40314 ( .A(n34154), .B(n42671), .Y(n43954) );
  XOR2XL U40315 ( .A(n34206), .B(n42616), .Y(n44706) );
  XOR2XL U40316 ( .A(n34148), .B(n42698), .Y(n44022) );
  XOR2XL U40317 ( .A(n34196), .B(n42698), .Y(n44114) );
  XOR2XL U40318 ( .A(n34172), .B(n42697), .Y(n43929) );
  XOR2XL U40319 ( .A(n34236), .B(n42698), .Y(n44685) );
  XOR2XL U40320 ( .A(n34164), .B(n42697), .Y(n43960) );
  XOR2XL U40321 ( .A(n34140), .B(n42698), .Y(n43898) );
  XOR2XL U40322 ( .A(n34188), .B(n42698), .Y(n44083) );
  XNOR2XL U40323 ( .A(n42472), .B(n34264), .Y(n47367) );
  XOR2XL U40324 ( .A(n41314), .B(n34423), .Y(n46597) );
  XOR2XL U40325 ( .A(n34236), .B(n42637), .Y(n44830) );
  XOR2XL U40326 ( .A(n34252), .B(n42637), .Y(n44799) );
  XOR2XL U40327 ( .A(n34220), .B(n42637), .Y(n44646) );
  XOR2XL U40328 ( .A(n34212), .B(n42637), .Y(n44737) );
  XOR2XL U40329 ( .A(n34244), .B(n42637), .Y(n44768) );
  XOR2XL U40330 ( .A(n34264), .B(net219434), .Y(n44803) );
  XOR2XL U40331 ( .A(n34336), .B(net219468), .Y(n45425) );
  XOR2XL U40332 ( .A(n34344), .B(net219468), .Y(n45176) );
  XOR2XL U40333 ( .A(n34248), .B(net219434), .Y(n44834) );
  XOR2XL U40334 ( .A(n34296), .B(net219434), .Y(n45355) );
  XOR2XL U40335 ( .A(n34328), .B(n42592), .Y(n45417) );
  XOR2XL U40336 ( .A(n34288), .B(net219468), .Y(n45297) );
  XOR2XL U40337 ( .A(n34336), .B(n34450), .Y(n45168) );
  XOR2XL U40338 ( .A(n34332), .B(n42638), .Y(n45172) );
  XOR2XL U40339 ( .A(n34312), .B(net219434), .Y(n45500) );
  XOR2XL U40340 ( .A(n34240), .B(n42592), .Y(n44826) );
  XOR2XL U40341 ( .A(n34288), .B(n42592), .Y(n45347) );
  XOR2XL U40342 ( .A(n34284), .B(n42638), .Y(n45351) );
  XOR2XL U40343 ( .A(n34272), .B(net219434), .Y(n44861) );
  XOR2XL U40344 ( .A(n34280), .B(net219468), .Y(n45328) );
  XOR2XL U40345 ( .A(n34280), .B(n42592), .Y(n45289) );
  XOR2XL U40346 ( .A(n34276), .B(n42638), .Y(n45293) );
  XOR2XL U40347 ( .A(n34240), .B(net219434), .Y(n44681) );
  XOR2XL U40348 ( .A(n34224), .B(net219434), .Y(n44741) );
  XOR2XL U40349 ( .A(n34256), .B(net219434), .Y(n44772) );
  XOR2XL U40350 ( .A(n34256), .B(n42592), .Y(n44795) );
  XOR2XL U40351 ( .A(n34224), .B(n42592), .Y(n44642) );
  XOR2XL U40352 ( .A(n34216), .B(n42592), .Y(n44733) );
  XOR2XL U40353 ( .A(n34152), .B(net219494), .Y(n44018) );
  XOR2XL U40354 ( .A(n34232), .B(net219468), .Y(n44650) );
  XOR2XL U40355 ( .A(n34192), .B(net219460), .Y(n44079) );
  XOR2XL U40356 ( .A(n34216), .B(net219468), .Y(n44712) );
  XOR2XL U40357 ( .A(n34172), .B(n42637), .Y(n44044) );
  XOR2XL U40358 ( .A(n34188), .B(n42637), .Y(n44106) );
  XOR2XL U40359 ( .A(n34144), .B(n34450), .Y(n44010) );
  XOR2XL U40360 ( .A(n34176), .B(n34450), .Y(n44040) );
  XOR2XL U40361 ( .A(n34164), .B(n42637), .Y(n43921) );
  XOR2XL U40362 ( .A(n34192), .B(n34450), .Y(n44102) );
  XOR2XL U40363 ( .A(n34156), .B(n42638), .Y(n43952) );
  XOR2XL U40364 ( .A(n34168), .B(n42586), .Y(n43917) );
  XOR2XL U40365 ( .A(n34160), .B(n36863), .Y(n43948) );
  XOR2XL U40366 ( .A(n34180), .B(n42637), .Y(n44075) );
  XOR2XL U40367 ( .A(n34204), .B(n42638), .Y(n44708) );
  XNOR2XL U40368 ( .A(n36772), .B(n33993), .Y(n47034) );
  XOR2XL U40369 ( .A(n34364), .B(n36821), .Y(n44947) );
  XOR2XL U40370 ( .A(n33660), .B(n36823), .Y(n44449) );
  XOR2XL U40371 ( .A(n33794), .B(n42560), .Y(n44293) );
  XOR2XL U40372 ( .A(n33642), .B(n42560), .Y(n44494) );
  XOR2XL U40373 ( .A(n34332), .B(n36825), .Y(n45222) );
  XOR2XL U40374 ( .A(n34356), .B(n36821), .Y(n44989) );
  XOR2XL U40375 ( .A(n34186), .B(n42559), .Y(n44159) );
  XOR2XL U40376 ( .A(n34354), .B(n42557), .Y(n44990) );
  XOR2XL U40377 ( .A(n34366), .B(n42533), .Y(n44943) );
  XOR2XL U40378 ( .A(n34138), .B(n42558), .Y(n44005) );
  XOR2XL U40379 ( .A(n34162), .B(n42558), .Y(n44066) );
  XOR2XL U40380 ( .A(n34202), .B(n42557), .Y(n44759) );
  XOR2XL U40381 ( .A(n34362), .B(n42557), .Y(n44946) );
  XOR2XL U40382 ( .A(n34314), .B(n41630), .Y(n45411) );
  XOR2XL U40383 ( .A(n36784), .B(n34417), .Y(n46604) );
  XOR2XL U40384 ( .A(n34361), .B(n42575), .Y(n44944) );
  XOR2XL U40385 ( .A(n33644), .B(n36824), .Y(n44495) );
  XOR2XL U40386 ( .A(n36839), .B(n34418), .Y(n46603) );
  XOR2XL U40387 ( .A(n34169), .B(n36709), .Y(n43932) );
  XOR2XL U40388 ( .A(n34170), .B(n42704), .Y(n43931) );
  XOR2XL U40389 ( .A(n42094), .B(n36883), .Y(n43930) );
  XOR2XL U40390 ( .A(n34233), .B(n36875), .Y(n44688) );
  XOR2XL U40391 ( .A(n34234), .B(n42704), .Y(n44687) );
  XOR2XL U40392 ( .A(n42086), .B(n36885), .Y(n44686) );
  XOR2XL U40393 ( .A(n34217), .B(n42718), .Y(n44748) );
  XOR2XL U40394 ( .A(n34218), .B(n42704), .Y(n44747) );
  XOR2XL U40395 ( .A(n34220), .B(n36871), .Y(n44745) );
  XOR2XL U40396 ( .A(n42060), .B(n42722), .Y(n43901) );
  XOR2XL U40397 ( .A(n34138), .B(n41641), .Y(n43900) );
  XOR2XL U40398 ( .A(n42098), .B(n36887), .Y(n43899) );
  XOR2XL U40399 ( .A(n34185), .B(n42717), .Y(n44086) );
  XOR2XL U40400 ( .A(n34186), .B(n42705), .Y(n44085) );
  XOR2XL U40401 ( .A(n42092), .B(n36880), .Y(n44084) );
  XOR2XL U40402 ( .A(n34249), .B(n42718), .Y(n44779) );
  XOR2XL U40403 ( .A(n34250), .B(n42707), .Y(n44778) );
  XOR2XL U40404 ( .A(n42084), .B(n36885), .Y(n44777) );
  XNOR2XL U40405 ( .A(n42473), .B(n34304), .Y(n47323) );
  XNOR2XL U40406 ( .A(n34209), .B(n42717), .Y(n41720) );
  XNOR2XL U40407 ( .A(n34210), .B(n41641), .Y(n41721) );
  NOR4X2 U40408 ( .A(n44461), .B(n44460), .C(n25096), .D(n25095), .Y(n44462)
         );
  XNOR2XL U40409 ( .A(n36858), .B(n34296), .Y(n46341) );
  XOR2XL U40410 ( .A(n34190), .B(n42535), .Y(n44154) );
  XOR2XL U40411 ( .A(n36747), .B(n34396), .Y(n47701) );
  XOR2XL U40412 ( .A(n41303), .B(n34396), .Y(n46591) );
  XNOR2XL U40413 ( .A(n36857), .B(n34376), .Y(n46471) );
  XOR2XL U40414 ( .A(n42470), .B(n34400), .Y(n47698) );
  XNOR2XL U40415 ( .A(n36854), .B(n34392), .Y(n46576) );
  XOR2XL U40416 ( .A(n41305), .B(n34388), .Y(n46582) );
  XOR2XL U40417 ( .A(n34025), .B(n36785), .Y(n45690) );
  NOR2XL U40418 ( .A(n12723), .B(n46177), .Y(net212716) );
  XOR2XL U40419 ( .A(n33769), .B(n36780), .Y(n46177) );
  XOR2XL U40420 ( .A(n41299), .B(n33812), .Y(n46163) );
  NOR2X2 U40421 ( .A(n11722), .B(n44489), .Y(net214879) );
  XOR2XL U40422 ( .A(n33732), .B(n36831), .Y(n44267) );
  XOR2XL U40423 ( .A(n33921), .B(n36782), .Y(n46093) );
  XOR2XL U40424 ( .A(n33521), .B(n36778), .Y(n45818) );
  XOR2XL U40425 ( .A(n41305), .B(n33980), .Y(n45694) );
  XOR2XL U40426 ( .A(n33724), .B(n36828), .Y(n44266) );
  XOR2XL U40427 ( .A(n36748), .B(n33940), .Y(n47044) );
  XOR2XL U40428 ( .A(n36746), .B(n34068), .Y(n47291) );
  XOR2XL U40429 ( .A(n34001), .B(n36782), .Y(n45665) );
  XOR2XL U40430 ( .A(n33897), .B(n36776), .Y(n46123) );
  XOR2XL U40431 ( .A(n33956), .B(n36823), .Y(n44229) );
  XOR2XL U40432 ( .A(n36750), .B(n33684), .Y(n47174) );
  XOR2XL U40433 ( .A(n33980), .B(n36827), .Y(n44217) );
  NOR2XL U40434 ( .A(n10863), .B(n47043), .Y(net211478) );
  XOR2XL U40435 ( .A(n36742), .B(n33948), .Y(n47043) );
  XOR2XL U40436 ( .A(n36735), .B(n33986), .Y(n47026) );
  XOR2XL U40437 ( .A(n41304), .B(n33684), .Y(n46168) );
  XOR2XL U40438 ( .A(n33833), .B(n36786), .Y(n46153) );
  XNOR2XL U40439 ( .A(n36776), .B(n34377), .Y(n46487) );
  XOR2XL U40440 ( .A(n33940), .B(n36831), .Y(n44228) );
  XOR2XL U40441 ( .A(n33828), .B(n36831), .Y(n43648) );
  XOR2XL U40442 ( .A(n42067), .B(n36883), .Y(n44923) );
  XOR2XL U40443 ( .A(n34274), .B(n41641), .Y(n45334) );
  XOR2XL U40444 ( .A(n42081), .B(n36887), .Y(n45333) );
  XOR2XL U40445 ( .A(n34004), .B(n36828), .Y(n44188) );
  XOR2XL U40446 ( .A(n33748), .B(n36823), .Y(n44307) );
  XOR2XL U40447 ( .A(n36771), .B(n33761), .Y(n47216) );
  NOR2X2 U40448 ( .A(n10378), .B(n43644), .Y(net216020) );
  XOR2XL U40449 ( .A(n33876), .B(n36827), .Y(n43644) );
  XOR2XL U40450 ( .A(n36918), .B(n33708), .Y(n46170) );
  XOR2XL U40451 ( .A(n36749), .B(n33444), .Y(n47068) );
  XNOR2XL U40452 ( .A(n42471), .B(n34352), .Y(n47643) );
  XOR2XL U40453 ( .A(n33788), .B(n36825), .Y(n45644) );
  XOR2XL U40454 ( .A(n33780), .B(n36822), .Y(n46172) );
  XOR2XL U40455 ( .A(n36766), .B(n34001), .Y(n47022) );
  XOR2XL U40456 ( .A(n33628), .B(n36822), .Y(n44427) );
  XOR2XL U40457 ( .A(n33609), .B(n36783), .Y(n45722) );
  NOR2X2 U40458 ( .A(n11731), .B(n44256), .Y(n44260) );
  XOR2XL U40459 ( .A(n33700), .B(n36829), .Y(n44256) );
  XOR2XL U40460 ( .A(n36740), .B(n33708), .Y(n47179) );
  XOR2XL U40461 ( .A(n36742), .B(n33956), .Y(n47041) );
  XOR2XL U40462 ( .A(n36736), .B(n33922), .Y(n47243) );
  XOR2XL U40463 ( .A(n36771), .B(n34081), .Y(n47281) );
  XOR2XL U40464 ( .A(n33881), .B(n36777), .Y(n46108) );
  XOR2XL U40465 ( .A(n33804), .B(n36830), .Y(n44282) );
  XOR2XL U40466 ( .A(n36733), .B(n33730), .Y(n47154) );
  XOR2XL U40467 ( .A(n33996), .B(n36829), .Y(n44202) );
  XOR2XL U40468 ( .A(n33692), .B(n36829), .Y(n44247) );
  NOR2XL U40469 ( .A(n12062), .B(n47199), .Y(n47203) );
  XOR2XL U40470 ( .A(n33460), .B(n36824), .Y(n43755) );
  XOR2XL U40471 ( .A(n34100), .B(n36825), .Y(n43837) );
  NOR2X2 U40472 ( .A(n46184), .B(n48188), .Y(n46188) );
  XOR2XL U40473 ( .A(n34089), .B(n36785), .Y(n46179) );
  XOR2XL U40474 ( .A(n34020), .B(n36824), .Y(n44164) );
  XOR2XL U40475 ( .A(n41304), .B(n33724), .Y(n45628) );
  XOR2XL U40476 ( .A(n34092), .B(n36828), .Y(n43829) );
  XOR2XL U40477 ( .A(n33593), .B(n36783), .Y(n45733) );
  XOR2XL U40478 ( .A(n33892), .B(n36823), .Y(n43630) );
  XOR2XL U40479 ( .A(n36743), .B(n33980), .Y(n47892) );
  XOR2XL U40480 ( .A(n33865), .B(n36785), .Y(n46133) );
  XOR2XL U40481 ( .A(n33900), .B(n36825), .Y(n43639) );
  XOR2XL U40482 ( .A(n34028), .B(n36825), .Y(n44173) );
  NOR2X2 U40483 ( .A(n12311), .B(n47882), .Y(n47886) );
  XOR2XL U40484 ( .A(n36744), .B(n33716), .Y(n47882) );
  XOR2XL U40485 ( .A(n34049), .B(n36764), .Y(n47002) );
  XOR2XL U40486 ( .A(n33577), .B(n36779), .Y(n45773) );
  XOR2XL U40487 ( .A(n36766), .B(n33873), .Y(n47253) );
  NOR2XL U40488 ( .A(n12726), .B(n45649), .Y(n45653) );
  XOR2XL U40489 ( .A(n33777), .B(n36777), .Y(n45649) );
  XOR2XL U40490 ( .A(n33772), .B(n36825), .Y(n44313) );
  XOR2XL U40491 ( .A(n36778), .B(n34113), .Y(n46205) );
  NOR2XL U40492 ( .A(n11138), .B(n47031), .Y(n47035) );
  XOR2XL U40493 ( .A(n36733), .B(n33994), .Y(n47031) );
  XOR2XL U40494 ( .A(n33964), .B(n36830), .Y(n44222) );
  XOR2XL U40495 ( .A(n33844), .B(n36830), .Y(n43559) );
  XOR2XL U40496 ( .A(n41304), .B(n33932), .Y(n46088) );
  XOR2XL U40497 ( .A(n36772), .B(n34017), .Y(n47024) );
  XOR2XL U40498 ( .A(n34418), .B(n42669), .Y(n45036) );
  XOR2XL U40499 ( .A(n41299), .B(n33948), .Y(n45705) );
  NOR2X2 U40500 ( .A(n10845), .B(n47169), .Y(n47173) );
  XOR2XL U40501 ( .A(n36743), .B(n33700), .Y(n47169) );
  XOR2XL U40502 ( .A(n36767), .B(n34025), .Y(n47023) );
  XOR2XL U40503 ( .A(n36740), .B(n33972), .Y(n47887) );
  XOR2XL U40504 ( .A(n34097), .B(n36785), .Y(n46195) );
  NOR2XL U40505 ( .A(n12079), .B(n46098), .Y(n46102) );
  XOR2XL U40506 ( .A(n33913), .B(n36783), .Y(n46098) );
  XOR2XL U40507 ( .A(n36734), .B(n34114), .Y(n47562) );
  XOR2XL U40508 ( .A(n36764), .B(n34097), .Y(n47552) );
  XOR2XL U40509 ( .A(n34225), .B(n42717), .Y(n44657) );
  XOR2XL U40510 ( .A(n34226), .B(n42707), .Y(n44656) );
  XOR2XL U40511 ( .A(n34228), .B(n42698), .Y(n44654) );
  XOR2X1 U40512 ( .A(n34329), .B(n34435), .Y(n45432) );
  XOR2XL U40513 ( .A(n42074), .B(n36883), .Y(n45430) );
  XNOR2XL U40514 ( .A(n34337), .B(n36875), .Y(n41726) );
  XOR2XL U40515 ( .A(n34345), .B(n34435), .Y(n45212) );
  XOR2XL U40516 ( .A(n34346), .B(n42706), .Y(n45211) );
  XOR2XL U40517 ( .A(n42072), .B(n36882), .Y(n45210) );
  XNOR2XL U40518 ( .A(n34241), .B(n34435), .Y(n41728) );
  XNOR2XL U40519 ( .A(n34242), .B(n42704), .Y(n41729) );
  XNOR2XL U40520 ( .A(n34321), .B(n34435), .Y(n41732) );
  XNOR2XL U40521 ( .A(n34322), .B(n41641), .Y(n41733) );
  XOR2XL U40522 ( .A(n34281), .B(n34435), .Y(n45304) );
  XOR2XL U40523 ( .A(n34282), .B(n42704), .Y(n45303) );
  XOR2XL U40524 ( .A(n34313), .B(n36875), .Y(n45481) );
  XOR2X1 U40525 ( .A(n34314), .B(n41641), .Y(n45480) );
  XOR2XL U40526 ( .A(n42076), .B(n36885), .Y(n45479) );
  XOR2XL U40527 ( .A(n34265), .B(n34435), .Y(n44868) );
  XOR2XL U40528 ( .A(n34266), .B(n41641), .Y(n44867) );
  XOR2XL U40529 ( .A(n42082), .B(n36886), .Y(n44866) );
  XOR2XL U40530 ( .A(n34108), .B(n36825), .Y(n43850) );
  XNOR2XL U40531 ( .A(n34256), .B(n42506), .Y(net214390) );
  XNOR2XL U40532 ( .A(n42471), .B(n34336), .Y(n47599) );
  NOR4X2 U40533 ( .A(n46517), .B(n46516), .C(n46515), .D(n46514), .Y(n46518)
         );
  XNOR2XL U40534 ( .A(n36767), .B(n34385), .Y(n47688) );
  XOR2XL U40535 ( .A(n41296), .B(n34422), .Y(n46600) );
  NOR2X1 U40536 ( .A(n45282), .B(n45281), .Y(n45286) );
  XOR2XL U40537 ( .A(n34378), .B(n41642), .Y(n44960) );
  XNOR2X1 U40538 ( .A(n34377), .B(n42579), .Y(n44902) );
  XNOR2XL U40539 ( .A(n36736), .B(n33810), .Y(n47142) );
  XNOR2XL U40540 ( .A(n36735), .B(n33554), .Y(n46913) );
  XNOR2XL U40541 ( .A(n36838), .B(n33586), .Y(n45720) );
  NAND4X2 U40542 ( .A(n46162), .B(n46161), .C(n46160), .D(n46159), .Y(n11117)
         );
  XNOR2XL U40543 ( .A(n36847), .B(n33826), .Y(n46161) );
  XNOR2XL U40544 ( .A(n36843), .B(n33514), .Y(n45801) );
  XNOR2XL U40545 ( .A(n33434), .B(n34452), .Y(n43730) );
  NAND4X2 U40546 ( .A(n45787), .B(n45786), .C(n45785), .D(n45784), .Y(n11083)
         );
  XNOR2XL U40547 ( .A(n36843), .B(n33562), .Y(n45786) );
  NAND4X2 U40548 ( .A(n47082), .B(n47081), .C(n47080), .D(n47079), .Y(n11372)
         );
  XNOR2XL U40549 ( .A(n36733), .B(n33538), .Y(n47081) );
  NAND4X2 U40550 ( .A(n45909), .B(n45908), .C(n45907), .D(n45906), .Y(n11054)
         );
  XNOR2XL U40551 ( .A(n36845), .B(n33394), .Y(n45908) );
  XNOR2XL U40552 ( .A(n36733), .B(n33362), .Y(n46747) );
  XNOR2XL U40553 ( .A(n36841), .B(n33938), .Y(n45698) );
  XNOR2XL U40554 ( .A(n36839), .B(n33554), .Y(n45771) );
  XNOR2XL U40555 ( .A(n36736), .B(n33394), .Y(n46722) );
  XNOR2XL U40556 ( .A(n33418), .B(n36725), .Y(n43217) );
  XNOR2XL U40557 ( .A(n36840), .B(n33482), .Y(net213116) );
  XNOR2XL U40558 ( .A(n36838), .B(n33546), .Y(n45826) );
  XNOR2XL U40559 ( .A(n36734), .B(n33746), .Y(net211262) );
  XNOR2XL U40560 ( .A(n33450), .B(n34452), .Y(n43712) );
  XNOR2XL U40561 ( .A(n36837), .B(n33530), .Y(n45836) );
  XNOR2XL U40562 ( .A(n33522), .B(n42569), .Y(n43785) );
  XNOR2XL U40563 ( .A(n33506), .B(n34452), .Y(n43703) );
  XNOR2XL U40564 ( .A(n36846), .B(n33874), .Y(n46116) );
  XNOR2XL U40565 ( .A(n36839), .B(n33858), .Y(n46131) );
  XNOR2XL U40566 ( .A(n36844), .B(n33426), .Y(n45841) );
  XNOR2XL U40567 ( .A(n33386), .B(n42569), .Y(n43279) );
  XNOR2XL U40568 ( .A(n36845), .B(n33458), .Y(n45862) );
  XNOR2XL U40569 ( .A(n36733), .B(n33850), .Y(n47231) );
  NAND4X2 U40570 ( .A(n47077), .B(n47076), .C(n47075), .D(n47074), .Y(n11371)
         );
  XNOR2XL U40571 ( .A(n36735), .B(n33546), .Y(n47076) );
  XNOR2XL U40572 ( .A(n36735), .B(n33386), .Y(n46762) );
  NAND4X2 U40573 ( .A(n47067), .B(n47066), .C(n47065), .D(n47064), .Y(n11358)
         );
  XNOR2XL U40574 ( .A(n36733), .B(n33450), .Y(n47066) );
  XNOR2XL U40575 ( .A(n33578), .B(n41630), .Y(n44559) );
  XNOR2XL U40576 ( .A(n36735), .B(n33834), .Y(n47137) );
  XNOR2XL U40577 ( .A(n36736), .B(n33578), .Y(n46918) );
  XNOR2XL U40578 ( .A(n36735), .B(n33378), .Y(n46772) );
  XNOR2XL U40579 ( .A(n36734), .B(n33458), .Y(n47121) );
  XNOR2XL U40580 ( .A(n33594), .B(n41630), .Y(n44515) );
  XNOR2XL U40581 ( .A(n36736), .B(n33562), .Y(n46908) );
  XNOR2XL U40582 ( .A(n36733), .B(n33818), .Y(n47147) );
  NAND4X2 U40583 ( .A(n47168), .B(n47167), .C(n47166), .D(n47165), .Y(n11397)
         );
  XNOR2XL U40584 ( .A(n36735), .B(n33690), .Y(n47167) );
  XNOR2XL U40585 ( .A(n36733), .B(n33402), .Y(n46717) );
  XNOR2XL U40586 ( .A(n36734), .B(n33410), .Y(n46712) );
  XNOR2XL U40587 ( .A(n36735), .B(n33370), .Y(n46757) );
  XNOR2XL U40588 ( .A(n36847), .B(n33842), .Y(n46141) );
  XNOR2XL U40589 ( .A(n36844), .B(n33410), .Y(n45918) );
  XNOR2XL U40590 ( .A(n36845), .B(n33730), .Y(n45626) );
  XNOR2XL U40591 ( .A(n36840), .B(n33442), .Y(n45851) );
  XOR2XL U40592 ( .A(n34321), .B(n42575), .Y(n45190) );
  XOR2XL U40593 ( .A(n42554), .B(n34117), .Y(n43877) );
  XOR2XL U40594 ( .A(n36846), .B(n34202), .Y(n46407) );
  XOR2XL U40595 ( .A(n36844), .B(n34210), .Y(n46396) );
  XOR2XL U40596 ( .A(n36733), .B(n34210), .Y(n47397) );
  XOR2XL U40597 ( .A(n36734), .B(n34202), .Y(n47408) );
  XOR2XL U40598 ( .A(n42544), .B(n34118), .Y(n43876) );
  XOR2XL U40599 ( .A(n36780), .B(n34201), .Y(n46405) );
  XOR2XL U40600 ( .A(n36765), .B(n34201), .Y(n47406) );
  XOR2XL U40601 ( .A(n36734), .B(n34370), .Y(n47618) );
  XOR2XL U40602 ( .A(n36843), .B(n34346), .Y(n46550) );
  XOR2XL U40603 ( .A(n36843), .B(n34314), .Y(n46349) );
  XOR2XL U40604 ( .A(n36838), .B(n34338), .Y(n46539) );
  XOR2XL U40605 ( .A(n36844), .B(n34330), .Y(n46517) );
  XOR2XL U40606 ( .A(n36843), .B(n34258), .Y(n46382) );
  XOR2XL U40607 ( .A(n36734), .B(n34362), .Y(n47607) );
  XOR2XL U40608 ( .A(n36838), .B(n34282), .Y(n46360) );
  XOR2XL U40609 ( .A(n36847), .B(n34322), .Y(n46528) );
  XOR2XL U40610 ( .A(n36733), .B(n34346), .Y(n47640) );
  XOR2XL U40611 ( .A(n36846), .B(n34274), .Y(n46371) );
  XOR2XL U40612 ( .A(n36839), .B(n34290), .Y(n46338) );
  XOR2XL U40613 ( .A(n36736), .B(n34354), .Y(n47629) );
  XOR2XL U40614 ( .A(n36839), .B(n34298), .Y(n46327) );
  XOR2XL U40615 ( .A(n36841), .B(n34242), .Y(n46469) );
  XOR2XL U40616 ( .A(n36837), .B(n34266), .Y(n46389) );
  XOR2XL U40617 ( .A(n36735), .B(n34322), .Y(n47585) );
  XOR2XL U40618 ( .A(n36734), .B(n34298), .Y(n47320) );
  XOR2XL U40619 ( .A(n36734), .B(n34282), .Y(n47342) );
  XOR2XL U40620 ( .A(n36734), .B(n34266), .Y(n47375) );
  XOR2XL U40621 ( .A(n36735), .B(n34274), .Y(n47353) );
  XOR2XL U40622 ( .A(n36735), .B(n34330), .Y(n47596) );
  XOR2XL U40623 ( .A(n36733), .B(n34258), .Y(n47364) );
  XOR2XL U40624 ( .A(n36736), .B(n34242), .Y(n47441) );
  XNOR2XL U40625 ( .A(n36734), .B(n33418), .Y(n46707) );
  XOR2XL U40626 ( .A(n42471), .B(n34168), .Y(n47508) );
  XOR2XL U40627 ( .A(n36735), .B(n34178), .Y(n47485) );
  XOR2XL U40628 ( .A(n36780), .B(n34329), .Y(n46515) );
  XOR2XL U40629 ( .A(n41299), .B(n34228), .Y(n46438) );
  XOR2XL U40630 ( .A(n41302), .B(n34260), .Y(n46380) );
  XOR2XL U40631 ( .A(n36785), .B(n34321), .Y(n46526) );
  XOR2XL U40632 ( .A(n36774), .B(n34337), .Y(n47646) );
  XOR2XL U40633 ( .A(n36774), .B(n34305), .Y(n47305) );
  XOR2XL U40634 ( .A(n36771), .B(n34321), .Y(n47583) );
  XOR2XL U40635 ( .A(n36778), .B(n34209), .Y(n46394) );
  XOR2XL U40636 ( .A(n36744), .B(n34228), .Y(n47461) );
  XOR2XL U40637 ( .A(n36766), .B(n34209), .Y(n47395) );
  XOR2XL U40638 ( .A(n36770), .B(n34329), .Y(n47594) );
  XOR2XL U40639 ( .A(n36746), .B(n34260), .Y(n47362) );
  XOR2XL U40640 ( .A(n36845), .B(n34226), .Y(n46440) );
  XOR2XL U40641 ( .A(n36841), .B(n34170), .Y(n46255) );
  XOR2XL U40642 ( .A(n36847), .B(n34234), .Y(n46451) );
  XOR2XL U40643 ( .A(n36845), .B(n34154), .Y(n46300) );
  XOR2XL U40644 ( .A(n36837), .B(n34218), .Y(n46429) );
  XOR2XL U40645 ( .A(n36847), .B(n34146), .Y(n46227) );
  XOR2XL U40646 ( .A(n36715), .B(n34341), .Y(n47652) );
  XOR2XL U40647 ( .A(n36837), .B(n34138), .Y(n46277) );
  XOR2XL U40648 ( .A(n36843), .B(n34162), .Y(n46266) );
  XOR2XL U40649 ( .A(n36840), .B(n34194), .Y(n46418) );
  XOR2XL U40650 ( .A(n36846), .B(n34186), .Y(n46238) );
  XOR2XL U40651 ( .A(n36840), .B(n34250), .Y(n46462) );
  XOR2XL U40652 ( .A(n36733), .B(n34170), .Y(n47496) );
  XOR2XL U40653 ( .A(n36734), .B(n34250), .Y(n47430) );
  XOR2XL U40654 ( .A(n36733), .B(n34226), .Y(n47463) );
  XOR2XL U40655 ( .A(n36734), .B(n34234), .Y(n47452) );
  XOR2XL U40656 ( .A(n36736), .B(n34218), .Y(n47386) );
  XOR2XL U40657 ( .A(n36733), .B(n34146), .Y(n47516) );
  XOR2XL U40658 ( .A(n36736), .B(n34138), .Y(n47538) );
  XOR2XL U40659 ( .A(n36733), .B(n34154), .Y(n47527) );
  XOR2XL U40660 ( .A(n36736), .B(n34194), .Y(n47419) );
  XOR2XL U40661 ( .A(n36735), .B(n34186), .Y(n47474) );
  XOR2XL U40662 ( .A(n36777), .B(n34345), .Y(n46549) );
  XOR2XL U40663 ( .A(n36778), .B(n34353), .Y(n46494) );
  XOR2XL U40664 ( .A(n36782), .B(n34337), .Y(n46538) );
  XOR2XL U40665 ( .A(n36776), .B(n34305), .Y(n46315) );
  XOR2XL U40666 ( .A(n36777), .B(n34257), .Y(n46381) );
  XOR2XL U40667 ( .A(n36783), .B(n34281), .Y(n46359) );
  XOR2XL U40668 ( .A(n36765), .B(n34345), .Y(n47639) );
  XOR2XL U40669 ( .A(n36777), .B(n34273), .Y(n46370) );
  XOR2XL U40670 ( .A(n36776), .B(n34289), .Y(n46337) );
  XOR2XL U40671 ( .A(n36773), .B(n34353), .Y(n47628) );
  XOR2XL U40672 ( .A(n36786), .B(n34297), .Y(n46326) );
  XOR2XL U40673 ( .A(n36782), .B(n34241), .Y(n46468) );
  XOR2XL U40674 ( .A(n36786), .B(n34265), .Y(n46388) );
  XOR2XL U40675 ( .A(n36736), .B(n34338), .Y(n47647) );
  XOR2XL U40676 ( .A(n36735), .B(n34306), .Y(n47306) );
  XOR2XL U40677 ( .A(n36773), .B(n34297), .Y(n47319) );
  XOR2XL U40678 ( .A(n36770), .B(n34281), .Y(n47341) );
  XOR2XL U40679 ( .A(n36770), .B(n34265), .Y(n47374) );
  XOR2XL U40680 ( .A(n36767), .B(n34273), .Y(n47352) );
  XOR2XL U40681 ( .A(n36772), .B(n34289), .Y(n47330) );
  XOR2XL U40682 ( .A(n36771), .B(n34257), .Y(n47363) );
  XOR2XL U40683 ( .A(n36768), .B(n34241), .Y(n47440) );
  XOR2XL U40684 ( .A(n36750), .B(n34180), .Y(n47483) );
  XOR2XL U40685 ( .A(n41303), .B(n34172), .Y(n46253) );
  XOR2XL U40686 ( .A(n36918), .B(n34236), .Y(n46449) );
  XOR2XL U40687 ( .A(n41299), .B(n34156), .Y(n46298) );
  XOR2XL U40688 ( .A(n41304), .B(n34220), .Y(n46427) );
  XOR2XL U40689 ( .A(n41301), .B(n34148), .Y(n46225) );
  XOR2XL U40690 ( .A(n41305), .B(n34284), .Y(n46358) );
  XOR2XL U40691 ( .A(n41302), .B(n34124), .Y(n46214) );
  XOR2XL U40692 ( .A(n41300), .B(n34140), .Y(n46275) );
  XOR2XL U40693 ( .A(n41299), .B(n34164), .Y(n46264) );
  XOR2XL U40694 ( .A(n41305), .B(n34292), .Y(n46336) );
  XOR2XL U40695 ( .A(n36779), .B(n34193), .Y(n46416) );
  XOR2XL U40696 ( .A(n36780), .B(n34185), .Y(n46236) );
  XOR2XL U40697 ( .A(n41301), .B(n34244), .Y(n46467) );
  XOR2XL U40698 ( .A(n41303), .B(n34252), .Y(n46460) );
  XOR2XL U40699 ( .A(n36764), .B(n34161), .Y(n47502) );
  XOR2XL U40700 ( .A(n36795), .B(n34166), .Y(n47506) );
  XOR2XL U40701 ( .A(n36742), .B(n34172), .Y(n47494) );
  XOR2XL U40702 ( .A(n36750), .B(n34252), .Y(n47428) );
  XOR2XL U40703 ( .A(n36749), .B(n34148), .Y(n47514) );
  XOR2XL U40704 ( .A(n36747), .B(n34284), .Y(n47340) );
  XOR2XL U40705 ( .A(n36749), .B(n34236), .Y(n47450) );
  XOR2XL U40706 ( .A(n36743), .B(n34220), .Y(n47384) );
  XOR2XL U40707 ( .A(n36746), .B(n34140), .Y(n47536) );
  XOR2XL U40708 ( .A(n36748), .B(n34156), .Y(n47525) );
  XOR2XL U40709 ( .A(n36796), .B(n34310), .Y(n47309) );
  XOR2XL U40710 ( .A(n36774), .B(n34193), .Y(n47417) );
  XOR2XL U40711 ( .A(n36748), .B(n34292), .Y(n47329) );
  XOR2XL U40712 ( .A(n36768), .B(n34185), .Y(n47472) );
  XOR2XL U40713 ( .A(n36743), .B(n34244), .Y(n47439) );
  XOR2XL U40714 ( .A(n36766), .B(n34177), .Y(n47484) );
  XOR2XL U40715 ( .A(n41304), .B(n34316), .Y(n46348) );
  XOR2XL U40716 ( .A(n36776), .B(n34169), .Y(n46254) );
  XOR2XL U40717 ( .A(n36777), .B(n34225), .Y(n46439) );
  XOR2XL U40718 ( .A(n36780), .B(n34153), .Y(n46299) );
  XOR2XL U40719 ( .A(n36779), .B(n34233), .Y(n46450) );
  XOR2XL U40720 ( .A(n36784), .B(n34217), .Y(n46428) );
  XOR2XL U40721 ( .A(n36777), .B(n34145), .Y(n46226) );
  XOR2XL U40722 ( .A(n36778), .B(n34161), .Y(n46265) );
  XOR2XL U40723 ( .A(n41301), .B(n34204), .Y(n46406) );
  XOR2XL U40724 ( .A(n36792), .B(n34342), .Y(n47651) );
  XOR2XL U40725 ( .A(n41300), .B(n34196), .Y(n46417) );
  XOR2XL U40726 ( .A(n41300), .B(n34188), .Y(n46237) );
  XOR2XL U40727 ( .A(n36778), .B(n34249), .Y(n46461) );
  XOR2XL U40728 ( .A(n36746), .B(n34324), .Y(n47584) );
  XOR2XL U40729 ( .A(n41303), .B(n34212), .Y(n46395) );
  XOR2XL U40730 ( .A(n36721), .B(n34165), .Y(n47507) );
  XOR2XL U40731 ( .A(n36772), .B(n34169), .Y(n47495) );
  XOR2XL U40732 ( .A(n36766), .B(n34249), .Y(n47429) );
  XOR2XL U40733 ( .A(n36767), .B(n34225), .Y(n47462) );
  XOR2XL U40734 ( .A(n36750), .B(n34316), .Y(n47298) );
  XOR2XL U40735 ( .A(n36765), .B(n34145), .Y(n47515) );
  XOR2XL U40736 ( .A(n36773), .B(n34233), .Y(n47451) );
  XOR2XL U40737 ( .A(n36764), .B(n34217), .Y(n47385) );
  XOR2XL U40738 ( .A(n36740), .B(n34212), .Y(n47396) );
  XOR2XL U40739 ( .A(n36774), .B(n34153), .Y(n47526) );
  XOR2XL U40740 ( .A(n36740), .B(n34196), .Y(n47418) );
  XOR2XL U40741 ( .A(n36743), .B(n34188), .Y(n47473) );
  XOR2XL U40742 ( .A(n36749), .B(n34204), .Y(n47407) );
  XOR2XL U40743 ( .A(n36744), .B(n34164), .Y(n47505) );
  XOR2XL U40744 ( .A(n36841), .B(n34370), .Y(n46476) );
  XOR2XL U40745 ( .A(n36837), .B(n34362), .Y(n46508) );
  XOR2XL U40746 ( .A(n36718), .B(n34373), .Y(n47614) );
  XOR2XL U40747 ( .A(n36718), .B(n34181), .Y(n47481) );
  XOR2XL U40748 ( .A(n41333), .B(n34357), .Y(n46491) );
  XOR2XL U40749 ( .A(n41327), .B(n34349), .Y(n46546) );
  XOR2XL U40750 ( .A(n41329), .B(n34341), .Y(n46535) );
  XOR2XL U40751 ( .A(n36913), .B(n34333), .Y(n46513) );
  XOR2XL U40752 ( .A(n41330), .B(n34229), .Y(n46436) );
  XOR2XL U40753 ( .A(n36716), .B(n34365), .Y(n47603) );
  XOR2XL U40754 ( .A(n41327), .B(n34173), .Y(n46251) );
  XOR2XL U40755 ( .A(n41332), .B(n34261), .Y(n46378) );
  XOR2XL U40756 ( .A(n41329), .B(n34237), .Y(n46447) );
  XOR2XL U40757 ( .A(n36913), .B(n34157), .Y(n46296) );
  XOR2XL U40758 ( .A(n41330), .B(n34309), .Y(n46312) );
  XOR2XL U40759 ( .A(n41331), .B(n34221), .Y(n46425) );
  XOR2XL U40760 ( .A(n41328), .B(n34325), .Y(n46524) );
  XOR2XL U40761 ( .A(n41331), .B(n34285), .Y(n46356) );
  XOR2XL U40762 ( .A(n36715), .B(n34349), .Y(n47636) );
  XOR2XL U40763 ( .A(n41332), .B(n34165), .Y(n46262) );
  XOR2XL U40764 ( .A(n41330), .B(n34125), .Y(n46212) );
  XOR2XL U40765 ( .A(n41329), .B(n34277), .Y(n46367) );
  XOR2XL U40766 ( .A(n41333), .B(n34293), .Y(n46334) );
  XOR2XL U40767 ( .A(n41331), .B(n34205), .Y(n46403) );
  XOR2XL U40768 ( .A(n41330), .B(n34245), .Y(n46465) );
  XOR2XL U40769 ( .A(n36718), .B(n34357), .Y(n47625) );
  XOR2XL U40770 ( .A(n41331), .B(n34301), .Y(n46323) );
  XOR2XL U40771 ( .A(n41327), .B(n34197), .Y(n46414) );
  XOR2XL U40772 ( .A(n41327), .B(n34269), .Y(n46385) );
  XOR2XL U40773 ( .A(n41332), .B(n34253), .Y(n46458) );
  XOR2XL U40774 ( .A(n41328), .B(n34149), .Y(n46223) );
  XOR2XL U40775 ( .A(n41328), .B(n34213), .Y(n46392) );
  XOR2XL U40776 ( .A(n36717), .B(n34173), .Y(n47492) );
  XOR2XL U40777 ( .A(n36716), .B(n34325), .Y(n47581) );
  XOR2XL U40778 ( .A(n36714), .B(n34253), .Y(n47426) );
  XOR2XL U40779 ( .A(n36714), .B(n34229), .Y(n47459) );
  XOR2XL U40780 ( .A(n36717), .B(n34317), .Y(n47295) );
  XOR2XL U40781 ( .A(n36721), .B(n34285), .Y(n47338) );
  XOR2XL U40782 ( .A(n36718), .B(n34237), .Y(n47448) );
  XOR2XL U40783 ( .A(n36716), .B(n34221), .Y(n47382) );
  XOR2XL U40784 ( .A(n36720), .B(n34269), .Y(n47371) );
  XOR2XL U40785 ( .A(n36722), .B(n34149), .Y(n47512) );
  XOR2XL U40786 ( .A(n36722), .B(n34333), .Y(n47592) );
  XOR2XL U40787 ( .A(n41331), .B(n34189), .Y(n46234) );
  XOR2XL U40788 ( .A(n36716), .B(n34277), .Y(n47349) );
  XOR2XL U40789 ( .A(n36722), .B(n34213), .Y(n47393) );
  XOR2XL U40790 ( .A(n36715), .B(n34157), .Y(n47523) );
  XOR2XL U40791 ( .A(n36717), .B(n34189), .Y(n47470) );
  XOR2XL U40792 ( .A(n36718), .B(n34197), .Y(n47415) );
  XOR2XL U40793 ( .A(n36720), .B(n34293), .Y(n47327) );
  XOR2XL U40794 ( .A(n36722), .B(n34261), .Y(n47360) );
  XOR2XL U40795 ( .A(n36721), .B(n34245), .Y(n47437) );
  XOR2XL U40796 ( .A(n36720), .B(n34205), .Y(n47404) );
  XNOR2XL U40797 ( .A(n42471), .B(n34128), .Y(n47576) );
  XOR2XL U40798 ( .A(n34124), .B(n36831), .Y(n43911) );
  XOR2XL U40799 ( .A(n34116), .B(n36827), .Y(n43880) );
  XOR2XL U40800 ( .A(n34261), .B(n42630), .Y(n44856) );
  XOR2XL U40801 ( .A(n36790), .B(n34374), .Y(n47613) );
  XOR2XL U40802 ( .A(n34320), .B(n36731), .Y(n45416) );
  XOR2XL U40803 ( .A(n34194), .B(n42560), .Y(n44728) );
  XNOR2XL U40804 ( .A(n36764), .B(n34377), .Y(n47653) );
  XOR2XL U40805 ( .A(n34309), .B(n42629), .Y(n45469) );
  XOR2XL U40806 ( .A(n34297), .B(n41319), .Y(n45499) );
  XOR2XL U40807 ( .A(n34309), .B(n41282), .Y(n45503) );
  XOR2XL U40808 ( .A(n34269), .B(n42624), .Y(n45323) );
  XOR2XL U40809 ( .A(n34257), .B(n36905), .Y(n44860) );
  XOR2XL U40810 ( .A(n34277), .B(n41283), .Y(n45331) );
  XOR2XL U40811 ( .A(n34289), .B(n42684), .Y(n45385) );
  XOR2XL U40812 ( .A(n34253), .B(n41282), .Y(n44775) );
  XOR2XL U40813 ( .A(n34241), .B(n41379), .Y(n44771) );
  XNOR2XL U40814 ( .A(n36733), .B(n33434), .Y(n47061) );
  XNOR2XL U40815 ( .A(n36779), .B(n34177), .Y(n46246) );
  XNOR2XL U40816 ( .A(n41296), .B(n34182), .Y(n46242) );
  XNOR2XL U40817 ( .A(n36722), .B(n34381), .Y(n47658) );
  XOR2XL U40818 ( .A(n34189), .B(n41282), .Y(n44082) );
  XOR2XL U40819 ( .A(n34213), .B(n41282), .Y(n44715) );
  XOR2XL U40820 ( .A(n34177), .B(n36905), .Y(n44078) );
  XOR2XL U40821 ( .A(n34201), .B(n41319), .Y(n44711) );
  XNOR2XL U40822 ( .A(n41305), .B(n34180), .Y(n46241) );
  XOR2XL U40823 ( .A(n36720), .B(n34389), .Y(n47685) );
  XOR2XL U40824 ( .A(n36799), .B(n34182), .Y(n47480) );
  XOR2XL U40825 ( .A(n34298), .B(n42672), .Y(n45498) );
  XOR2XL U40826 ( .A(n34266), .B(n42669), .Y(n45326) );
  XOR2XL U40827 ( .A(n34281), .B(n42576), .Y(n45402) );
  XOR2XL U40828 ( .A(n34257), .B(n42576), .Y(n45340) );
  XOR2XL U40829 ( .A(n34289), .B(n42576), .Y(n45516) );
  XOR2XL U40830 ( .A(n34297), .B(n42576), .Y(n45489) );
  XOR2XL U40831 ( .A(n41297), .B(n34318), .Y(n46344) );
  XOR2XL U40832 ( .A(n41291), .B(n34342), .Y(n46534) );
  XOR2XL U40833 ( .A(n36916), .B(n34334), .Y(n46512) );
  XOR2XL U40834 ( .A(n41291), .B(n34230), .Y(n46435) );
  XOR2XL U40835 ( .A(n36797), .B(n34366), .Y(n47602) );
  XOR2XL U40836 ( .A(n41293), .B(n34262), .Y(n46377) );
  XOR2XL U40837 ( .A(n41293), .B(n34238), .Y(n46446) );
  XOR2XL U40838 ( .A(n41294), .B(n34158), .Y(n46295) );
  XOR2XL U40839 ( .A(n41295), .B(n34310), .Y(n46311) );
  XOR2XL U40840 ( .A(n41295), .B(n34222), .Y(n46424) );
  XOR2XL U40841 ( .A(n41294), .B(n34326), .Y(n46523) );
  XOR2XL U40842 ( .A(n36789), .B(n34350), .Y(n47635) );
  XOR2XL U40843 ( .A(n41294), .B(n34286), .Y(n46355) );
  XOR2XL U40844 ( .A(n41292), .B(n34166), .Y(n46261) );
  XOR2XL U40845 ( .A(n41292), .B(n34278), .Y(n46366) );
  XOR2XL U40846 ( .A(n41296), .B(n34294), .Y(n46333) );
  XOR2XL U40847 ( .A(n41294), .B(n34246), .Y(n46464) );
  XOR2XL U40848 ( .A(n41291), .B(n34206), .Y(n46402) );
  XOR2XL U40849 ( .A(n36796), .B(n34358), .Y(n47624) );
  XOR2XL U40850 ( .A(n41293), .B(n34302), .Y(n46322) );
  XOR2XL U40851 ( .A(n41290), .B(n34198), .Y(n46413) );
  XOR2XL U40852 ( .A(n36916), .B(n34270), .Y(n46384) );
  XOR2XL U40853 ( .A(n41296), .B(n34254), .Y(n46457) );
  XOR2XL U40854 ( .A(n41293), .B(n34174), .Y(n46250) );
  XOR2XL U40855 ( .A(n41294), .B(n34150), .Y(n46222) );
  XOR2XL U40856 ( .A(n41297), .B(n34214), .Y(n46391) );
  XOR2XL U40857 ( .A(n36791), .B(n34174), .Y(n47491) );
  XOR2XL U40858 ( .A(n36798), .B(n34326), .Y(n47580) );
  XOR2XL U40859 ( .A(n36790), .B(n34254), .Y(n47425) );
  XOR2XL U40860 ( .A(n36799), .B(n34302), .Y(n47315) );
  XOR2XL U40861 ( .A(n36793), .B(n34230), .Y(n47458) );
  XOR2XL U40862 ( .A(n36799), .B(n34318), .Y(n47294) );
  XOR2XL U40863 ( .A(n36793), .B(n34286), .Y(n47337) );
  XOR2XL U40864 ( .A(n36797), .B(n34238), .Y(n47447) );
  XOR2XL U40865 ( .A(n36796), .B(n34222), .Y(n47381) );
  XOR2XL U40866 ( .A(n36792), .B(n34270), .Y(n47370) );
  XOR2XL U40867 ( .A(n36796), .B(n34150), .Y(n47511) );
  XOR2XL U40868 ( .A(n36795), .B(n34334), .Y(n47591) );
  XOR2XL U40869 ( .A(n41296), .B(n34190), .Y(n46233) );
  XOR2XL U40870 ( .A(n36791), .B(n34278), .Y(n47348) );
  XOR2XL U40871 ( .A(n36790), .B(n34214), .Y(n47392) );
  XOR2XL U40872 ( .A(n36797), .B(n34158), .Y(n47522) );
  XOR2XL U40873 ( .A(n36789), .B(n34190), .Y(n47469) );
  XOR2XL U40874 ( .A(n36798), .B(n34198), .Y(n47414) );
  XOR2XL U40875 ( .A(n36797), .B(n34294), .Y(n47326) );
  XOR2XL U40876 ( .A(n36792), .B(n34262), .Y(n47359) );
  XOR2XL U40877 ( .A(n36789), .B(n34206), .Y(n47403) );
  XOR2XL U40878 ( .A(n36791), .B(n34246), .Y(n47436) );
  XOR2XL U40879 ( .A(n34302), .B(n40039), .Y(n45388) );
  XOR2XL U40880 ( .A(n34310), .B(net219310), .Y(n45502) );
  XOR2XL U40881 ( .A(n34270), .B(n36868), .Y(n45322) );
  XOR2XL U40882 ( .A(n34270), .B(net219310), .Y(n44863) );
  XOR2XL U40883 ( .A(n34258), .B(n42672), .Y(n44859) );
  XOR2XL U40884 ( .A(n34278), .B(net219330), .Y(n45330) );
  XOR2XL U40885 ( .A(n34254), .B(net219310), .Y(n44774) );
  XOR2XL U40886 ( .A(n34242), .B(n42669), .Y(n44770) );
  XOR2XL U40887 ( .A(n36838), .B(n34122), .Y(n46216) );
  XOR2XL U40888 ( .A(n34190), .B(net219308), .Y(n44081) );
  XOR2XL U40889 ( .A(n34214), .B(net219314), .Y(n44714) );
  XOR2XL U40890 ( .A(n34178), .B(n42671), .Y(n44077) );
  XOR2XL U40891 ( .A(n34202), .B(n36907), .Y(n44710) );
  XNOR2XL U40892 ( .A(n36793), .B(n34382), .Y(n47657) );
  XOR2XL U40893 ( .A(n42584), .B(n34121), .Y(n43910) );
  XNOR2XL U40894 ( .A(n41331), .B(n34181), .Y(n46239) );
  XOR2XL U40895 ( .A(n34304), .B(n34450), .Y(n45492) );
  XOR2XL U40896 ( .A(n36782), .B(n34121), .Y(n46215) );
  XOR2XL U40897 ( .A(n34313), .B(n42576), .Y(n45413) );
  XOR2XL U40898 ( .A(n34296), .B(n34450), .Y(n45378) );
  XOR2XL U40899 ( .A(n34308), .B(n42638), .Y(n45470) );
  XOR2XL U40900 ( .A(n34312), .B(n36863), .Y(n45466) );
  XOR2XL U40901 ( .A(n34268), .B(n42638), .Y(n45324) );
  XOR2XL U40902 ( .A(n34272), .B(n34450), .Y(n45320) );
  XOR2XL U40903 ( .A(n34264), .B(n42592), .Y(n44853) );
  XOR2XL U40904 ( .A(n34161), .B(n42584), .Y(n44064) );
  XOR2XL U40905 ( .A(n34177), .B(n42577), .Y(n44126) );
  XOR2XL U40906 ( .A(n34217), .B(n42575), .Y(n44697) );
  XOR2XL U40907 ( .A(n34201), .B(n42583), .Y(n44757) );
  XOR2XL U40908 ( .A(n34153), .B(n42577), .Y(n43941) );
  XOR2XL U40909 ( .A(n34225), .B(n42577), .Y(n44846) );
  XOR2XL U40910 ( .A(n34145), .B(n42580), .Y(n43972) );
  XOR2XL U40911 ( .A(n34169), .B(n42581), .Y(n44095) );
  XOR2XL U40912 ( .A(n34193), .B(n42581), .Y(n44726) );
  XOR2XL U40913 ( .A(n34125), .B(n41281), .Y(n43844) );
  XOR2XL U40914 ( .A(n34184), .B(n34450), .Y(n44071) );
  XOR2XL U40915 ( .A(n34208), .B(n34450), .Y(n44704) );
  NAND4X2 U40916 ( .A(n46929), .B(n46928), .C(n46927), .D(n46926), .Y(
        net210259) );
  XNOR2XL U40917 ( .A(n36772), .B(n33609), .Y(n46928) );
  XNOR2XL U40918 ( .A(n36733), .B(n33722), .Y(n47880) );
  XOR2XL U40919 ( .A(n34252), .B(n36830), .Y(n44878) );
  XOR2XL U40920 ( .A(n34164), .B(n36830), .Y(n44065) );
  XOR2XL U40921 ( .A(n34180), .B(n36822), .Y(n44127) );
  XOR2XL U40922 ( .A(n34308), .B(n36821), .Y(n45460) );
  XOR2XL U40923 ( .A(n34148), .B(n36823), .Y(n43973) );
  XOR2XL U40924 ( .A(n34212), .B(n36821), .Y(n44667) );
  XOR2XL U40925 ( .A(n34276), .B(n36821), .Y(n45372) );
  XOR2XL U40926 ( .A(n34268), .B(n36823), .Y(n45314) );
  XOR2XL U40927 ( .A(n34284), .B(n36828), .Y(n45403) );
  XOR2XL U40928 ( .A(n34172), .B(n36830), .Y(n44096) );
  XOR2XL U40929 ( .A(n34196), .B(n36829), .Y(n44727) );
  XOR2XL U40930 ( .A(n34260), .B(n36830), .Y(n45341) );
  XOR2XL U40931 ( .A(n34292), .B(n36824), .Y(n45517) );
  XOR2XL U40932 ( .A(n34300), .B(n36824), .Y(n45490) );
  XOR2XL U40933 ( .A(n34338), .B(n41630), .Y(n45132) );
  XOR2XL U40934 ( .A(n34346), .B(n41630), .Y(n45163) );
  XOR2XL U40935 ( .A(n34154), .B(n42558), .Y(n43943) );
  XOR2XL U40936 ( .A(n34226), .B(n42557), .Y(n44848) );
  XOR2XL U40937 ( .A(n34234), .B(n42557), .Y(n44790) );
  XOR2XL U40938 ( .A(n34122), .B(n42558), .Y(n43912) );
  XOR2XL U40939 ( .A(n34146), .B(n42558), .Y(n43974) );
  XOR2XL U40940 ( .A(n34210), .B(n42557), .Y(n44668) );
  XOR2XL U40941 ( .A(n34274), .B(n41630), .Y(n45373) );
  XOR2XL U40942 ( .A(n34170), .B(n42558), .Y(n44097) );
  XOR2XL U40943 ( .A(n34266), .B(n41630), .Y(n45315) );
  XOR2XL U40944 ( .A(n34282), .B(n41630), .Y(n45404) );
  XOR2XL U40945 ( .A(n34114), .B(n41630), .Y(n43881) );
  XOR2XL U40946 ( .A(n34258), .B(n41630), .Y(n45342) );
  XOR2XL U40947 ( .A(n34298), .B(n42558), .Y(n45491) );
  XOR2XL U40948 ( .A(n34250), .B(n42559), .Y(n44879) );
  XOR2XL U40949 ( .A(n34325), .B(n42549), .Y(n45188) );
  XOR2XL U40950 ( .A(n34269), .B(n42549), .Y(n45311) );
  XOR2XL U40951 ( .A(n34285), .B(n42549), .Y(n45400) );
  XOR2XL U40952 ( .A(n34277), .B(n42549), .Y(n45369) );
  XOR2XL U40953 ( .A(n34301), .B(n42549), .Y(n45487) );
  XOR2XL U40954 ( .A(n34293), .B(n42549), .Y(n45514) );
  XOR2XL U40955 ( .A(n34353), .B(n42575), .Y(n44988) );
  XOR2XL U40956 ( .A(n34241), .B(n42575), .Y(n44819) );
  XOR2XL U40957 ( .A(n34305), .B(n42575), .Y(n45459) );
  XOR2XL U40958 ( .A(n34233), .B(n42575), .Y(n44788) );
  XOR2XL U40959 ( .A(n34273), .B(n42575), .Y(n45371) );
  XOR2XL U40960 ( .A(n34265), .B(n42575), .Y(n45313) );
  XOR2XL U40961 ( .A(n34249), .B(n42575), .Y(n44877) );
  XNOR2XL U40962 ( .A(n33908), .B(n36821), .Y(n43614) );
  XNOR2XL U40963 ( .A(n33916), .B(n36823), .Y(n43601) );
  XOR2XL U40964 ( .A(n34334), .B(n42534), .Y(n45218) );
  XOR2XL U40965 ( .A(n34286), .B(n42534), .Y(n45399) );
  XOR2XL U40966 ( .A(n34302), .B(n42534), .Y(n45486) );
  XOR2XL U40967 ( .A(n34262), .B(n42534), .Y(n45337) );
  XOR2XL U40968 ( .A(n34294), .B(n42534), .Y(n45513) );
  XOR2XL U40969 ( .A(n42544), .B(n34126), .Y(n43907) );
  XOR2XL U40970 ( .A(n41294), .B(n34126), .Y(n46211) );
  XOR2XL U40971 ( .A(n42584), .B(n34113), .Y(n43879) );
  XOR2XL U40972 ( .A(n34357), .B(n36832), .Y(n44986) );
  XOR2XL U40973 ( .A(n34333), .B(n36832), .Y(n45219) );
  XOR2XL U40974 ( .A(n34221), .B(n42547), .Y(n44695) );
  XOR2XL U40975 ( .A(n34205), .B(n42547), .Y(n44755) );
  XOR2XL U40976 ( .A(n34245), .B(n36832), .Y(n44817) );
  XOR2XL U40977 ( .A(n34165), .B(n42547), .Y(n44062) );
  XOR2XL U40978 ( .A(n34157), .B(n42547), .Y(n43939) );
  XOR2XL U40979 ( .A(n34181), .B(n42547), .Y(n44124) );
  XOR2XL U40980 ( .A(n34125), .B(n42547), .Y(n43908) );
  XOR2XL U40981 ( .A(n34229), .B(n36832), .Y(n44844) );
  XOR2XL U40982 ( .A(n34149), .B(n42547), .Y(n43970) );
  XOR2XL U40983 ( .A(n34173), .B(n42547), .Y(n44093) );
  XOR2XL U40984 ( .A(n34213), .B(n42547), .Y(n44664) );
  XOR2XL U40985 ( .A(n34197), .B(n42547), .Y(n44724) );
  XOR2XL U40986 ( .A(n34261), .B(n36832), .Y(n45338) );
  XOR2XL U40987 ( .A(n34253), .B(n36832), .Y(n44875) );
  XOR2XL U40988 ( .A(n34222), .B(n42533), .Y(n44694) );
  XOR2XL U40989 ( .A(n34206), .B(n42536), .Y(n44754) );
  XOR2XL U40990 ( .A(n34246), .B(n42533), .Y(n44816) );
  XOR2XL U40991 ( .A(n34166), .B(n42540), .Y(n44061) );
  XOR2XL U40992 ( .A(n34158), .B(n42535), .Y(n43938) );
  XOR2XL U40993 ( .A(n34182), .B(n42535), .Y(n44123) );
  XOR2XL U40994 ( .A(n34238), .B(n42533), .Y(n44785) );
  XOR2XL U40995 ( .A(n34230), .B(n42535), .Y(n44843) );
  XOR2XL U40996 ( .A(n34310), .B(n42533), .Y(n45456) );
  XOR2XL U40997 ( .A(n34174), .B(n42541), .Y(n44092) );
  XOR2XL U40998 ( .A(n34270), .B(n42533), .Y(n45310) );
  XOR2XL U40999 ( .A(n34150), .B(n42536), .Y(n43969) );
  XOR2XL U41000 ( .A(n34278), .B(n42533), .Y(n45368) );
  XOR2XL U41001 ( .A(n34198), .B(n42539), .Y(n44723) );
  XOR2XL U41002 ( .A(n42471), .B(n34312), .Y(n47311) );
  XOR2XL U41003 ( .A(n42471), .B(n34344), .Y(n47650) );
  XOR2XL U41004 ( .A(n36746), .B(n34372), .Y(n47616) );
  XOR2XL U41005 ( .A(n36744), .B(n34348), .Y(n47638) );
  XOR2XL U41006 ( .A(n36743), .B(n34332), .Y(n47595) );
  XOR2XL U41007 ( .A(n41304), .B(n34348), .Y(n46548) );
  XOR2XL U41008 ( .A(n41305), .B(n34356), .Y(n46493) );
  XOR2XL U41009 ( .A(n41302), .B(n34340), .Y(n46537) );
  XOR2XL U41010 ( .A(n36740), .B(n34356), .Y(n47627) );
  XOR2XL U41011 ( .A(n41300), .B(n34276), .Y(n46369) );
  XOR2XL U41012 ( .A(n41303), .B(n34300), .Y(n46325) );
  XOR2XL U41013 ( .A(n41300), .B(n34268), .Y(n46387) );
  XOR2XL U41014 ( .A(n36742), .B(n34276), .Y(n47351) );
  XOR2XL U41015 ( .A(n41301), .B(n34332), .Y(n46516) );
  XOR2XL U41016 ( .A(n36741), .B(n34340), .Y(n47649) );
  XNOR2XL U41017 ( .A(n36859), .B(n34368), .Y(n46503) );
  XOR2XL U41018 ( .A(n36918), .B(n34364), .Y(n46507) );
  XOR2XL U41019 ( .A(n42470), .B(n34392), .Y(n47686) );
  NOR2X2 U41020 ( .A(n11685), .B(n43718), .Y(n43722) );
  XOR2XL U41021 ( .A(n33444), .B(n36821), .Y(n43718) );
  XOR2XL U41022 ( .A(n33740), .B(n36829), .Y(n44277) );
  XNOR2XL U41023 ( .A(n36747), .B(n34380), .Y(n47656) );
  NOR2XL U41024 ( .A(n10555), .B(n46171), .Y(net212726) );
  XOR2XL U41025 ( .A(n33761), .B(n36778), .Y(n46171) );
  XOR2XL U41026 ( .A(n36741), .B(n33508), .Y(n47093) );
  XOR2XL U41027 ( .A(n41303), .B(n33492), .Y(n45813) );
  XOR2XL U41028 ( .A(n36743), .B(n33492), .Y(n47108) );
  XOR2XL U41029 ( .A(n36773), .B(n33841), .Y(n47233) );
  XOR2XL U41030 ( .A(n41305), .B(n33444), .Y(n45848) );
  XOR2XL U41031 ( .A(n33841), .B(n36782), .Y(n46138) );
  XOR2XL U41032 ( .A(n36767), .B(n33633), .Y(n46950) );
  NOR2XL U41033 ( .A(n12292), .B(n47088), .Y(n47092) );
  XOR2XL U41034 ( .A(n36768), .B(n33521), .Y(n47088) );
  XOR2XL U41035 ( .A(n36774), .B(n33529), .Y(n47083) );
  XOR2XL U41036 ( .A(n33633), .B(n36782), .Y(n45748) );
  NOR2XL U41037 ( .A(n12711), .B(n45758), .Y(n45762) );
  XOR2XL U41038 ( .A(n33617), .B(n36778), .Y(n45758) );
  NOR2XL U41039 ( .A(n12703), .B(n45778), .Y(n45782) );
  XOR2XL U41040 ( .A(n41305), .B(n33572), .Y(n45778) );
  NOR2XL U41041 ( .A(n12535), .B(n43629), .Y(net216047) );
  XOR2XL U41042 ( .A(n33884), .B(n36830), .Y(n43629) );
  XOR2XL U41043 ( .A(n41302), .B(n33508), .Y(n45803) );
  NOR2X2 U41044 ( .A(n12493), .B(n43223), .Y(n43227) );
  XOR2XL U41045 ( .A(n33556), .B(n36824), .Y(n44547) );
  XOR2XL U41046 ( .A(n33756), .B(n36828), .Y(n44314) );
  XOR2XL U41047 ( .A(n33492), .B(n36829), .Y(n43691) );
  NOR2XL U41048 ( .A(n10554), .B(n46178), .Y(net212711) );
  XOR2XL U41049 ( .A(n33753), .B(n36783), .Y(n46178) );
  XOR2XL U41050 ( .A(n33540), .B(n36828), .Y(n43809) );
  XOR2XL U41051 ( .A(n33860), .B(n36828), .Y(n43573) );
  XOR2XL U41052 ( .A(n33948), .B(n36827), .Y(n44223) );
  XOR2XL U41053 ( .A(n33745), .B(n36784), .Y(n45654) );
  XOR2XL U41054 ( .A(n41300), .B(n33732), .Y(n45623) );
  XOR2XL U41055 ( .A(n33428), .B(n36830), .Y(n43736) );
  XOR2XL U41056 ( .A(n36771), .B(n34009), .Y(n47025) );
  XOR2XL U41057 ( .A(n41305), .B(n33700), .Y(n46169) );
  XOR2XL U41058 ( .A(n33852), .B(n36829), .Y(n43550) );
  XOR2XL U41059 ( .A(n36918), .B(n33556), .Y(n45768) );
  XOR2XL U41060 ( .A(n36770), .B(n33577), .Y(n46915) );
  XOR2XL U41061 ( .A(n41302), .B(n33804), .Y(n47189) );
  XOR2XL U41062 ( .A(n33657), .B(n36786), .Y(n45743) );
  XOR2XL U41063 ( .A(n33812), .B(n36828), .Y(n43673) );
  XOR2XL U41064 ( .A(n33857), .B(n36777), .Y(n46128) );
  XOR2XL U41065 ( .A(n36748), .B(n33812), .Y(n47139) );
  XOR2XL U41066 ( .A(n36741), .B(n33820), .Y(n47144) );
  NOR2XL U41067 ( .A(n12303), .B(n46965), .Y(net211657) );
  XOR2XL U41068 ( .A(n36772), .B(n33657), .Y(n46965) );
  XOR2XL U41069 ( .A(n33452), .B(n36831), .Y(n43709) );
  XOR2XL U41070 ( .A(n36918), .B(n33428), .Y(n45838) );
  XOR2XL U41071 ( .A(n33836), .B(n36830), .Y(n43656) );
  XOR2XL U41072 ( .A(n33580), .B(n36822), .Y(n44556) );
  XOR2XL U41073 ( .A(n33516), .B(n36828), .Y(n43773) );
  XOR2XL U41074 ( .A(n33596), .B(n36823), .Y(n44512) );
  XOR2XL U41075 ( .A(n33385), .B(n36772), .Y(n46759) );
  XOR2XL U41076 ( .A(n36736), .B(n33930), .Y(n47238) );
  XOR2XL U41077 ( .A(n36742), .B(n33548), .Y(n47073) );
  XOR2XL U41078 ( .A(n33825), .B(n36786), .Y(n46158) );
  XOR2XL U41079 ( .A(n33564), .B(n36829), .Y(n44538) );
  XOR2XL U41080 ( .A(n33436), .B(n36827), .Y(n43727) );
  XOR2XL U41081 ( .A(n36765), .B(n33369), .Y(n46754) );
  XOR2XL U41082 ( .A(n33649), .B(n36786), .Y(n45738) );
  NOR2X2 U41083 ( .A(n12280), .B(n46719), .Y(n46723) );
  XOR2XL U41084 ( .A(n36768), .B(n33393), .Y(n46719) );
  XOR2XL U41085 ( .A(n36774), .B(n33785), .Y(n47204) );
  NOR2XL U41086 ( .A(n10243), .B(n47113), .Y(n47117) );
  XOR2XL U41087 ( .A(n36746), .B(n33476), .Y(n47113) );
  XOR2XL U41088 ( .A(n36774), .B(n33905), .Y(n47897) );
  XOR2XL U41089 ( .A(n33468), .B(n36827), .Y(n43750) );
  NOR2X2 U41090 ( .A(n43205), .B(net214729), .Y(n43209) );
  XOR2XL U41091 ( .A(n33396), .B(n36828), .Y(n43205) );
  XOR2XL U41092 ( .A(n33513), .B(n36784), .Y(n45798) );
  XOR2XL U41093 ( .A(n33601), .B(n36784), .Y(n45728) );
  XOR2XL U41094 ( .A(n36773), .B(n33649), .Y(n46966) );
  XOR2XL U41095 ( .A(n33353), .B(n36784), .Y(n45930) );
  XOR2XL U41096 ( .A(n41300), .B(n33500), .Y(n45808) );
  XOR2XL U41097 ( .A(n36733), .B(n33866), .Y(n47223) );
  XOR2XL U41098 ( .A(n36766), .B(n33849), .Y(n47228) );
  XOR2XL U41099 ( .A(n33369), .B(n36782), .Y(n45895) );
  XOR2XL U41100 ( .A(n33377), .B(n36783), .Y(n46749) );
  XOR2XL U41101 ( .A(n36765), .B(n34105), .Y(n47557) );
  NOR2XL U41102 ( .A(n10529), .B(n45858), .Y(net213125) );
  XOR2XL U41103 ( .A(n41302), .B(n33468), .Y(n45858) );
  NOR2XL U41104 ( .A(n10853), .B(n47217), .Y(net211246) );
  XOR2XL U41105 ( .A(n36772), .B(n33753), .Y(n47217) );
  XOR2XL U41106 ( .A(n36736), .B(n33674), .Y(n46955) );
  XOR2XL U41107 ( .A(n36740), .B(n33420), .Y(n46704) );
  NOR2XL U41108 ( .A(n12063), .B(n45639), .Y(n45643) );
  XOR2XL U41109 ( .A(n33785), .B(n36785), .Y(n45639) );
  XOR2XL U41110 ( .A(n36733), .B(n33738), .Y(n47159) );
  XOR2XL U41111 ( .A(n36740), .B(n33452), .Y(n47063) );
  NOR2XL U41112 ( .A(n12151), .B(n45753), .Y(n45757) );
  XOR2XL U41113 ( .A(n33641), .B(n36784), .Y(n45753) );
  XOR2XL U41114 ( .A(n41303), .B(n33460), .Y(n45859) );
  XOR2XL U41115 ( .A(n33484), .B(n36827), .Y(n43764) );
  NOR2XL U41116 ( .A(n12024), .B(n47128), .Y(n47132) );
  XOR2XL U41117 ( .A(n41302), .B(n33476), .Y(n47128) );
  XOR2XL U41118 ( .A(n36771), .B(n33617), .Y(n46935) );
  XOR2XL U41119 ( .A(n33585), .B(n36786), .Y(n45717) );
  NOR2X2 U41120 ( .A(n11051), .B(n46744), .Y(n46748) );
  XOR2XL U41121 ( .A(n36766), .B(n33361), .Y(n46744) );
  XOR2XL U41122 ( .A(n33364), .B(n36823), .Y(n43294) );
  XOR2XL U41123 ( .A(n33668), .B(n36830), .Y(n44480) );
  XOR2XL U41124 ( .A(n33377), .B(n36770), .Y(n46769) );
  XOR2XL U41125 ( .A(n33508), .B(n36829), .Y(n43700) );
  XOR2XL U41126 ( .A(n33793), .B(n36774), .Y(n47194) );
  XOR2XL U41127 ( .A(n33380), .B(n36823), .Y(n43267) );
  XOR2XL U41128 ( .A(n33889), .B(n36786), .Y(n46118) );
  XOR2XL U41129 ( .A(n33665), .B(n36765), .Y(n46972) );
  XOR2XL U41130 ( .A(n33524), .B(n36831), .Y(n43782) );
  NOR2XL U41131 ( .A(n12342), .B(n47012), .Y(n47016) );
  XOR2XL U41132 ( .A(n36767), .B(n34041), .Y(n47012) );
  NOR2X2 U41133 ( .A(n11710), .B(n44565), .Y(n44569) );
  XOR2XL U41134 ( .A(n33572), .B(n36830), .Y(n44565) );
  NOR2XL U41135 ( .A(n11094), .B(n46940), .Y(n46944) );
  XOR2XL U41136 ( .A(n36772), .B(n33625), .Y(n46940) );
  XOR2XL U41137 ( .A(n36748), .B(n33564), .Y(n46905) );
  XOR2XL U41138 ( .A(n41302), .B(n33436), .Y(n45843) );
  XOR2XL U41139 ( .A(n41301), .B(n33548), .Y(n45823) );
  XOR2XL U41140 ( .A(n36746), .B(n33692), .Y(n47164) );
  XOR2XL U41141 ( .A(n36765), .B(n33513), .Y(n47098) );
  XOR2XL U41142 ( .A(n36766), .B(n33833), .Y(n47134) );
  XOR2XL U41143 ( .A(n33849), .B(n36785), .Y(n46143) );
  NOR2XL U41144 ( .A(n10543), .B(n45763), .Y(n45767) );
  XOR2XL U41145 ( .A(n33625), .B(n36780), .Y(n45763) );
  XOR2XL U41146 ( .A(n36734), .B(n33610), .Y(n46925) );
  XOR2XL U41147 ( .A(n36768), .B(n33593), .Y(n47848) );
  XOR2XL U41148 ( .A(n36768), .B(n33913), .Y(n47902) );
  XOR2XL U41149 ( .A(n41304), .B(n33420), .Y(n45910) );
  XOR2XL U41150 ( .A(n33385), .B(n36785), .Y(n46764) );
  XOR2XL U41151 ( .A(n36743), .B(n34060), .Y(n46992) );
  XOR2XL U41152 ( .A(n41302), .B(n33940), .Y(n45695) );
  XOR2XL U41153 ( .A(n33708), .B(n36831), .Y(n44261) );
  XOR2XL U41154 ( .A(n36747), .B(n33724), .Y(n47877) );
  NOR2XL U41155 ( .A(n11115), .B(n47184), .Y(n47188) );
  XOR2XL U41156 ( .A(n36747), .B(n33804), .Y(n47184) );
  XOR2XL U41157 ( .A(n33868), .B(n36831), .Y(n43564) );
  XOR2XL U41158 ( .A(n36744), .B(n33436), .Y(n47058) );
  XOR2XL U41159 ( .A(n36768), .B(n33641), .Y(n46945) );
  XOR2XL U41160 ( .A(n33684), .B(n36827), .Y(n44238) );
  NOR2XL U41161 ( .A(n47248), .B(net209249), .Y(n47252) );
  XOR2XL U41162 ( .A(n36772), .B(n33881), .Y(n47248) );
  NOR2XL U41163 ( .A(n47215), .B(net209242), .Y(net211256) );
  XOR2XL U41164 ( .A(n36771), .B(n33769), .Y(n47215) );
  XOR2XL U41165 ( .A(n36747), .B(n33428), .Y(n47053) );
  XOR2XL U41166 ( .A(n33873), .B(n36777), .Y(n46113) );
  XOR2XL U41167 ( .A(n33420), .B(n36831), .Y(n43214) );
  XOR2XL U41168 ( .A(n41302), .B(n33484), .Y(n45864) );
  XOR2XL U41169 ( .A(n33388), .B(n36829), .Y(n43276) );
  XOR2XL U41170 ( .A(n36774), .B(n33777), .Y(n47209) );
  XOR2XL U41171 ( .A(n34260), .B(n42637), .Y(n44857) );
  XNOR2XL U41172 ( .A(n36837), .B(n33298), .Y(n45948) );
  XNOR2XL U41173 ( .A(n36845), .B(n33346), .Y(n45938) );
  XNOR2XL U41174 ( .A(n33370), .B(n36725), .Y(n43288) );
  XOR2XL U41175 ( .A(n36744), .B(n34124), .Y(n47571) );
  XOR2XL U41176 ( .A(n36714), .B(n34125), .Y(n47569) );
  XOR2XL U41177 ( .A(n36735), .B(n34122), .Y(n47573) );
  XOR2XL U41178 ( .A(n36771), .B(n34121), .Y(n47572) );
  XNOR2XL U41179 ( .A(n36736), .B(n33338), .Y(n47925) );
  XOR2XL U41180 ( .A(n36797), .B(n34126), .Y(n47568) );
  NOR2XL U41181 ( .A(n12287), .B(n47133), .Y(net211348) );
  XOR2XL U41182 ( .A(n36742), .B(n33468), .Y(n47133) );
  XOR2XL U41183 ( .A(n33340), .B(n36828), .Y(n43232) );
  NOR2X2 U41184 ( .A(n11668), .B(n43303), .Y(n43307) );
  XOR2XL U41185 ( .A(n33324), .B(n36828), .Y(n43303) );
  XOR2XL U41186 ( .A(n36734), .B(n33322), .Y(n46729) );
  XOR2XL U41187 ( .A(n36770), .B(n33329), .Y(n47917) );
  XOR2XL U41188 ( .A(n36772), .B(n33337), .Y(n47922) );
  XOR2XL U41189 ( .A(n33361), .B(n36778), .Y(n45900) );
  XOR2XL U41190 ( .A(n33321), .B(n36776), .Y(n45953) );
  NOR2XL U41191 ( .A(n10233), .B(n46724), .Y(n46728) );
  XOR2XL U41192 ( .A(n36735), .B(n33314), .Y(n46724) );
  XOR2XL U41193 ( .A(n33372), .B(n36830), .Y(n43285) );
  XOR2XL U41194 ( .A(n33356), .B(n36821), .Y(n43250) );
  XOR2XL U41195 ( .A(n33300), .B(n36831), .Y(n43321) );
  XOR2XL U41196 ( .A(n36735), .B(n33354), .Y(n46774) );
  NOR2XL U41197 ( .A(n11073), .B(n47123), .Y(n47127) );
  XOR2XL U41198 ( .A(n36744), .B(n33484), .Y(n47123) );
  NOR2XL U41199 ( .A(n11075), .B(n47103), .Y(n47107) );
  XOR2XL U41200 ( .A(n36740), .B(n33500), .Y(n47103) );
  XOR2XL U41201 ( .A(n33316), .B(n36821), .Y(n43312) );
  XOR2XL U41202 ( .A(n33329), .B(n36779), .Y(n45925) );
  NOR2XL U41203 ( .A(n11046), .B(n46734), .Y(n46738) );
  XOR2XL U41204 ( .A(n36742), .B(n33308), .Y(n46734) );
  XNOR2XL U41205 ( .A(n36841), .B(n33234), .Y(n45988) );
  XNOR2XL U41206 ( .A(n33313), .B(n36785), .Y(n22879) );
  XNOR2XL U41207 ( .A(n33314), .B(n36844), .Y(n22880) );
  NOR2XL U41208 ( .A(n11041), .B(n46686), .Y(net211997) );
  XOR2XL U41209 ( .A(n36747), .B(n33292), .Y(n46686) );
  XOR2XL U41210 ( .A(n36771), .B(n33265), .Y(n46688) );
  XOR2XL U41211 ( .A(n33217), .B(n36777), .Y(n45880) );
  XOR2XL U41212 ( .A(n33228), .B(n36827), .Y(n43335) );
  XOR2XL U41213 ( .A(n36765), .B(n33257), .Y(n46675) );
  XOR2XL U41214 ( .A(n36774), .B(n33225), .Y(n46895) );
  XOR2XL U41215 ( .A(n36772), .B(n33273), .Y(n46685) );
  XOR2XL U41216 ( .A(n36774), .B(n33209), .Y(n46885) );
  XOR2XL U41217 ( .A(n33260), .B(n36829), .Y(n43177) );
  XOR2XL U41218 ( .A(n33281), .B(n36782), .Y(n45969) );
  XOR2XL U41219 ( .A(n33249), .B(n36777), .Y(n45959) );
  XOR2XL U41220 ( .A(n36774), .B(n33249), .Y(n46680) );
  XOR2XL U41221 ( .A(n36768), .B(n33241), .Y(n47932) );
  XOR2XL U41222 ( .A(n33284), .B(n36823), .Y(n43168) );
  XNOR2XL U41223 ( .A(n36843), .B(n33154), .Y(n46038) );
  XNOR2XL U41224 ( .A(n36736), .B(n33194), .Y(n46863) );
  XNOR2XL U41225 ( .A(n36733), .B(n33178), .Y(n46873) );
  XOR2XL U41226 ( .A(n33129), .B(n36786), .Y(n46015) );
  NOR2XL U41227 ( .A(n11029), .B(n46860), .Y(n46864) );
  XOR2XL U41228 ( .A(n36768), .B(n33193), .Y(n46860) );
  XOR2XL U41229 ( .A(n33196), .B(n36824), .Y(n43369) );
  XOR2XL U41230 ( .A(n33145), .B(n36784), .Y(n46040) );
  XOR2XL U41231 ( .A(n36767), .B(n33145), .Y(n46784) );
  XOR2XL U41232 ( .A(n36750), .B(n33180), .Y(n46870) );
  XOR2XL U41233 ( .A(n33172), .B(n36824), .Y(n43396) );
  XOR2XL U41234 ( .A(n41301), .B(n33188), .Y(n45870) );
  XOR2XL U41235 ( .A(n33164), .B(n36828), .Y(n43087) );
  XOR2XL U41236 ( .A(n36743), .B(n33164), .Y(n46799) );
  XNOR2XL U41237 ( .A(n36840), .B(n33114), .Y(n46013) );
  XNOR2XL U41238 ( .A(n36847), .B(n33106), .Y(n46023) );
  XNOR2XL U41239 ( .A(n36838), .B(n33122), .Y(n46028) );
  XNOR2XL U41240 ( .A(n36736), .B(n33074), .Y(n47940) );
  XOR2XL U41241 ( .A(n33108), .B(n36827), .Y(n43131) );
  XOR2XL U41242 ( .A(n33116), .B(n36823), .Y(n43150) );
  XOR2XL U41243 ( .A(n33137), .B(n36786), .Y(n46045) );
  XOR2XL U41244 ( .A(n33121), .B(n36785), .Y(n46025) );
  XOR2XL U41245 ( .A(n33105), .B(n36786), .Y(n46020) );
  XOR2XL U41246 ( .A(n33124), .B(n36828), .Y(n43122) );
  XOR2XL U41247 ( .A(n36765), .B(n33073), .Y(n47937) );
  XOR2XL U41248 ( .A(n36764), .B(n33129), .Y(n46809) );
  NOR2XL U41249 ( .A(n11217), .B(n46829), .Y(n46833) );
  XOR2XL U41250 ( .A(n36733), .B(n33098), .Y(n46829) );
  XOR2XL U41251 ( .A(n36767), .B(n33113), .Y(n47829) );
  XOR2XL U41252 ( .A(n33113), .B(n36783), .Y(n46010) );
  XOR2XL U41253 ( .A(n36773), .B(n33081), .Y(n47942) );
  XOR2XL U41254 ( .A(n33148), .B(n36823), .Y(n43104) );
  XOR2XL U41255 ( .A(n33089), .B(n36783), .Y(n46000) );
  XOR2XL U41256 ( .A(n33132), .B(n36830), .Y(n43136) );
  XOR2XL U41257 ( .A(n33081), .B(n36779), .Y(n46005) );
  XOR2XL U41258 ( .A(n33100), .B(n36822), .Y(n43059) );
  XOR2XL U41259 ( .A(n36735), .B(n33090), .Y(n46834) );
  XOR2XL U41260 ( .A(n33092), .B(n36825), .Y(n43068) );
  XOR2XL U41261 ( .A(n33097), .B(n36784), .Y(n45995) );
  XNOR2XL U41262 ( .A(n36734), .B(n33010), .Y(net211968) );
  XNOR2XL U41263 ( .A(n36736), .B(n33026), .Y(n46693) );
  XNOR2XL U41264 ( .A(n36734), .B(n33050), .Y(n46842) );
  XNOR2XL U41265 ( .A(n36735), .B(n33042), .Y(n46847) );
  XOR2XL U41266 ( .A(n33065), .B(n36785), .Y(n46051) );
  XOR2XL U41267 ( .A(n41303), .B(n33044), .Y(n46050) );
  XOR2XL U41268 ( .A(n33044), .B(n36823), .Y(n43082) );
  NOR2XL U41269 ( .A(n9676), .B(net266151), .Y(n47952) );
  XOR2XL U41270 ( .A(n33057), .B(n36782), .Y(n46053) );
  XOR2XL U41271 ( .A(n33060), .B(n36823), .Y(n43077) );
  XOR2XL U41272 ( .A(n41305), .B(n33052), .Y(n46052) );
  XOR2XL U41273 ( .A(n33012), .B(n36821), .Y(n43408) );
  XOR2XL U41274 ( .A(n36768), .B(n33009), .Y(n46696) );
  XOR2XL U41275 ( .A(n33009), .B(n36785), .Y(n46069) );
  XOR2XL U41276 ( .A(n36767), .B(n32993), .Y(n46698) );
  XOR2XL U41277 ( .A(n33001), .B(n36782), .Y(n46074) );
  NOR2XL U41278 ( .A(n10997), .B(n46697), .Y(net211962) );
  XOR2XL U41279 ( .A(n36771), .B(n33001), .Y(n46697) );
  XOR2XL U41280 ( .A(n36765), .B(n33017), .Y(n46695) );
  XOR2XL U41281 ( .A(n36736), .B(n33066), .Y(n46819) );
  XOR2XL U41282 ( .A(n33017), .B(n36780), .Y(n46064) );
  XOR2XL U41283 ( .A(n33073), .B(n36776), .Y(n45990) );
  XOR2XL U41284 ( .A(n33020), .B(n36827), .Y(n43407) );
  XOR2XL U41285 ( .A(n36765), .B(n33025), .Y(n46690) );
  XOR2XL U41286 ( .A(n33025), .B(n36776), .Y(n46059) );
  XOR2XL U41287 ( .A(n36743), .B(n33036), .Y(n46689) );
  XOR2XL U41288 ( .A(n36747), .B(n33044), .Y(n46844) );
  XOR2XL U41289 ( .A(n33084), .B(n36831), .Y(n43049) );
  XOR2XL U41290 ( .A(n41300), .B(n33036), .Y(n46054) );
  XOR2XL U41291 ( .A(n33052), .B(n36822), .Y(n43141) );
  NOR2XL U41292 ( .A(n10272), .B(n46824), .Y(n46828) );
  XOR2XL U41293 ( .A(n36733), .B(n33058), .Y(n46824) );
  XOR2XL U41294 ( .A(n33049), .B(n36770), .Y(n46839) );
  XOR2XL U41295 ( .A(n33068), .B(n36829), .Y(n44626) );
  XNOR2XL U41296 ( .A(n32850), .B(n42568), .Y(net216320) );
  XNOR2XL U41297 ( .A(n32986), .B(n42567), .Y(n43426) );
  XNOR2XL U41298 ( .A(n32890), .B(n42568), .Y(net216347) );
  XNOR2XL U41299 ( .A(n32978), .B(n42567), .Y(n43421) );
  XNOR2XL U41300 ( .A(n32858), .B(n42565), .Y(net212155) );
  XNOR2XL U41301 ( .A(n32962), .B(n42567), .Y(n43471) );
  XNOR2XL U41302 ( .A(n32930), .B(n42567), .Y(n43451) );
  XNOR2XL U41303 ( .A(n32898), .B(n42567), .Y(net216365) );
  XNOR2XL U41304 ( .A(n36845), .B(n32922), .Y(n47756) );
  XNOR2XL U41305 ( .A(n36844), .B(n32850), .Y(n46631) );
  XNOR2XL U41306 ( .A(n36733), .B(n32986), .Y(n46702) );
  XNOR2XL U41307 ( .A(n36733), .B(n32906), .Y(net212185) );
  XNOR2XL U41308 ( .A(n36733), .B(n32970), .Y(net211794) );
  XNOR2XL U41309 ( .A(n32906), .B(n42567), .Y(n43480) );
  XNOR2XL U41310 ( .A(n33002), .B(n42567), .Y(n43431) );
  XNOR2XL U41311 ( .A(n36733), .B(n32890), .Y(net212175) );
  XNOR2XL U41312 ( .A(n32938), .B(n42567), .Y(net216428) );
  XNOR2XL U41313 ( .A(n36736), .B(n32874), .Y(net212160) );
  XNOR2XL U41314 ( .A(n36847), .B(n32986), .Y(n47795) );
  XNOR2XL U41315 ( .A(n32858), .B(n36846), .Y(n46613) );
  XNOR2XL U41316 ( .A(n32922), .B(n42567), .Y(n43445) );
  XNOR2XL U41317 ( .A(n36840), .B(n32938), .Y(n46083) );
  XNOR2XL U41318 ( .A(n32970), .B(n42567), .Y(n43460) );
  XNOR2XL U41319 ( .A(n32914), .B(n42567), .Y(n43440) );
  XNOR2XL U41320 ( .A(n36734), .B(n32882), .Y(net212170) );
  XNOR2XL U41321 ( .A(n32874), .B(n42568), .Y(net216329) );
  XNOR2XL U41322 ( .A(n32866), .B(n42568), .Y(net216338) );
  XNOR2XL U41323 ( .A(n36735), .B(n32962), .Y(n46852) );
  XNOR2XL U41324 ( .A(n36734), .B(n32898), .Y(n46621) );
  XNOR2XL U41325 ( .A(n36736), .B(n32866), .Y(net212165) );
  XNOR2XL U41326 ( .A(n36735), .B(n32850), .Y(net212195) );
  XNOR2XL U41327 ( .A(n36735), .B(n32834), .Y(n46637) );
  OAI211XL U41328 ( .A0(n41808), .A1(n42816), .B0(n19126), .C0(n49568), .Y(
        n36548) );
  OA22XL U41329 ( .A0(net262532), .A1(n41810), .B0(n41809), .B1(net218800),
        .Y(n19126) );
  INVX1 U41330 ( .A(n19128), .Y(n49568) );
  OAI211XL U41331 ( .A0(n42066), .A1(n42816), .B0(n19114), .C0(n49569), .Y(
        n36544) );
  OA22XL U41332 ( .A0(net262532), .A1(n42068), .B0(n42067), .B1(net218752),
        .Y(n19114) );
  INVX1 U41333 ( .A(n19116), .Y(n49569) );
  OAI211XL U41334 ( .A0(n33708), .A1(n42754), .B0(n17053), .C0(n17054), .Y(
        n35857) );
  OA22XL U41335 ( .A0(net261924), .A1(n33692), .B0(n33700), .B1(n40148), .Y(
        n17053) );
  OAI211XL U41336 ( .A0(n33692), .A1(n42756), .B0(n17005), .C0(n17006), .Y(
        n35841) );
  OA22XL U41337 ( .A0(net261943), .A1(n33676), .B0(n33684), .B1(n40147), .Y(
        n17005) );
  OAI211XL U41338 ( .A0(n33684), .A1(n42757), .B0(n16981), .C0(n16982), .Y(
        n35833) );
  OA22XL U41339 ( .A0(net261943), .A1(n33668), .B0(n33676), .B1(n40146), .Y(
        n16981) );
  OAI211XL U41340 ( .A0(n33676), .A1(n42758), .B0(n16957), .C0(n16958), .Y(
        n35825) );
  OA22XL U41341 ( .A0(net261943), .A1(n33660), .B0(n33668), .B1(n40146), .Y(
        n16957) );
  OAI211XL U41342 ( .A0(n33668), .A1(n42759), .B0(n16933), .C0(n16934), .Y(
        n35817) );
  OA22XL U41343 ( .A0(net218446), .A1(n33652), .B0(n33660), .B1(n40145), .Y(
        n16933) );
  OAI211XL U41344 ( .A0(n33660), .A1(n42761), .B0(n16909), .C0(n16910), .Y(
        n35809) );
  OA22XL U41345 ( .A0(net218480), .A1(n33644), .B0(n33652), .B1(n40145), .Y(
        n16909) );
  OAI211XL U41346 ( .A0(n33484), .A1(n42786), .B0(n16381), .C0(n16382), .Y(
        n35633) );
  OA22XL U41347 ( .A0(net262152), .A1(n33468), .B0(n33476), .B1(n40136), .Y(
        n16381) );
  OAI211XL U41348 ( .A0(n33476), .A1(n42787), .B0(n16357), .C0(n16358), .Y(
        n35625) );
  OA22XL U41349 ( .A0(net262171), .A1(n33460), .B0(n33468), .B1(n40135), .Y(
        n16357) );
  OAI211XL U41350 ( .A0(n33468), .A1(n42788), .B0(n16333), .C0(n16334), .Y(
        n35617) );
  OA22XL U41351 ( .A0(net262171), .A1(n33452), .B0(n33460), .B1(n40135), .Y(
        n16333) );
  OAI211XL U41352 ( .A0(n33020), .A1(n42981), .B0(n14989), .C0(n14990), .Y(
        n35169) );
  OA22XL U41353 ( .A0(net263995), .A1(n33004), .B0(n33012), .B1(n40040), .Y(
        n14989) );
  OAI211XL U41354 ( .A0(n34066), .A1(n42799), .B0(n18127), .C0(n18128), .Y(
        n36215) );
  OA22XL U41355 ( .A0(net262893), .A1(n34050), .B0(n34058), .B1(net218670),
        .Y(n18127) );
  OAI211XL U41356 ( .A0(n34058), .A1(n42800), .B0(n18103), .C0(n18104), .Y(
        n36207) );
  OA22XL U41357 ( .A0(net262893), .A1(n34042), .B0(n34050), .B1(net218832),
        .Y(n18103) );
  OAI211XL U41358 ( .A0(n34018), .A1(n42806), .B0(n17983), .C0(n17984), .Y(
        n36167) );
  OA22XL U41359 ( .A0(net262665), .A1(n34002), .B0(n34010), .B1(n40111), .Y(
        n17983) );
  OAI211XL U41360 ( .A0(n34010), .A1(n42807), .B0(n17959), .C0(n17960), .Y(
        n36159) );
  OA22XL U41361 ( .A0(net218442), .A1(n33994), .B0(n34002), .B1(n40111), .Y(
        n17959) );
  OAI211XL U41362 ( .A0(n33706), .A1(n42754), .B0(n17047), .C0(n17048), .Y(
        n35855) );
  OA22XL U41363 ( .A0(net261924), .A1(n33690), .B0(n33698), .B1(n40148), .Y(
        n17047) );
  OAI211XL U41364 ( .A0(n33690), .A1(n42756), .B0(n16999), .C0(n17000), .Y(
        n35839) );
  OA22XL U41365 ( .A0(net261943), .A1(n33674), .B0(n33682), .B1(n40147), .Y(
        n16999) );
  OAI211XL U41366 ( .A0(n33682), .A1(n42757), .B0(n16975), .C0(n16976), .Y(
        n35831) );
  OA22XL U41367 ( .A0(net261943), .A1(n33666), .B0(n33674), .B1(n40146), .Y(
        n16975) );
  OAI211XL U41368 ( .A0(n33674), .A1(n42759), .B0(n16951), .C0(n16952), .Y(
        n35823) );
  OA22XL U41369 ( .A0(net218440), .A1(n33658), .B0(n33666), .B1(n40146), .Y(
        n16951) );
  OAI211XL U41370 ( .A0(n33666), .A1(n42760), .B0(n16927), .C0(n16928), .Y(
        n35815) );
  OA22XL U41371 ( .A0(net218438), .A1(n33650), .B0(n33658), .B1(n40145), .Y(
        n16927) );
  OAI211XL U41372 ( .A0(n33658), .A1(n42761), .B0(n16903), .C0(n16904), .Y(
        n35807) );
  OA22XL U41373 ( .A0(net218446), .A1(n33642), .B0(n33650), .B1(n40145), .Y(
        n16903) );
  OAI211XL U41374 ( .A0(n33570), .A1(n42741), .B0(n16639), .C0(n16640), .Y(
        n35719) );
  OA22XL U41375 ( .A0(net262342), .A1(n33554), .B0(n33562), .B1(n40126), .Y(
        n16639) );
  OAI211XL U41376 ( .A0(n33562), .A1(n42743), .B0(n16615), .C0(n16616), .Y(
        n35711) );
  OA22XL U41377 ( .A0(net262342), .A1(n33546), .B0(n33554), .B1(n40126), .Y(
        n16615) );
  OAI211XL U41378 ( .A0(n33554), .A1(n42744), .B0(n16591), .C0(n16592), .Y(
        n35703) );
  OA22XL U41379 ( .A0(net262342), .A1(n33538), .B0(n33546), .B1(n40125), .Y(
        n16591) );
  OAI211XL U41380 ( .A0(n33490), .A1(n42785), .B0(n16399), .C0(n16400), .Y(
        n35639) );
  OA22XL U41381 ( .A0(net262152), .A1(n33474), .B0(n33482), .B1(n40136), .Y(
        n16399) );
  OAI211XL U41382 ( .A0(n33482), .A1(n42786), .B0(n16375), .C0(n16376), .Y(
        n35631) );
  OA22XL U41383 ( .A0(net262152), .A1(n33466), .B0(n33474), .B1(n40136), .Y(
        n16375) );
  OAI211XL U41384 ( .A0(n33474), .A1(n42787), .B0(n16351), .C0(n16352), .Y(
        n35623) );
  OA22XL U41385 ( .A0(net262171), .A1(n33458), .B0(n33466), .B1(n40135), .Y(
        n16351) );
  OAI211XL U41386 ( .A0(n33466), .A1(n42788), .B0(n16327), .C0(n16328), .Y(
        n35615) );
  OA22XL U41387 ( .A0(net262171), .A1(n33450), .B0(n33458), .B1(n40135), .Y(
        n16327) );
  OAI211XL U41388 ( .A0(n33386), .A1(n42768), .B0(n16087), .C0(n16088), .Y(
        n35535) );
  OA22XL U41389 ( .A0(net263615), .A1(n33370), .B0(n33378), .B1(n40061), .Y(
        n16087) );
  OAI211XL U41390 ( .A0(n33322), .A1(n42777), .B0(n15895), .C0(n15896), .Y(
        n35471) );
  OA22XL U41391 ( .A0(net263672), .A1(n33306), .B0(n33314), .B1(n40065), .Y(
        n15895) );
  OAI211XL U41392 ( .A0(n33314), .A1(n42778), .B0(n15871), .C0(n15872), .Y(
        n35463) );
  OA22XL U41393 ( .A0(net263691), .A1(n33298), .B0(n33306), .B1(n40057), .Y(
        n15871) );
  OAI211XL U41394 ( .A0(n33242), .A1(n42949), .B0(n15655), .C0(n15656), .Y(
        n35391) );
  OA22XL U41395 ( .A0(net218370), .A1(n33226), .B0(n33234), .B1(n40068), .Y(
        n15655) );
  OA22XL U41396 ( .A0(net218524), .A1(n32994), .B0(n33002), .B1(net218866),
        .Y(n14959) );
  OA22XL U41397 ( .A0(net263292), .A1(n42707), .B0(n32402), .B1(n40079), .Y(
        n13159) );
  OA22XL U41398 ( .A0(net263292), .A1(n36907), .B0(n42707), .B1(n40078), .Y(
        n13135) );
  OAI211XL U41399 ( .A0(n33948), .A1(n42848), .B0(n17773), .C0(n17774), .Y(
        n36097) );
  OA22XL U41400 ( .A0(net262741), .A1(n33932), .B0(n33940), .B1(n40108), .Y(
        n17773) );
  OAI211XL U41401 ( .A0(n33940), .A1(n42849), .B0(n17749), .C0(n17750), .Y(
        n36089) );
  OA22XL U41402 ( .A0(net218458), .A1(n33924), .B0(n33932), .B1(n40058), .Y(
        n17749) );
  OAI211XL U41403 ( .A0(n33932), .A1(n42851), .B0(n17725), .C0(n17726), .Y(
        n36081) );
  OA22XL U41404 ( .A0(net218456), .A1(n33916), .B0(n33924), .B1(n40130), .Y(
        n17725) );
  OAI211XL U41405 ( .A0(n33796), .A1(n42838), .B0(n17317), .C0(n17318), .Y(
        n35945) );
  OA22XL U41406 ( .A0(net262095), .A1(n33780), .B0(n33788), .B1(net218870),
        .Y(n17317) );
  OAI211XL U41407 ( .A0(n33788), .A1(n42839), .B0(n17293), .C0(n17294), .Y(
        n35937) );
  OA22XL U41408 ( .A0(net262095), .A1(n33772), .B0(n33780), .B1(n40139), .Y(
        n17293) );
  OAI211XL U41409 ( .A0(n33780), .A1(n42840), .B0(n17269), .C0(n17270), .Y(
        n35929) );
  OA22XL U41410 ( .A0(net262114), .A1(n33764), .B0(n33772), .B1(n40139), .Y(
        n17269) );
  OAI211XL U41411 ( .A0(n34074), .A1(n42830), .B0(n18151), .C0(n18152), .Y(
        n36223) );
  OA22XL U41412 ( .A0(net262874), .A1(n34058), .B0(n34066), .B1(n40102), .Y(
        n18151) );
  OAI211XL U41413 ( .A0(n33978), .A1(n42812), .B0(n17863), .C0(n17864), .Y(
        n36127) );
  OA22XL U41414 ( .A0(net262703), .A1(n33962), .B0(n33970), .B1(n40109), .Y(
        n17863) );
  OAI211XL U41415 ( .A0(n33946), .A1(n42849), .B0(n17767), .C0(n17768), .Y(
        n36095) );
  OA22XL U41416 ( .A0(net262741), .A1(n33930), .B0(n33938), .B1(n40108), .Y(
        n17767) );
  OAI211XL U41417 ( .A0(n33938), .A1(n42850), .B0(n17743), .C0(n17744), .Y(
        n36087) );
  OA22XL U41418 ( .A0(net218476), .A1(n33922), .B0(n33930), .B1(n40058), .Y(
        n17743) );
  OAI211XL U41419 ( .A0(n33930), .A1(n42851), .B0(n17719), .C0(n17720), .Y(
        n36079) );
  OA22XL U41420 ( .A0(net218478), .A1(n33914), .B0(n33922), .B1(n40130), .Y(
        n17719) );
  OAI211XL U41421 ( .A0(n33922), .A1(n42852), .B0(n17695), .C0(n17696), .Y(
        n36071) );
  OA22XL U41422 ( .A0(net262779), .A1(n33906), .B0(n33914), .B1(n40107), .Y(
        n17695) );
  OAI211XL U41423 ( .A0(n33914), .A1(n42853), .B0(n17671), .C0(n17672), .Y(
        n36063) );
  OA22XL U41424 ( .A0(net262779), .A1(n33898), .B0(n33906), .B1(n40107), .Y(
        n17671) );
  OAI211XL U41425 ( .A0(n33850), .A1(n42862), .B0(n17479), .C0(n17480), .Y(
        n35999) );
  OA22XL U41426 ( .A0(net262038), .A1(n33834), .B0(n33842), .B1(n40142), .Y(
        n17479) );
  OAI211XL U41427 ( .A0(n33842), .A1(n42831), .B0(n17455), .C0(n17456), .Y(
        n35991) );
  OA22XL U41428 ( .A0(net262038), .A1(n33826), .B0(n33834), .B1(n40141), .Y(
        n17455) );
  OAI211XL U41429 ( .A0(n33834), .A1(n42832), .B0(n17431), .C0(n17432), .Y(
        n35983) );
  OA22XL U41430 ( .A0(net262057), .A1(n33818), .B0(n33826), .B1(n40141), .Y(
        n17431) );
  OAI211XL U41431 ( .A0(n33826), .A1(n42834), .B0(n17407), .C0(n17408), .Y(
        n35975) );
  OA22XL U41432 ( .A0(net262057), .A1(n33810), .B0(n33818), .B1(n40140), .Y(
        n17407) );
  OAI211XL U41433 ( .A0(n33818), .A1(n42835), .B0(n17383), .C0(n17384), .Y(
        n35967) );
  OA22XL U41434 ( .A0(net218574), .A1(n33802), .B0(n33810), .B1(n40140), .Y(
        n17383) );
  OAI211XL U41435 ( .A0(n33810), .A1(n42836), .B0(n17359), .C0(n17360), .Y(
        n35959) );
  OA22XL U41436 ( .A0(net218458), .A1(n33794), .B0(n33802), .B1(net218842),
        .Y(n17359) );
  OAI211XL U41437 ( .A0(n33802), .A1(n42837), .B0(n17335), .C0(n17336), .Y(
        n35951) );
  OA22XL U41438 ( .A0(net262095), .A1(n33786), .B0(n33794), .B1(net218856),
        .Y(n17335) );
  OAI211XL U41439 ( .A0(n33794), .A1(n42838), .B0(n17311), .C0(n17312), .Y(
        n35943) );
  OA22XL U41440 ( .A0(net262095), .A1(n33778), .B0(n33786), .B1(n40139), .Y(
        n17311) );
  OAI211XL U41441 ( .A0(n33786), .A1(n42839), .B0(n17287), .C0(n17288), .Y(
        n35935) );
  OA22XL U41442 ( .A0(net262095), .A1(n33770), .B0(n33778), .B1(n40139), .Y(
        n17287) );
  OAI211XL U41443 ( .A0(n33778), .A1(n42841), .B0(n17263), .C0(n17264), .Y(
        n35927) );
  OA22XL U41444 ( .A0(net262114), .A1(n33762), .B0(n33770), .B1(n40138), .Y(
        n17263) );
  OAI211XL U41445 ( .A0(n33770), .A1(n42842), .B0(n17239), .C0(n17240), .Y(
        n35919) );
  OA22XL U41446 ( .A0(net218294), .A1(n33754), .B0(n33762), .B1(net218610),
        .Y(n17239) );
  OAI211XL U41447 ( .A0(n33762), .A1(n42843), .B0(n17215), .C0(n17216), .Y(
        n35911) );
  OA22XL U41448 ( .A0(net261867), .A1(n33746), .B0(n33754), .B1(n40151), .Y(
        n17215) );
  OAI211XL U41449 ( .A0(n33754), .A1(n42844), .B0(n17191), .C0(n17192), .Y(
        n35903) );
  OA22XL U41450 ( .A0(net261867), .A1(n33738), .B0(n33746), .B1(n40151), .Y(
        n17191) );
  OAI211XL U41451 ( .A0(n9654), .A1(n9754), .B0(net218294), .C0(n42735), .Y(
        n34517) );
  OAI211XL U41452 ( .A0(n41806), .A1(n42735), .B0(n19174), .C0(n49559), .Y(
        n36564) );
  OA22XL U41453 ( .A0(net262646), .A1(n41808), .B0(n41807), .B1(n40065), .Y(
        n19174) );
  OAI211XL U41454 ( .A0(n33578), .A1(n42740), .B0(n16663), .C0(n16664), .Y(
        n35727) );
  OA22XL U41455 ( .A0(net262323), .A1(n33562), .B0(n33570), .B1(n40127), .Y(
        n16663) );
  XOR2XL U41456 ( .A(n32977), .B(n36783), .Y(n46075) );
  OAI211XL U41457 ( .A0(n32946), .A1(n42991), .B0(n14767), .C0(n14768), .Y(
        n35095) );
  XOR2XL U41458 ( .A(n32868), .B(n36823), .Y(n43493) );
  XOR2XL U41459 ( .A(n32876), .B(n36821), .Y(n43494) );
  OA22XL U41460 ( .A0(net263330), .A1(n34404), .B0(n41798), .B1(n40077), .Y(
        n13040) );
  INVX1 U41461 ( .A(n13042), .Y(n50077) );
  OAI211XL U41462 ( .A0(n41798), .A1(n42815), .B0(n19165), .C0(n49562), .Y(
        n36561) );
  OA22XL U41463 ( .A0(net262513), .A1(n34396), .B0(n34404), .B1(net218754),
        .Y(n19165) );
  OA22XL U41464 ( .A0(net263330), .A1(n34405), .B0(n41800), .B1(n40077), .Y(
        n13037) );
  INVX1 U41465 ( .A(n13039), .Y(n50078) );
  OAI211XL U41466 ( .A0(n41800), .A1(n42823), .B0(n19168), .C0(n49561), .Y(
        n36562) );
  OA22XL U41467 ( .A0(net262513), .A1(n34397), .B0(n34405), .B1(net218750),
        .Y(n19168) );
  OA22XL U41468 ( .A0(net263330), .A1(n34406), .B0(n41803), .B1(n40077), .Y(
        n13034) );
  INVX1 U41469 ( .A(n13036), .Y(n50079) );
  OAI211XL U41470 ( .A0(n41803), .A1(n42831), .B0(n19171), .C0(n49560), .Y(
        n36563) );
  OA22XL U41471 ( .A0(net262589), .A1(n34398), .B0(n34406), .B1(n40115), .Y(
        n19171) );
  OA22XL U41472 ( .A0(net263463), .A1(n41807), .B0(n41806), .B1(n40069), .Y(
        n13031) );
  INVX1 U41473 ( .A(n13033), .Y(n50080) );
  OAI211XL U41474 ( .A0(n41807), .A1(n42815), .B0(n19150), .C0(n49566), .Y(
        n36556) );
  OA22XL U41475 ( .A0(net262532), .A1(n41809), .B0(n41808), .B1(net218768),
        .Y(n19150) );
  OA22XL U41476 ( .A0(net218294), .A1(n34408), .B0(n42057), .B1(net218610),
        .Y(n13028) );
  INVX1 U41477 ( .A(n13030), .Y(n50081) );
  OAI211XL U41478 ( .A0(n42057), .A1(n42863), .B0(n19177), .C0(n49558), .Y(
        n36565) );
  OA22XL U41479 ( .A0(net262931), .A1(n34400), .B0(n34408), .B1(n40100), .Y(
        n19177) );
  OA22XL U41480 ( .A0(net263330), .A1(n34401), .B0(n42059), .B1(net218656),
        .Y(n13049) );
  INVX1 U41481 ( .A(n13051), .Y(n50074) );
  OAI211XL U41482 ( .A0(n42059), .A1(n42815), .B0(n19156), .C0(n49565), .Y(
        n36558) );
  OA22XL U41483 ( .A0(net262532), .A1(n34393), .B0(n34401), .B1(net218756),
        .Y(n19156) );
  OA22XL U41484 ( .A0(net263330), .A1(n34402), .B0(n42062), .B1(net218654),
        .Y(n13046) );
  INVX1 U41485 ( .A(n13048), .Y(n50075) );
  OAI211XL U41486 ( .A0(n42062), .A1(n42815), .B0(n19159), .C0(n49564), .Y(
        n36559) );
  OA22XL U41487 ( .A0(net262532), .A1(n34394), .B0(n34402), .B1(net218866),
        .Y(n19159) );
  OA22XL U41488 ( .A0(net263330), .A1(n42065), .B0(n42064), .B1(n40077), .Y(
        n13043) );
  INVX1 U41489 ( .A(n13045), .Y(n50076) );
  OAI211XL U41490 ( .A0(n42064), .A1(n42815), .B0(n19162), .C0(n49563), .Y(
        n36560) );
  OA22XL U41491 ( .A0(net262532), .A1(n42066), .B0(n42065), .B1(net218866),
        .Y(n19162) );
  OAI211XL U41492 ( .A0(n42065), .A1(n42815), .B0(n19138), .C0(n49567), .Y(
        n36552) );
  OA22XL U41493 ( .A0(net262532), .A1(n42067), .B0(n42066), .B1(net218770),
        .Y(n19138) );
  OAI211XL U41494 ( .A0(n34068), .A1(n42799), .B0(n18133), .C0(n18134), .Y(
        n36217) );
  OA22XL U41495 ( .A0(net262893), .A1(n34052), .B0(n34060), .B1(n40102), .Y(
        n18133) );
  OAI211XL U41496 ( .A0(n34060), .A1(n42800), .B0(n18109), .C0(n18110), .Y(
        n36209) );
  OA22XL U41497 ( .A0(net262893), .A1(n34044), .B0(n34052), .B1(n40124), .Y(
        n18109) );
  OAI211XL U41498 ( .A0(n34052), .A1(n42801), .B0(n18085), .C0(n18086), .Y(
        n36201) );
  OA22XL U41499 ( .A0(net262912), .A1(n34036), .B0(n34044), .B1(net218900),
        .Y(n18085) );
  OAI211XL U41500 ( .A0(n34028), .A1(n42805), .B0(n18013), .C0(n18014), .Y(
        n36177) );
  OA22XL U41501 ( .A0(net262665), .A1(n34012), .B0(n34020), .B1(n40086), .Y(
        n18013) );
  OAI211XL U41502 ( .A0(n34020), .A1(n42806), .B0(n17989), .C0(n17990), .Y(
        n36169) );
  OA22XL U41503 ( .A0(net262665), .A1(n34004), .B0(n34012), .B1(n40072), .Y(
        n17989) );
  OAI211XL U41504 ( .A0(n34012), .A1(n42807), .B0(n17965), .C0(n17966), .Y(
        n36161) );
  OA22XL U41505 ( .A0(net218310), .A1(n33996), .B0(n34004), .B1(n40111), .Y(
        n17965) );
  OAI211XL U41506 ( .A0(n34004), .A1(n42808), .B0(n17941), .C0(n17942), .Y(
        n36153) );
  OA22XL U41507 ( .A0(net218384), .A1(n33988), .B0(n33996), .B1(n40111), .Y(
        n17941) );
  OAI211XL U41508 ( .A0(n33996), .A1(n42809), .B0(n17917), .C0(n17918), .Y(
        n36145) );
  OA22XL U41509 ( .A0(net218314), .A1(n33980), .B0(n33988), .B1(n40110), .Y(
        n17917) );
  OAI211XL U41510 ( .A0(n33732), .A1(n42758), .B0(n17125), .C0(n17126), .Y(
        n35881) );
  OA22XL U41511 ( .A0(net261886), .A1(n33716), .B0(n33724), .B1(n40150), .Y(
        n17125) );
  OAI211XL U41512 ( .A0(n33724), .A1(n42751), .B0(n17101), .C0(n17102), .Y(
        n35873) );
  OA22XL U41513 ( .A0(net261905), .A1(n33708), .B0(n33716), .B1(n40149), .Y(
        n17101) );
  OAI211XL U41514 ( .A0(n33716), .A1(n42752), .B0(n17077), .C0(n17078), .Y(
        n35865) );
  OA22XL U41515 ( .A0(net261905), .A1(n33700), .B0(n33708), .B1(n40149), .Y(
        n17077) );
  OAI211XL U41516 ( .A0(n33644), .A1(n42763), .B0(n16861), .C0(n16862), .Y(
        n35793) );
  OA22XL U41517 ( .A0(net262247), .A1(n33628), .B0(n33636), .B1(n40130), .Y(
        n16861) );
  OAI211XL U41518 ( .A0(n33636), .A1(n42764), .B0(n16837), .C0(n16838), .Y(
        n35785) );
  OA22XL U41519 ( .A0(net262266), .A1(n33620), .B0(n33628), .B1(n40130), .Y(
        n16837) );
  OAI211XL U41520 ( .A0(n33628), .A1(n42765), .B0(n16813), .C0(n16814), .Y(
        n35777) );
  OA22XL U41521 ( .A0(net262266), .A1(n33612), .B0(n33620), .B1(n40129), .Y(
        n16813) );
  OAI211XL U41522 ( .A0(n33620), .A1(n42742), .B0(n16789), .C0(n16790), .Y(
        n35769) );
  OA22XL U41523 ( .A0(net262285), .A1(n33604), .B0(n33612), .B1(n40129), .Y(
        n16789) );
  OAI211XL U41524 ( .A0(n33572), .A1(n42741), .B0(n16645), .C0(n16646), .Y(
        n35721) );
  OA22XL U41525 ( .A0(net262323), .A1(n33556), .B0(n33564), .B1(n40126), .Y(
        n16645) );
  OAI211XL U41526 ( .A0(n33564), .A1(n42742), .B0(n16621), .C0(n16622), .Y(
        n35713) );
  OA22XL U41527 ( .A0(net262342), .A1(n33548), .B0(n33556), .B1(n40126), .Y(
        n16621) );
  OAI211XL U41528 ( .A0(n33556), .A1(n42743), .B0(n16597), .C0(n16598), .Y(
        n35705) );
  OA22XL U41529 ( .A0(net262342), .A1(n33540), .B0(n33548), .B1(n40125), .Y(
        n16597) );
  OAI211XL U41530 ( .A0(n33516), .A1(n42749), .B0(n16477), .C0(n16478), .Y(
        n35665) );
  OA22XL U41531 ( .A0(net262114), .A1(n33500), .B0(n33508), .B1(n40138), .Y(
        n16477) );
  OAI211XL U41532 ( .A0(n33508), .A1(n42790), .B0(n16453), .C0(n16454), .Y(
        n35657) );
  OA22XL U41533 ( .A0(net262133), .A1(n33492), .B0(n33500), .B1(n40137), .Y(
        n16453) );
  OAI211XL U41534 ( .A0(n33500), .A1(n42784), .B0(n16429), .C0(n16430), .Y(
        n35649) );
  OA22XL U41535 ( .A0(net262133), .A1(n33484), .B0(n33492), .B1(n40137), .Y(
        n16429) );
  OAI211XL U41536 ( .A0(n33492), .A1(n42785), .B0(n16405), .C0(n16406), .Y(
        n35641) );
  OA22XL U41537 ( .A0(net262152), .A1(n33476), .B0(n33484), .B1(n40136), .Y(
        n16405) );
  OAI211XL U41538 ( .A0(n33388), .A1(n42767), .B0(n16093), .C0(n16094), .Y(
        n35537) );
  OA22XL U41539 ( .A0(net263596), .A1(n33372), .B0(n33380), .B1(n40061), .Y(
        n16093) );
  OAI211XL U41540 ( .A0(n33380), .A1(n42769), .B0(n16069), .C0(n16070), .Y(
        n35529) );
  OA22XL U41541 ( .A0(net263615), .A1(n33364), .B0(n33372), .B1(n40061), .Y(
        n16069) );
  OAI211XL U41542 ( .A0(n33372), .A1(n42770), .B0(n16045), .C0(n16046), .Y(
        n35521) );
  OA22XL U41543 ( .A0(net263615), .A1(n33356), .B0(n33364), .B1(n40060), .Y(
        n16045) );
  OAI211XL U41544 ( .A0(n33364), .A1(n42771), .B0(n16021), .C0(n16022), .Y(
        n35513) );
  OA22XL U41545 ( .A0(net263634), .A1(n33348), .B0(n33356), .B1(n40060), .Y(
        n16021) );
  OAI211XL U41546 ( .A0(n33356), .A1(n42772), .B0(n15997), .C0(n15998), .Y(
        n35505) );
  OA22XL U41547 ( .A0(net263634), .A1(n33340), .B0(n33348), .B1(n40059), .Y(
        n15997) );
  OAI211XL U41548 ( .A0(n33348), .A1(n42773), .B0(n15973), .C0(n15974), .Y(
        n35497) );
  OA22XL U41549 ( .A0(net263653), .A1(n33332), .B0(n33340), .B1(n40059), .Y(
        n15973) );
  OAI211XL U41550 ( .A0(n33340), .A1(n42774), .B0(n15949), .C0(n15950), .Y(
        n35489) );
  OA22XL U41551 ( .A0(net263653), .A1(n33324), .B0(n33332), .B1(n40058), .Y(
        n15949) );
  OAI211XL U41552 ( .A0(n33332), .A1(n42776), .B0(n15925), .C0(n15926), .Y(
        n35481) );
  OA22XL U41553 ( .A0(net263672), .A1(n33316), .B0(n33324), .B1(n40058), .Y(
        n15925) );
  OAI211XL U41554 ( .A0(n33324), .A1(n42777), .B0(n15901), .C0(n15902), .Y(
        n35473) );
  OA22XL U41555 ( .A0(net263672), .A1(n33308), .B0(n33316), .B1(n40137), .Y(
        n15901) );
  OAI211XL U41556 ( .A0(n33316), .A1(n42778), .B0(n15877), .C0(n15878), .Y(
        n35465) );
  OA22XL U41557 ( .A0(net263672), .A1(n33300), .B0(n33308), .B1(n40138), .Y(
        n15877) );
  OAI211XL U41558 ( .A0(n33308), .A1(n42779), .B0(n15853), .C0(n15854), .Y(
        n35457) );
  OA22XL U41559 ( .A0(net263691), .A1(n33292), .B0(n33300), .B1(n40057), .Y(
        n15853) );
  OAI211XL U41560 ( .A0(n33300), .A1(n42780), .B0(n15829), .C0(n15830), .Y(
        n35449) );
  OA22XL U41561 ( .A0(net263691), .A1(n33284), .B0(n33292), .B1(n40057), .Y(
        n15829) );
  OAI211XL U41562 ( .A0(n33292), .A1(n42781), .B0(n15805), .C0(n15806), .Y(
        n35441) );
  OA22XL U41563 ( .A0(net263710), .A1(n33276), .B0(n33284), .B1(n40056), .Y(
        n15805) );
  OAI211XL U41564 ( .A0(n33260), .A1(n42947), .B0(n15709), .C0(n15710), .Y(
        n35409) );
  OA22XL U41565 ( .A0(net263463), .A1(n33244), .B0(n33252), .B1(n40069), .Y(
        n15709) );
  OAI211XL U41566 ( .A0(n33252), .A1(n42948), .B0(n15685), .C0(n15686), .Y(
        n35401) );
  OA22XL U41567 ( .A0(net218430), .A1(n33236), .B0(n33244), .B1(n40069), .Y(
        n15685) );
  OAI211XL U41568 ( .A0(n33244), .A1(n42949), .B0(n15661), .C0(n15662), .Y(
        n35393) );
  OA22XL U41569 ( .A0(net218538), .A1(n33228), .B0(n33236), .B1(n40068), .Y(
        n15661) );
  OAI211XL U41570 ( .A0(n33236), .A1(n42950), .B0(n15637), .C0(n15638), .Y(
        n35385) );
  OA22XL U41571 ( .A0(net263501), .A1(n33220), .B0(n33228), .B1(n40068), .Y(
        n15637) );
  OAI211XL U41572 ( .A0(n33228), .A1(n42951), .B0(n15613), .C0(n15614), .Y(
        n35377) );
  OA22XL U41573 ( .A0(net263501), .A1(n33212), .B0(n33220), .B1(n40067), .Y(
        n15613) );
  OAI211XL U41574 ( .A0(n33220), .A1(n42952), .B0(n15589), .C0(n15590), .Y(
        n35369) );
  OA22XL U41575 ( .A0(net218308), .A1(n33204), .B0(n33212), .B1(n40067), .Y(
        n15589) );
  OAI211XL U41576 ( .A0(n33212), .A1(n42954), .B0(n15565), .C0(n15566), .Y(
        n35361) );
  OA22XL U41577 ( .A0(net218484), .A1(n33196), .B0(n33204), .B1(n40066), .Y(
        n15565) );
  OAI211XL U41578 ( .A0(n33204), .A1(n42955), .B0(n15541), .C0(n15542), .Y(
        n35353) );
  OA22XL U41579 ( .A0(net218384), .A1(n33188), .B0(n33196), .B1(n40066), .Y(
        n15541) );
  OAI211XL U41580 ( .A0(n33196), .A1(n42956), .B0(n15517), .C0(n15518), .Y(
        n35345) );
  OA22XL U41581 ( .A0(net263539), .A1(n33180), .B0(n33188), .B1(n40065), .Y(
        n15517) );
  OAI211XL U41582 ( .A0(n33188), .A1(n42957), .B0(n15493), .C0(n15494), .Y(
        n35337) );
  OA22XL U41583 ( .A0(net263539), .A1(n33172), .B0(n33180), .B1(n40064), .Y(
        n15493) );
  OAI211XL U41584 ( .A0(n33180), .A1(n42958), .B0(n15469), .C0(n15470), .Y(
        n35329) );
  OA22XL U41585 ( .A0(net263558), .A1(n33164), .B0(n33172), .B1(n40064), .Y(
        n15469) );
  OAI211XL U41586 ( .A0(n33172), .A1(n42959), .B0(n15445), .C0(n15446), .Y(
        n35321) );
  OA22XL U41587 ( .A0(net263558), .A1(n33156), .B0(n33164), .B1(n40063), .Y(
        n15445) );
  OAI211XL U41588 ( .A0(n33132), .A1(n42933), .B0(n15325), .C0(n15326), .Y(
        n35281) );
  OA22XL U41589 ( .A0(net263881), .A1(n33116), .B0(n33124), .B1(n40046), .Y(
        n15325) );
  OAI211XL U41590 ( .A0(n33124), .A1(n42934), .B0(n15301), .C0(n15302), .Y(
        n35273) );
  OA22XL U41591 ( .A0(net263881), .A1(n33108), .B0(n33116), .B1(n40046), .Y(
        n15301) );
  OAI211XL U41592 ( .A0(n33116), .A1(n42935), .B0(n15277), .C0(n15278), .Y(
        n35265) );
  OA22XL U41593 ( .A0(net263900), .A1(n33100), .B0(n33108), .B1(n40045), .Y(
        n15277) );
  OAI211XL U41594 ( .A0(n33108), .A1(n42936), .B0(n15253), .C0(n15254), .Y(
        n35257) );
  OA22XL U41595 ( .A0(net263900), .A1(n33092), .B0(n33100), .B1(n40045), .Y(
        n15253) );
  OAI211XL U41596 ( .A0(n33100), .A1(n42937), .B0(n15229), .C0(n15230), .Y(
        n35249) );
  OA22XL U41597 ( .A0(net263900), .A1(n33084), .B0(n33092), .B1(n40044), .Y(
        n15229) );
  OAI211XL U41598 ( .A0(n33092), .A1(n42939), .B0(n15205), .C0(n15206), .Y(
        n35241) );
  OA22XL U41599 ( .A0(net263919), .A1(n33076), .B0(n33084), .B1(n40044), .Y(
        n15205) );
  OAI211XL U41600 ( .A0(n33084), .A1(n42940), .B0(n15181), .C0(n15182), .Y(
        n35233) );
  OA22XL U41601 ( .A0(net263919), .A1(n33068), .B0(n33076), .B1(n40043), .Y(
        n15181) );
  OAI211XL U41602 ( .A0(n33076), .A1(n42941), .B0(n15157), .C0(n15158), .Y(
        n35225) );
  OA22XL U41603 ( .A0(net263805), .A1(n33060), .B0(n33068), .B1(n40043), .Y(
        n15157) );
  OAI211XL U41604 ( .A0(n33068), .A1(n42942), .B0(n15133), .C0(n15134), .Y(
        n35217) );
  OA22XL U41605 ( .A0(net218354), .A1(n33052), .B0(n33060), .B1(n40072), .Y(
        n15133) );
  OAI211XL U41606 ( .A0(n33060), .A1(n42943), .B0(n15109), .C0(n15110), .Y(
        n35209) );
  OA22XL U41607 ( .A0(net263957), .A1(n33044), .B0(n33052), .B1(n40042), .Y(
        n15109) );
  OAI211XL U41608 ( .A0(n33052), .A1(n42977), .B0(n15085), .C0(n15086), .Y(
        n35201) );
  OA22XL U41609 ( .A0(net263957), .A1(n33036), .B0(n33044), .B1(n40042), .Y(
        n15085) );
  OAI211XL U41610 ( .A0(n33044), .A1(n42978), .B0(n15061), .C0(n15062), .Y(
        n35193) );
  OA22XL U41611 ( .A0(net263976), .A1(n33028), .B0(n33036), .B1(n40041), .Y(
        n15061) );
  OAI211XL U41612 ( .A0(n33036), .A1(n42979), .B0(n15037), .C0(n15038), .Y(
        n35185) );
  OA22XL U41613 ( .A0(net263976), .A1(n33020), .B0(n33028), .B1(n40041), .Y(
        n15037) );
  OAI211XL U41614 ( .A0(n33028), .A1(n42980), .B0(n15013), .C0(n15014), .Y(
        n35177) );
  OA22XL U41615 ( .A0(net263995), .A1(n33012), .B0(n33020), .B1(n40040), .Y(
        n15013) );
  OAI211XL U41616 ( .A0(n33004), .A1(n42983), .B0(n14941), .C0(n14942), .Y(
        n35153) );
  OA22XL U41617 ( .A0(net263748), .A1(n32988), .B0(n32996), .B1(n40054), .Y(
        n14941) );
  OAI211XL U41618 ( .A0(n32996), .A1(n42985), .B0(n14917), .C0(n14918), .Y(
        n35145) );
  OA22XL U41619 ( .A0(net263748), .A1(n32980), .B0(n32988), .B1(n40053), .Y(
        n14917) );
  OAI211XL U41620 ( .A0(n32988), .A1(n42986), .B0(n14893), .C0(n14894), .Y(
        n35137) );
  OA22XL U41621 ( .A0(net263767), .A1(n32972), .B0(n32980), .B1(n40053), .Y(
        n14893) );
  OAI211XL U41622 ( .A0(n32980), .A1(n42987), .B0(n14869), .C0(n14870), .Y(
        n35129) );
  OA22XL U41623 ( .A0(net263767), .A1(n32964), .B0(n32972), .B1(n40052), .Y(
        n14869) );
  OA22XL U41624 ( .A0(net263292), .A1(n42691), .B0(n32404), .B1(n40079), .Y(
        n13165) );
  OA22XL U41625 ( .A0(net263292), .A1(n42644), .B0(n42691), .B1(n40078), .Y(
        n13141) );
  OAI211XL U41626 ( .A0(n34069), .A1(n42799), .B0(n18136), .C0(n18137), .Y(
        n36218) );
  OA22XL U41627 ( .A0(net262893), .A1(n34053), .B0(n34061), .B1(n40102), .Y(
        n18136) );
  OAI211XL U41628 ( .A0(n34061), .A1(n42800), .B0(n18112), .C0(n18113), .Y(
        n36210) );
  OA22XL U41629 ( .A0(net262893), .A1(n34045), .B0(n34053), .B1(n40131), .Y(
        n18112) );
  OAI211XL U41630 ( .A0(n34053), .A1(n42801), .B0(n18088), .C0(n18089), .Y(
        n36202) );
  OA22XL U41631 ( .A0(net262912), .A1(n34037), .B0(n34045), .B1(n40055), .Y(
        n18088) );
  OAI211XL U41632 ( .A0(n34045), .A1(n42802), .B0(n18064), .C0(n18065), .Y(
        n36194) );
  OA22XL U41633 ( .A0(net262912), .A1(n34029), .B0(n34037), .B1(n40101), .Y(
        n18064) );
  OAI211XL U41634 ( .A0(n34037), .A1(n42803), .B0(n18040), .C0(n18041), .Y(
        n36186) );
  OA22XL U41635 ( .A0(net262912), .A1(n34021), .B0(n34029), .B1(n40101), .Y(
        n18040) );
  OAI211XL U41636 ( .A0(n34029), .A1(n42804), .B0(n18016), .C0(n18017), .Y(
        n36178) );
  OA22XL U41637 ( .A0(net262665), .A1(n34013), .B0(n34021), .B1(n40095), .Y(
        n18016) );
  OAI211XL U41638 ( .A0(n34021), .A1(n42806), .B0(n17992), .C0(n17993), .Y(
        n36170) );
  OA22XL U41639 ( .A0(net262665), .A1(n34005), .B0(n34013), .B1(n40088), .Y(
        n17992) );
  OAI211XL U41640 ( .A0(n34013), .A1(n42807), .B0(n17968), .C0(n17969), .Y(
        n36162) );
  OA22XL U41641 ( .A0(net218364), .A1(n33997), .B0(n34005), .B1(n40111), .Y(
        n17968) );
  OAI211XL U41642 ( .A0(n34005), .A1(n42808), .B0(n17944), .C0(n17945), .Y(
        n36154) );
  OA22XL U41643 ( .A0(net218496), .A1(n33989), .B0(n33997), .B1(n40111), .Y(
        n17944) );
  OAI211XL U41644 ( .A0(n33997), .A1(n42809), .B0(n17920), .C0(n17921), .Y(
        n36146) );
  OA22XL U41645 ( .A0(net218372), .A1(n33981), .B0(n33989), .B1(n40110), .Y(
        n17920) );
  OAI211XL U41646 ( .A0(n33733), .A1(n42766), .B0(n17128), .C0(n17129), .Y(
        n35882) );
  OA22XL U41647 ( .A0(net261886), .A1(n33717), .B0(n33725), .B1(n40150), .Y(
        n17128) );
  OAI211XL U41648 ( .A0(n33725), .A1(n42751), .B0(n17104), .C0(n17105), .Y(
        n35874) );
  OA22XL U41649 ( .A0(net261905), .A1(n33709), .B0(n33717), .B1(n40149), .Y(
        n17104) );
  OAI211XL U41650 ( .A0(n33717), .A1(n42752), .B0(n17080), .C0(n17081), .Y(
        n35866) );
  OA22XL U41651 ( .A0(net261905), .A1(n33701), .B0(n33709), .B1(n40149), .Y(
        n17080) );
  OAI211XL U41652 ( .A0(n33709), .A1(n42753), .B0(n17056), .C0(n17057), .Y(
        n35858) );
  OA22XL U41653 ( .A0(net261924), .A1(n33693), .B0(n33701), .B1(n40148), .Y(
        n17056) );
  OAI211XL U41654 ( .A0(n33701), .A1(n42755), .B0(n17032), .C0(n17033), .Y(
        n35850) );
  OA22XL U41655 ( .A0(net261924), .A1(n33685), .B0(n33693), .B1(n40148), .Y(
        n17032) );
  OAI211XL U41656 ( .A0(n33693), .A1(n42756), .B0(n17008), .C0(n17009), .Y(
        n35842) );
  OA22XL U41657 ( .A0(net261924), .A1(n33677), .B0(n33685), .B1(n40147), .Y(
        n17008) );
  OAI211XL U41658 ( .A0(n33685), .A1(n42757), .B0(n16984), .C0(n16985), .Y(
        n35834) );
  OA22XL U41659 ( .A0(net261943), .A1(n33669), .B0(n33677), .B1(n40147), .Y(
        n16984) );
  OAI211XL U41660 ( .A0(n33677), .A1(n42758), .B0(n16960), .C0(n16961), .Y(
        n35826) );
  OA22XL U41661 ( .A0(net261943), .A1(n33661), .B0(n33669), .B1(n40146), .Y(
        n16960) );
  OAI211XL U41662 ( .A0(n33669), .A1(n42759), .B0(n16936), .C0(n16937), .Y(
        n35818) );
  OA22XL U41663 ( .A0(net218500), .A1(n33653), .B0(n33661), .B1(n40146), .Y(
        n16936) );
  OAI211XL U41664 ( .A0(n33661), .A1(n42760), .B0(n16912), .C0(n16913), .Y(
        n35810) );
  OA22XL U41665 ( .A0(net218482), .A1(n33645), .B0(n33653), .B1(n40145), .Y(
        n16912) );
  OAI211XL U41666 ( .A0(n33653), .A1(n42762), .B0(n16888), .C0(n16889), .Y(
        n35802) );
  OA22XL U41667 ( .A0(net261981), .A1(n33637), .B0(n33645), .B1(n40145), .Y(
        n16888) );
  OAI211XL U41668 ( .A0(n33645), .A1(n42763), .B0(n16864), .C0(n16865), .Y(
        n35794) );
  OA22XL U41669 ( .A0(net262247), .A1(n33629), .B0(n33637), .B1(n40130), .Y(
        n16864) );
  OAI211XL U41670 ( .A0(n33637), .A1(n42764), .B0(n16840), .C0(n16841), .Y(
        n35786) );
  OA22XL U41671 ( .A0(net262266), .A1(n33621), .B0(n33629), .B1(n40130), .Y(
        n16840) );
  OAI211XL U41672 ( .A0(n33629), .A1(n42765), .B0(n16816), .C0(n16817), .Y(
        n35778) );
  OA22XL U41673 ( .A0(net262266), .A1(n33613), .B0(n33621), .B1(n40129), .Y(
        n16816) );
  OAI211XL U41674 ( .A0(n33621), .A1(n42766), .B0(n16792), .C0(n16793), .Y(
        n35770) );
  OA22XL U41675 ( .A0(net262285), .A1(n33605), .B0(n33613), .B1(n40129), .Y(
        n16792) );
  OAI211XL U41676 ( .A0(n33573), .A1(n42741), .B0(n16648), .C0(n16649), .Y(
        n35722) );
  OA22XL U41677 ( .A0(net262323), .A1(n33557), .B0(n33565), .B1(n40127), .Y(
        n16648) );
  OAI211XL U41678 ( .A0(n33565), .A1(n42742), .B0(n16624), .C0(n16625), .Y(
        n35714) );
  OA22XL U41679 ( .A0(net262342), .A1(n33549), .B0(n33557), .B1(n40126), .Y(
        n16624) );
  OAI211XL U41680 ( .A0(n33557), .A1(n42743), .B0(n16600), .C0(n16601), .Y(
        n35706) );
  OA22XL U41681 ( .A0(net262342), .A1(n33541), .B0(n33549), .B1(n40126), .Y(
        n16600) );
  OAI211XL U41682 ( .A0(n33549), .A1(n42744), .B0(n16576), .C0(n16577), .Y(
        n35698) );
  OA22XL U41683 ( .A0(net262361), .A1(n33533), .B0(n33541), .B1(n40125), .Y(
        n16576) );
  OAI211XL U41684 ( .A0(n33541), .A1(n42746), .B0(n16552), .C0(n16553), .Y(
        n35690) );
  OA22XL U41685 ( .A0(net262361), .A1(n33525), .B0(n33533), .B1(n40125), .Y(
        n16552) );
  OAI211XL U41686 ( .A0(n33533), .A1(n42747), .B0(n16528), .C0(n16529), .Y(
        n35682) );
  OA22XL U41687 ( .A0(net262380), .A1(n33517), .B0(n33525), .B1(n40124), .Y(
        n16528) );
  OAI211XL U41688 ( .A0(n33525), .A1(n42748), .B0(n16504), .C0(n16505), .Y(
        n35674) );
  OA22XL U41689 ( .A0(net262380), .A1(n33509), .B0(n33517), .B1(n40124), .Y(
        n16504) );
  OAI211XL U41690 ( .A0(n33517), .A1(n42749), .B0(n16480), .C0(n16481), .Y(
        n35666) );
  OA22XL U41691 ( .A0(net262114), .A1(n33501), .B0(n33509), .B1(n40138), .Y(
        n16480) );
  OAI211XL U41692 ( .A0(n33509), .A1(n42750), .B0(n16456), .C0(n16457), .Y(
        n35658) );
  OA22XL U41693 ( .A0(net262133), .A1(n33493), .B0(n33501), .B1(n40138), .Y(
        n16456) );
  OAI211XL U41694 ( .A0(n33501), .A1(n42783), .B0(n16432), .C0(n16433), .Y(
        n35650) );
  OA22XL U41695 ( .A0(net262133), .A1(n33485), .B0(n33493), .B1(n40137), .Y(
        n16432) );
  OAI211XL U41696 ( .A0(n33493), .A1(n42785), .B0(n16408), .C0(n16409), .Y(
        n35642) );
  OA22XL U41697 ( .A0(net262152), .A1(n33477), .B0(n33485), .B1(n40137), .Y(
        n16408) );
  OAI211XL U41698 ( .A0(n33485), .A1(n42786), .B0(n16384), .C0(n16385), .Y(
        n35634) );
  OA22XL U41699 ( .A0(net262152), .A1(n33469), .B0(n33477), .B1(n40136), .Y(
        n16384) );
  OAI211XL U41700 ( .A0(n33477), .A1(n42787), .B0(n16360), .C0(n16361), .Y(
        n35626) );
  OA22XL U41701 ( .A0(net262152), .A1(n33461), .B0(n33469), .B1(n40136), .Y(
        n16360) );
  OAI211XL U41702 ( .A0(n33469), .A1(n42788), .B0(n16336), .C0(n16337), .Y(
        n35618) );
  OA22XL U41703 ( .A0(net262171), .A1(n33453), .B0(n33461), .B1(n40135), .Y(
        n16336) );
  OAI211XL U41704 ( .A0(n33461), .A1(n42789), .B0(n16312), .C0(n16313), .Y(
        n35610) );
  OA22XL U41705 ( .A0(net262171), .A1(n33445), .B0(n33453), .B1(n40135), .Y(
        n16312) );
  OAI211XL U41706 ( .A0(n33453), .A1(n42790), .B0(n16288), .C0(n16289), .Y(
        n35602) );
  OA22XL U41707 ( .A0(net262190), .A1(n33437), .B0(n33445), .B1(n40134), .Y(
        n16288) );
  OAI211XL U41708 ( .A0(n33445), .A1(n42792), .B0(n16264), .C0(n16265), .Y(
        n35594) );
  OA22XL U41709 ( .A0(net262190), .A1(n33429), .B0(n33437), .B1(n40133), .Y(
        n16264) );
  OAI211XL U41710 ( .A0(n33437), .A1(n42793), .B0(n16240), .C0(n16241), .Y(
        n35586) );
  OA22XL U41711 ( .A0(net262209), .A1(n33421), .B0(n33429), .B1(n40133), .Y(
        n16240) );
  OAI211XL U41712 ( .A0(n33429), .A1(n42794), .B0(n16216), .C0(n16217), .Y(
        n35578) );
  OA22XL U41713 ( .A0(net262209), .A1(n33413), .B0(n33421), .B1(n40132), .Y(
        n16216) );
  OAI211XL U41714 ( .A0(n33421), .A1(n42795), .B0(n16192), .C0(n16193), .Y(
        n35570) );
  OA22XL U41715 ( .A0(net262228), .A1(n33405), .B0(n33413), .B1(n40132), .Y(
        n16192) );
  OAI211XL U41716 ( .A0(n33413), .A1(n42796), .B0(n16168), .C0(n16169), .Y(
        n35562) );
  OA22XL U41717 ( .A0(net262228), .A1(n33397), .B0(n33405), .B1(n40131), .Y(
        n16168) );
  OAI211XL U41718 ( .A0(n33405), .A1(n42797), .B0(n16144), .C0(n16145), .Y(
        n35554) );
  OA22XL U41719 ( .A0(net262247), .A1(n33389), .B0(n33397), .B1(n40131), .Y(
        n16144) );
  OAI211XL U41720 ( .A0(n33397), .A1(n42798), .B0(n16120), .C0(n16121), .Y(
        n35546) );
  OA22XL U41721 ( .A0(net262247), .A1(n33381), .B0(n33389), .B1(n40130), .Y(
        n16120) );
  OAI211XL U41722 ( .A0(n33389), .A1(n42767), .B0(n16096), .C0(n16097), .Y(
        n35538) );
  OA22XL U41723 ( .A0(net263596), .A1(n33373), .B0(n33381), .B1(n40061), .Y(
        n16096) );
  OAI211XL U41724 ( .A0(n33381), .A1(n42768), .B0(n16072), .C0(n16073), .Y(
        n35530) );
  OA22XL U41725 ( .A0(net263615), .A1(n33365), .B0(n33373), .B1(n40061), .Y(
        n16072) );
  OAI211XL U41726 ( .A0(n33373), .A1(n42770), .B0(n16048), .C0(n16049), .Y(
        n35522) );
  OA22XL U41727 ( .A0(net263615), .A1(n33357), .B0(n33365), .B1(n40060), .Y(
        n16048) );
  OAI211XL U41728 ( .A0(n33365), .A1(n42771), .B0(n16024), .C0(n16025), .Y(
        n35514) );
  OA22XL U41729 ( .A0(net263634), .A1(n33349), .B0(n33357), .B1(n40060), .Y(
        n16024) );
  OAI211XL U41730 ( .A0(n33357), .A1(n42772), .B0(n16000), .C0(n16001), .Y(
        n35506) );
  OA22XL U41731 ( .A0(net263634), .A1(n33341), .B0(n33349), .B1(n40059), .Y(
        n16000) );
  OAI211XL U41732 ( .A0(n33349), .A1(n42773), .B0(n15976), .C0(n15977), .Y(
        n35498) );
  OA22XL U41733 ( .A0(net263653), .A1(n33333), .B0(n33341), .B1(n40059), .Y(
        n15976) );
  OAI211XL U41734 ( .A0(n33341), .A1(n42774), .B0(n15952), .C0(n15953), .Y(
        n35490) );
  OA22XL U41735 ( .A0(net263653), .A1(n33325), .B0(n33333), .B1(n40058), .Y(
        n15952) );
  OAI211XL U41736 ( .A0(n33333), .A1(n42775), .B0(n15928), .C0(n15929), .Y(
        n35482) );
  OA22XL U41737 ( .A0(net263653), .A1(n33317), .B0(n33325), .B1(n40058), .Y(
        n15928) );
  OAI211XL U41738 ( .A0(n33325), .A1(n42777), .B0(n15904), .C0(n15905), .Y(
        n35474) );
  OA22XL U41739 ( .A0(net263672), .A1(n33309), .B0(n33317), .B1(n40136), .Y(
        n15904) );
  OAI211XL U41740 ( .A0(n33317), .A1(n42778), .B0(n15880), .C0(n15881), .Y(
        n35466) );
  OA22XL U41741 ( .A0(net263672), .A1(n33301), .B0(n33309), .B1(n40135), .Y(
        n15880) );
  OAI211XL U41742 ( .A0(n33309), .A1(n42779), .B0(n15856), .C0(n15857), .Y(
        n35458) );
  OA22XL U41743 ( .A0(net263691), .A1(n33293), .B0(n33301), .B1(n40057), .Y(
        n15856) );
  OAI211XL U41744 ( .A0(n33301), .A1(n42780), .B0(n15832), .C0(n15833), .Y(
        n35450) );
  OA22XL U41745 ( .A0(net263691), .A1(n33285), .B0(n33293), .B1(n40057), .Y(
        n15832) );
  OAI211XL U41746 ( .A0(n33293), .A1(n42781), .B0(n15808), .C0(n15809), .Y(
        n35442) );
  OA22XL U41747 ( .A0(net263710), .A1(n33277), .B0(n33285), .B1(n40056), .Y(
        n15808) );
  OAI211XL U41748 ( .A0(n33285), .A1(n42782), .B0(n15784), .C0(n15785), .Y(
        n35434) );
  OA22XL U41749 ( .A0(net263710), .A1(n33269), .B0(n33277), .B1(n40056), .Y(
        n15784) );
  OAI211XL U41750 ( .A0(n33277), .A1(n42944), .B0(n15760), .C0(n15761), .Y(
        n35426) );
  OA22XL U41751 ( .A0(net218368), .A1(n33261), .B0(n33269), .B1(n40055), .Y(
        n15760) );
  OAI211XL U41752 ( .A0(n33269), .A1(n42945), .B0(n15736), .C0(n15737), .Y(
        n35418) );
  OA22XL U41753 ( .A0(net218380), .A1(n33253), .B0(n33261), .B1(n40055), .Y(
        n15736) );
  OAI211XL U41754 ( .A0(n33261), .A1(n42946), .B0(n15712), .C0(n15713), .Y(
        n35410) );
  OA22XL U41755 ( .A0(net263463), .A1(n33245), .B0(n33253), .B1(n40069), .Y(
        n15712) );
  OAI211XL U41756 ( .A0(n33253), .A1(n42948), .B0(n15688), .C0(n15689), .Y(
        n35402) );
  OA22XL U41757 ( .A0(net218432), .A1(n33237), .B0(n33245), .B1(n40069), .Y(
        n15688) );
  OAI211XL U41758 ( .A0(n33245), .A1(n42949), .B0(n15664), .C0(n15665), .Y(
        n35394) );
  OA22XL U41759 ( .A0(net263159), .A1(n33229), .B0(n33237), .B1(n40068), .Y(
        n15664) );
  OAI211XL U41760 ( .A0(n33237), .A1(n42950), .B0(n15640), .C0(n15641), .Y(
        n35386) );
  OA22XL U41761 ( .A0(net263501), .A1(n33221), .B0(n33229), .B1(n40068), .Y(
        n15640) );
  OAI211XL U41762 ( .A0(n33229), .A1(n42951), .B0(n15616), .C0(n15617), .Y(
        n35378) );
  OA22XL U41763 ( .A0(net263501), .A1(n33213), .B0(n33221), .B1(n40067), .Y(
        n15616) );
  OAI211XL U41764 ( .A0(n33221), .A1(n42952), .B0(n15592), .C0(n15593), .Y(
        n35370) );
  OA22XL U41765 ( .A0(net218532), .A1(n33205), .B0(n33213), .B1(n40067), .Y(
        n15592) );
  OAI211XL U41766 ( .A0(n33213), .A1(n42953), .B0(n15568), .C0(n15569), .Y(
        n35362) );
  OA22XL U41767 ( .A0(net218302), .A1(n33197), .B0(n33205), .B1(n40066), .Y(
        n15568) );
  OAI211XL U41768 ( .A0(n33205), .A1(n42955), .B0(n15544), .C0(n15545), .Y(
        n35354) );
  OA22XL U41769 ( .A0(net218486), .A1(n33189), .B0(n33197), .B1(n40066), .Y(
        n15544) );
  OAI211XL U41770 ( .A0(n33197), .A1(n42956), .B0(n15520), .C0(n15521), .Y(
        n35346) );
  OA22XL U41771 ( .A0(net263539), .A1(n33181), .B0(n33189), .B1(n40065), .Y(
        n15520) );
  OAI211XL U41772 ( .A0(n33189), .A1(n42957), .B0(n15496), .C0(n15497), .Y(
        n35338) );
  OA22XL U41773 ( .A0(net263539), .A1(n33173), .B0(n33181), .B1(n40065), .Y(
        n15496) );
  OAI211XL U41774 ( .A0(n33181), .A1(n42958), .B0(n15472), .C0(n15473), .Y(
        n35330) );
  OA22XL U41775 ( .A0(net263558), .A1(n33165), .B0(n33173), .B1(n40064), .Y(
        n15472) );
  OAI211XL U41776 ( .A0(n33173), .A1(n42959), .B0(n15448), .C0(n15449), .Y(
        n35322) );
  OA22XL U41777 ( .A0(net263558), .A1(n33157), .B0(n33165), .B1(n40064), .Y(
        n15448) );
  OAI211XL U41778 ( .A0(n33165), .A1(n42928), .B0(n15424), .C0(n15425), .Y(
        n35314) );
  OA22XL U41779 ( .A0(net263577), .A1(n33149), .B0(n33157), .B1(n40063), .Y(
        n15424) );
  OAI211XL U41780 ( .A0(n33157), .A1(n42929), .B0(n15400), .C0(n15401), .Y(
        n35306) );
  OA22XL U41781 ( .A0(net263577), .A1(n33141), .B0(n33149), .B1(n40063), .Y(
        n15400) );
  OAI211XL U41782 ( .A0(n33149), .A1(n42930), .B0(n15376), .C0(n15377), .Y(
        n35298) );
  OA22XL U41783 ( .A0(net263596), .A1(n33133), .B0(n33141), .B1(n40062), .Y(
        n15376) );
  OAI211XL U41784 ( .A0(n33141), .A1(n42931), .B0(n15352), .C0(n15353), .Y(
        n35290) );
  OA22XL U41785 ( .A0(net263596), .A1(n33125), .B0(n33133), .B1(n40062), .Y(
        n15352) );
  OAI211XL U41786 ( .A0(n33133), .A1(n42933), .B0(n15328), .C0(n15329), .Y(
        n35282) );
  OA22XL U41787 ( .A0(net263881), .A1(n33117), .B0(n33125), .B1(n40046), .Y(
        n15328) );
  OAI211XL U41788 ( .A0(n33125), .A1(n42934), .B0(n15304), .C0(n15305), .Y(
        n35274) );
  OA22XL U41789 ( .A0(net263881), .A1(n33109), .B0(n33117), .B1(n40046), .Y(
        n15304) );
  OAI211XL U41790 ( .A0(n33117), .A1(n42935), .B0(n15280), .C0(n15281), .Y(
        n35266) );
  OA22XL U41791 ( .A0(net263900), .A1(n33101), .B0(n33109), .B1(n40045), .Y(
        n15280) );
  OAI211XL U41792 ( .A0(n33109), .A1(n42936), .B0(n15256), .C0(n15257), .Y(
        n35258) );
  OA22XL U41793 ( .A0(net263900), .A1(n33093), .B0(n33101), .B1(n40045), .Y(
        n15256) );
  OAI211XL U41794 ( .A0(n33101), .A1(n42937), .B0(n15232), .C0(n15233), .Y(
        n35250) );
  OA22XL U41795 ( .A0(net263900), .A1(n33085), .B0(n33093), .B1(n40044), .Y(
        n15232) );
  OAI211XL U41796 ( .A0(n33093), .A1(n42938), .B0(n15208), .C0(n15209), .Y(
        n35242) );
  OA22XL U41797 ( .A0(net263919), .A1(n33077), .B0(n33085), .B1(n40044), .Y(
        n15208) );
  OAI211XL U41798 ( .A0(n33085), .A1(n42940), .B0(n15184), .C0(n15185), .Y(
        n35234) );
  OA22XL U41799 ( .A0(net263919), .A1(n33069), .B0(n33077), .B1(n40043), .Y(
        n15184) );
  OAI211XL U41800 ( .A0(n33077), .A1(n42941), .B0(n15160), .C0(n15161), .Y(
        n35226) );
  OA22XL U41801 ( .A0(net218504), .A1(n33061), .B0(n33069), .B1(n40043), .Y(
        n15160) );
  OAI211XL U41802 ( .A0(n33069), .A1(n42942), .B0(n15136), .C0(n15137), .Y(
        n35218) );
  OA22XL U41803 ( .A0(net218352), .A1(n33053), .B0(n33061), .B1(n40062), .Y(
        n15136) );
  OAI211XL U41804 ( .A0(n33061), .A1(n42943), .B0(n15112), .C0(n15113), .Y(
        n35210) );
  OA22XL U41805 ( .A0(net263957), .A1(n33045), .B0(n33053), .B1(n40133), .Y(
        n15112) );
  OAI211XL U41806 ( .A0(n33053), .A1(n42976), .B0(n15088), .C0(n15089), .Y(
        n35202) );
  OA22XL U41807 ( .A0(net263957), .A1(n33037), .B0(n33045), .B1(n40042), .Y(
        n15088) );
  OAI211XL U41808 ( .A0(n33045), .A1(n42978), .B0(n15064), .C0(n15065), .Y(
        n35194) );
  OA22XL U41809 ( .A0(net263976), .A1(n33029), .B0(n33037), .B1(n40042), .Y(
        n15064) );
  OAI211XL U41810 ( .A0(n33037), .A1(n42979), .B0(n15040), .C0(n15041), .Y(
        n35186) );
  OA22XL U41811 ( .A0(net263976), .A1(n33021), .B0(n33029), .B1(n40041), .Y(
        n15040) );
  OAI211XL U41812 ( .A0(n33029), .A1(n42984), .B0(n15016), .C0(n15017), .Y(
        n35178) );
  OA22XL U41813 ( .A0(net263976), .A1(n33013), .B0(n33021), .B1(n40041), .Y(
        n15016) );
  OAI211XL U41814 ( .A0(n33021), .A1(n42981), .B0(n14992), .C0(n14993), .Y(
        n35170) );
  OA22XL U41815 ( .A0(net263995), .A1(n33005), .B0(n33013), .B1(n40040), .Y(
        n14992) );
  OAI211XL U41816 ( .A0(n33013), .A1(n42982), .B0(n14968), .C0(n14969), .Y(
        n35162) );
  OA22XL U41817 ( .A0(net263995), .A1(n32997), .B0(n33005), .B1(n40040), .Y(
        n14968) );
  OAI211XL U41818 ( .A0(n33005), .A1(n42983), .B0(n14944), .C0(n14945), .Y(
        n35154) );
  OA22XL U41819 ( .A0(net263748), .A1(n32989), .B0(n32997), .B1(n40054), .Y(
        n14944) );
  OAI211XL U41820 ( .A0(n32997), .A1(n42984), .B0(n14920), .C0(n14921), .Y(
        n35146) );
  OA22XL U41821 ( .A0(net263748), .A1(n32981), .B0(n32989), .B1(n40054), .Y(
        n14920) );
  OA22XL U41822 ( .A0(net263767), .A1(n32965), .B0(n32973), .B1(n40053), .Y(
        n14872) );
  OA22XL U41823 ( .A0(net263292), .A1(n41283), .B0(n32405), .B1(n40079), .Y(
        n13168) );
  OA22XL U41824 ( .A0(net263292), .A1(n42626), .B0(n41281), .B1(n40078), .Y(
        n13144) );
  OAI211XL U41825 ( .A0(n34070), .A1(n42807), .B0(n18139), .C0(n18140), .Y(
        n36219) );
  OA22XL U41826 ( .A0(net262893), .A1(n34054), .B0(n34062), .B1(n40102), .Y(
        n18139) );
  OAI211XL U41827 ( .A0(n34062), .A1(n42800), .B0(n18115), .C0(n18116), .Y(
        n36211) );
  OA22XL U41828 ( .A0(net262893), .A1(n34046), .B0(n34054), .B1(n40132), .Y(
        n18115) );
  OAI211XL U41829 ( .A0(n34054), .A1(n42801), .B0(n18091), .C0(n18092), .Y(
        n36203) );
  OA22XL U41830 ( .A0(net262893), .A1(n34038), .B0(n34046), .B1(n40123), .Y(
        n18091) );
  OAI211XL U41831 ( .A0(n34046), .A1(n42802), .B0(n18067), .C0(n18068), .Y(
        n36195) );
  OA22XL U41832 ( .A0(net262912), .A1(n34030), .B0(n34038), .B1(n40101), .Y(
        n18067) );
  OAI211XL U41833 ( .A0(n34038), .A1(n42803), .B0(n18043), .C0(n18044), .Y(
        n36187) );
  OA22XL U41834 ( .A0(net262912), .A1(n34022), .B0(n34030), .B1(n40101), .Y(
        n18043) );
  OAI211XL U41835 ( .A0(n34030), .A1(n42804), .B0(n18019), .C0(n18020), .Y(
        n36179) );
  OA22XL U41836 ( .A0(net262665), .A1(n34014), .B0(n34022), .B1(n40089), .Y(
        n18019) );
  OAI211XL U41837 ( .A0(n34022), .A1(n42805), .B0(n17995), .C0(n17996), .Y(
        n36171) );
  OA22XL U41838 ( .A0(net262665), .A1(n34006), .B0(n34014), .B1(n40087), .Y(
        n17995) );
  OAI211XL U41839 ( .A0(n34014), .A1(n42807), .B0(n17971), .C0(n17972), .Y(
        n36163) );
  OA22XL U41840 ( .A0(net262665), .A1(n33998), .B0(n34006), .B1(n40111), .Y(
        n17971) );
  OAI211XL U41841 ( .A0(n34006), .A1(n42808), .B0(n17947), .C0(n17948), .Y(
        n36155) );
  OA22XL U41842 ( .A0(net218342), .A1(n33990), .B0(n33998), .B1(n40111), .Y(
        n17947) );
  OAI211XL U41843 ( .A0(n33998), .A1(n42809), .B0(n17923), .C0(n17924), .Y(
        n36147) );
  OA22XL U41844 ( .A0(net218402), .A1(n33982), .B0(n33990), .B1(n40110), .Y(
        n17923) );
  OAI211XL U41845 ( .A0(n33726), .A1(n42751), .B0(n17107), .C0(n17108), .Y(
        n35875) );
  OA22XL U41846 ( .A0(net261905), .A1(n33710), .B0(n33718), .B1(n40149), .Y(
        n17107) );
  OAI211XL U41847 ( .A0(n33718), .A1(n42752), .B0(n17083), .C0(n17084), .Y(
        n35867) );
  OA22XL U41848 ( .A0(net261905), .A1(n33702), .B0(n33710), .B1(n40149), .Y(
        n17083) );
  OAI211XL U41849 ( .A0(n33710), .A1(n42753), .B0(n17059), .C0(n17060), .Y(
        n35859) );
  OA22XL U41850 ( .A0(net261924), .A1(n33694), .B0(n33702), .B1(n40148), .Y(
        n17059) );
  OAI211XL U41851 ( .A0(n33702), .A1(n42754), .B0(n17035), .C0(n17036), .Y(
        n35851) );
  OA22XL U41852 ( .A0(net261924), .A1(n33686), .B0(n33694), .B1(n40148), .Y(
        n17035) );
  OAI211XL U41853 ( .A0(n33694), .A1(n42756), .B0(n17011), .C0(n17012), .Y(
        n35843) );
  OA22XL U41854 ( .A0(net261924), .A1(n33678), .B0(n33686), .B1(n40147), .Y(
        n17011) );
  OAI211XL U41855 ( .A0(n33686), .A1(n42757), .B0(n16987), .C0(n16988), .Y(
        n35835) );
  OA22XL U41856 ( .A0(net261943), .A1(n33670), .B0(n33678), .B1(n40147), .Y(
        n16987) );
  OAI211XL U41857 ( .A0(n33678), .A1(n42758), .B0(n16963), .C0(n16964), .Y(
        n35827) );
  OA22XL U41858 ( .A0(net261943), .A1(n33662), .B0(n33670), .B1(n40146), .Y(
        n16963) );
  OAI211XL U41859 ( .A0(n33670), .A1(n42759), .B0(n16939), .C0(n16940), .Y(
        n35819) );
  OA22XL U41860 ( .A0(net218502), .A1(n33654), .B0(n33662), .B1(n40146), .Y(
        n16939) );
  OAI211XL U41861 ( .A0(n33662), .A1(n42760), .B0(n16915), .C0(n16916), .Y(
        n35811) );
  OA22XL U41862 ( .A0(net218454), .A1(n33646), .B0(n33654), .B1(n40145), .Y(
        n16915) );
  OAI211XL U41863 ( .A0(n33654), .A1(n42761), .B0(n16891), .C0(n16892), .Y(
        n35803) );
  OA22XL U41864 ( .A0(net261981), .A1(n33638), .B0(n33646), .B1(n40145), .Y(
        n16891) );
  OAI211XL U41865 ( .A0(n33646), .A1(n42763), .B0(n16867), .C0(n16868), .Y(
        n35795) );
  OA22XL U41866 ( .A0(net262247), .A1(n33630), .B0(n33638), .B1(n40130), .Y(
        n16867) );
  OAI211XL U41867 ( .A0(n33638), .A1(n42764), .B0(n16843), .C0(n16844), .Y(
        n35787) );
  OA22XL U41868 ( .A0(net262266), .A1(n33622), .B0(n33630), .B1(n40130), .Y(
        n16843) );
  OAI211XL U41869 ( .A0(n33630), .A1(n42765), .B0(n16819), .C0(n16820), .Y(
        n35779) );
  OA22XL U41870 ( .A0(net262266), .A1(n33614), .B0(n33622), .B1(n40129), .Y(
        n16819) );
  OAI211XL U41871 ( .A0(n33622), .A1(n42766), .B0(n16795), .C0(n16796), .Y(
        n35771) );
  OA22XL U41872 ( .A0(net262285), .A1(n33606), .B0(n33614), .B1(n40129), .Y(
        n16795) );
  OAI211XL U41873 ( .A0(n33574), .A1(n42741), .B0(n16651), .C0(n16652), .Y(
        n35723) );
  OA22XL U41874 ( .A0(net262323), .A1(n33558), .B0(n33566), .B1(n40127), .Y(
        n16651) );
  OAI211XL U41875 ( .A0(n33566), .A1(n42742), .B0(n16627), .C0(n16628), .Y(
        n35715) );
  OA22XL U41876 ( .A0(net262342), .A1(n33550), .B0(n33558), .B1(n40126), .Y(
        n16627) );
  OAI211XL U41877 ( .A0(n33558), .A1(n42743), .B0(n16603), .C0(n16604), .Y(
        n35707) );
  OA22XL U41878 ( .A0(net262342), .A1(n33542), .B0(n33550), .B1(n40126), .Y(
        n16603) );
  OAI211XL U41879 ( .A0(n33550), .A1(n42744), .B0(n16579), .C0(n16580), .Y(
        n35699) );
  OA22XL U41880 ( .A0(net262361), .A1(n33534), .B0(n33542), .B1(n40125), .Y(
        n16579) );
  OAI211XL U41881 ( .A0(n33542), .A1(n42745), .B0(n16555), .C0(n16556), .Y(
        n35691) );
  OA22XL U41882 ( .A0(net262361), .A1(n33526), .B0(n33534), .B1(n40125), .Y(
        n16555) );
  OAI211XL U41883 ( .A0(n33534), .A1(n42747), .B0(n16531), .C0(n16532), .Y(
        n35683) );
  OA22XL U41884 ( .A0(net262380), .A1(n33518), .B0(n33526), .B1(n40124), .Y(
        n16531) );
  OAI211XL U41885 ( .A0(n33526), .A1(n42748), .B0(n16507), .C0(n16508), .Y(
        n35675) );
  OA22XL U41886 ( .A0(net262380), .A1(n33510), .B0(n33518), .B1(n40124), .Y(
        n16507) );
  OAI211XL U41887 ( .A0(n33518), .A1(n42749), .B0(n16483), .C0(n16484), .Y(
        n35667) );
  OA22XL U41888 ( .A0(net262114), .A1(n33502), .B0(n33510), .B1(n40138), .Y(
        n16483) );
  OAI211XL U41889 ( .A0(n33510), .A1(n42750), .B0(n16459), .C0(n16460), .Y(
        n35659) );
  OA22XL U41890 ( .A0(net262133), .A1(n33494), .B0(n33502), .B1(n40138), .Y(
        n16459) );
  OAI211XL U41891 ( .A0(n33502), .A1(n42783), .B0(n16435), .C0(n16436), .Y(
        n35651) );
  OA22XL U41892 ( .A0(net262133), .A1(n33486), .B0(n33494), .B1(n40137), .Y(
        n16435) );
  OAI211XL U41893 ( .A0(n33494), .A1(n42784), .B0(n16411), .C0(n16412), .Y(
        n35643) );
  OA22XL U41894 ( .A0(net262152), .A1(n33478), .B0(n33486), .B1(n40137), .Y(
        n16411) );
  OAI211XL U41895 ( .A0(n33486), .A1(n42786), .B0(n16387), .C0(n16388), .Y(
        n35635) );
  OA22XL U41896 ( .A0(net262152), .A1(n33470), .B0(n33478), .B1(n40136), .Y(
        n16387) );
  OAI211XL U41897 ( .A0(n33478), .A1(n42787), .B0(n16363), .C0(n16364), .Y(
        n35627) );
  OA22XL U41898 ( .A0(net262152), .A1(n33462), .B0(n33470), .B1(n40136), .Y(
        n16363) );
  OAI211XL U41899 ( .A0(n33470), .A1(n42788), .B0(n16339), .C0(n16340), .Y(
        n35619) );
  OA22XL U41900 ( .A0(net262171), .A1(n33454), .B0(n33462), .B1(n40135), .Y(
        n16339) );
  OAI211XL U41901 ( .A0(n33462), .A1(n42789), .B0(n16315), .C0(n16316), .Y(
        n35611) );
  OA22XL U41902 ( .A0(net262171), .A1(n33446), .B0(n33454), .B1(n40135), .Y(
        n16315) );
  OAI211XL U41903 ( .A0(n33454), .A1(n42790), .B0(n16291), .C0(n16292), .Y(
        n35603) );
  OA22XL U41904 ( .A0(net262190), .A1(n33438), .B0(n33446), .B1(n40134), .Y(
        n16291) );
  OAI211XL U41905 ( .A0(n33446), .A1(n42791), .B0(n16267), .C0(n16268), .Y(
        n35595) );
  OA22XL U41906 ( .A0(net262190), .A1(n33430), .B0(n33438), .B1(n40134), .Y(
        n16267) );
  OAI211XL U41907 ( .A0(n33438), .A1(n42793), .B0(n16243), .C0(n16244), .Y(
        n35587) );
  OA22XL U41908 ( .A0(net262209), .A1(n33422), .B0(n33430), .B1(n40133), .Y(
        n16243) );
  OAI211XL U41909 ( .A0(n33430), .A1(n42794), .B0(n16219), .C0(n16220), .Y(
        n35579) );
  OA22XL U41910 ( .A0(net262209), .A1(n33414), .B0(n33422), .B1(n40133), .Y(
        n16219) );
  OAI211XL U41911 ( .A0(n33422), .A1(n42795), .B0(n16195), .C0(n16196), .Y(
        n35571) );
  OA22XL U41912 ( .A0(net262228), .A1(n33406), .B0(n33414), .B1(n40132), .Y(
        n16195) );
  OAI211XL U41913 ( .A0(n33414), .A1(n42796), .B0(n16171), .C0(n16172), .Y(
        n35563) );
  OA22XL U41914 ( .A0(net262228), .A1(n33398), .B0(n33406), .B1(n40132), .Y(
        n16171) );
  OAI211XL U41915 ( .A0(n33406), .A1(n42797), .B0(n16147), .C0(n16148), .Y(
        n35555) );
  OA22XL U41916 ( .A0(net262228), .A1(n33390), .B0(n33398), .B1(n40131), .Y(
        n16147) );
  OAI211XL U41917 ( .A0(n33398), .A1(n42798), .B0(n16123), .C0(n16124), .Y(
        n35547) );
  OA22XL U41918 ( .A0(net262247), .A1(n33382), .B0(n33390), .B1(n40131), .Y(
        n16123) );
  OAI211XL U41919 ( .A0(n33390), .A1(n42767), .B0(n16099), .C0(n16100), .Y(
        n35539) );
  OA22XL U41920 ( .A0(net263596), .A1(n33374), .B0(n33382), .B1(n40061), .Y(
        n16099) );
  OAI211XL U41921 ( .A0(n33382), .A1(n42768), .B0(n16075), .C0(n16076), .Y(
        n35531) );
  OA22XL U41922 ( .A0(net263615), .A1(n33366), .B0(n33374), .B1(n40061), .Y(
        n16075) );
  OAI211XL U41923 ( .A0(n33374), .A1(n42769), .B0(n16051), .C0(n16052), .Y(
        n35523) );
  OA22XL U41924 ( .A0(net263615), .A1(n33358), .B0(n33366), .B1(n40060), .Y(
        n16051) );
  OAI211XL U41925 ( .A0(n33366), .A1(n42771), .B0(n16027), .C0(n16028), .Y(
        n35515) );
  OA22XL U41926 ( .A0(net263634), .A1(n33350), .B0(n33358), .B1(n40060), .Y(
        n16027) );
  OAI211XL U41927 ( .A0(n33358), .A1(n42772), .B0(n16003), .C0(n16004), .Y(
        n35507) );
  OA22XL U41928 ( .A0(net263634), .A1(n33342), .B0(n33350), .B1(n40059), .Y(
        n16003) );
  OAI211XL U41929 ( .A0(n33350), .A1(n42773), .B0(n15979), .C0(n15980), .Y(
        n35499) );
  OA22XL U41930 ( .A0(net263653), .A1(n33334), .B0(n33342), .B1(n40059), .Y(
        n15979) );
  OAI211XL U41931 ( .A0(n33342), .A1(n42774), .B0(n15955), .C0(n15956), .Y(
        n35491) );
  OA22XL U41932 ( .A0(net263653), .A1(n33326), .B0(n33334), .B1(n40058), .Y(
        n15955) );
  OAI211XL U41933 ( .A0(n33334), .A1(n42775), .B0(n15931), .C0(n15932), .Y(
        n35483) );
  OA22XL U41934 ( .A0(net263653), .A1(n33318), .B0(n33326), .B1(n40058), .Y(
        n15931) );
  OAI211XL U41935 ( .A0(n33326), .A1(n42776), .B0(n15907), .C0(n15908), .Y(
        n35475) );
  OA22XL U41936 ( .A0(net263672), .A1(n33310), .B0(n33318), .B1(n40135), .Y(
        n15907) );
  OAI211XL U41937 ( .A0(n33318), .A1(n42778), .B0(n15883), .C0(n15884), .Y(
        n35467) );
  OA22XL U41938 ( .A0(net263672), .A1(n33302), .B0(n33310), .B1(n40136), .Y(
        n15883) );
  OAI211XL U41939 ( .A0(n33310), .A1(n42779), .B0(n15859), .C0(n15860), .Y(
        n35459) );
  OA22XL U41940 ( .A0(net263691), .A1(n33294), .B0(n33302), .B1(n40057), .Y(
        n15859) );
  OAI211XL U41941 ( .A0(n33302), .A1(n42780), .B0(n15835), .C0(n15836), .Y(
        n35451) );
  OA22XL U41942 ( .A0(net263691), .A1(n33286), .B0(n33294), .B1(n40057), .Y(
        n15835) );
  OAI211XL U41943 ( .A0(n33294), .A1(n42781), .B0(n15811), .C0(n15812), .Y(
        n35443) );
  OA22XL U41944 ( .A0(net263710), .A1(n33278), .B0(n33286), .B1(n40056), .Y(
        n15811) );
  OAI211XL U41945 ( .A0(n33286), .A1(n42782), .B0(n15787), .C0(n15788), .Y(
        n35435) );
  OA22XL U41946 ( .A0(net263710), .A1(n33270), .B0(n33278), .B1(n40056), .Y(
        n15787) );
  OAI211XL U41947 ( .A0(n33278), .A1(n42944), .B0(n15763), .C0(n15764), .Y(
        n35427) );
  OA22XL U41948 ( .A0(net218472), .A1(n33262), .B0(n33270), .B1(n40055), .Y(
        n15763) );
  OAI211XL U41949 ( .A0(n33270), .A1(n42945), .B0(n15739), .C0(n15740), .Y(
        n35419) );
  OA22XL U41950 ( .A0(net218412), .A1(n33254), .B0(n33262), .B1(n40055), .Y(
        n15739) );
  OAI211XL U41951 ( .A0(n33262), .A1(n42946), .B0(n15715), .C0(n15716), .Y(
        n35411) );
  OA22XL U41952 ( .A0(net263463), .A1(n33246), .B0(n33254), .B1(n40069), .Y(
        n15715) );
  OAI211XL U41953 ( .A0(n33254), .A1(n42947), .B0(n15691), .C0(n15692), .Y(
        n35403) );
  OA22XL U41954 ( .A0(net218374), .A1(n33238), .B0(n33246), .B1(n40069), .Y(
        n15691) );
  OAI211XL U41955 ( .A0(n33246), .A1(n42949), .B0(n15667), .C0(n15668), .Y(
        n35395) );
  OA22XL U41956 ( .A0(net218396), .A1(n33230), .B0(n33238), .B1(n40068), .Y(
        n15667) );
  OAI211XL U41957 ( .A0(n33238), .A1(n42950), .B0(n15643), .C0(n15644), .Y(
        n35387) );
  OA22XL U41958 ( .A0(net263501), .A1(n33222), .B0(n33230), .B1(n40068), .Y(
        n15643) );
  OAI211XL U41959 ( .A0(n33230), .A1(n42951), .B0(n15619), .C0(n15620), .Y(
        n35379) );
  OA22XL U41960 ( .A0(net263501), .A1(n33214), .B0(n33222), .B1(n40067), .Y(
        n15619) );
  OAI211XL U41961 ( .A0(n33222), .A1(n42952), .B0(n15595), .C0(n15596), .Y(
        n35371) );
  OA22XL U41962 ( .A0(net263501), .A1(n33206), .B0(n33214), .B1(n40067), .Y(
        n15595) );
  OAI211XL U41963 ( .A0(n33214), .A1(n42953), .B0(n15571), .C0(n15572), .Y(
        n35363) );
  OA22XL U41964 ( .A0(net218386), .A1(n33198), .B0(n33206), .B1(n40066), .Y(
        n15571) );
  OAI211XL U41965 ( .A0(n33206), .A1(n42954), .B0(n15547), .C0(n15548), .Y(
        n35355) );
  OA22XL U41966 ( .A0(net218494), .A1(n33190), .B0(n33198), .B1(n40066), .Y(
        n15547) );
  OAI211XL U41967 ( .A0(n33198), .A1(n42956), .B0(n15523), .C0(n15524), .Y(
        n35347) );
  OA22XL U41968 ( .A0(net263539), .A1(n33182), .B0(n33190), .B1(n40065), .Y(
        n15523) );
  OAI211XL U41969 ( .A0(n33190), .A1(n42957), .B0(n15499), .C0(n15500), .Y(
        n35339) );
  OA22XL U41970 ( .A0(net263539), .A1(n33174), .B0(n33182), .B1(n40065), .Y(
        n15499) );
  OAI211XL U41971 ( .A0(n33182), .A1(n42958), .B0(n15475), .C0(n15476), .Y(
        n35331) );
  OA22XL U41972 ( .A0(net263558), .A1(n33166), .B0(n33174), .B1(n40064), .Y(
        n15475) );
  OAI211XL U41973 ( .A0(n33174), .A1(n42959), .B0(n15451), .C0(n15452), .Y(
        n35323) );
  OA22XL U41974 ( .A0(net263558), .A1(n33158), .B0(n33166), .B1(n40064), .Y(
        n15451) );
  OAI211XL U41975 ( .A0(n33166), .A1(n42928), .B0(n15427), .C0(n15428), .Y(
        n35315) );
  OA22XL U41976 ( .A0(net263577), .A1(n33150), .B0(n33158), .B1(n40063), .Y(
        n15427) );
  OAI211XL U41977 ( .A0(n33158), .A1(n42929), .B0(n15403), .C0(n15404), .Y(
        n35307) );
  OA22XL U41978 ( .A0(net263577), .A1(n33142), .B0(n33150), .B1(n40063), .Y(
        n15403) );
  OAI211XL U41979 ( .A0(n33150), .A1(n42930), .B0(n15379), .C0(n15380), .Y(
        n35299) );
  OA22XL U41980 ( .A0(net263596), .A1(n33134), .B0(n33142), .B1(n40062), .Y(
        n15379) );
  OAI211XL U41981 ( .A0(n33142), .A1(n42931), .B0(n15355), .C0(n15356), .Y(
        n35291) );
  OA22XL U41982 ( .A0(net263596), .A1(n33126), .B0(n33134), .B1(n40062), .Y(
        n15355) );
  OAI211XL U41983 ( .A0(n33134), .A1(n42932), .B0(n15331), .C0(n15332), .Y(
        n35283) );
  OA22XL U41984 ( .A0(net263881), .A1(n33118), .B0(n33126), .B1(n40046), .Y(
        n15331) );
  OAI211XL U41985 ( .A0(n33126), .A1(n42934), .B0(n15307), .C0(n15308), .Y(
        n35275) );
  OA22XL U41986 ( .A0(net263881), .A1(n33110), .B0(n33118), .B1(n40046), .Y(
        n15307) );
  OAI211XL U41987 ( .A0(n33118), .A1(n42935), .B0(n15283), .C0(n15284), .Y(
        n35267) );
  OA22XL U41988 ( .A0(net263881), .A1(n33102), .B0(n33110), .B1(n40045), .Y(
        n15283) );
  OAI211XL U41989 ( .A0(n33110), .A1(n42936), .B0(n15259), .C0(n15260), .Y(
        n35259) );
  OA22XL U41990 ( .A0(net263900), .A1(n33094), .B0(n33102), .B1(n40045), .Y(
        n15259) );
  OAI211XL U41991 ( .A0(n33102), .A1(n42937), .B0(n15235), .C0(n15236), .Y(
        n35251) );
  OA22XL U41992 ( .A0(net263900), .A1(n33086), .B0(n33094), .B1(n40044), .Y(
        n15235) );
  OAI211XL U41993 ( .A0(n33094), .A1(n42938), .B0(n15211), .C0(n15212), .Y(
        n35243) );
  OA22XL U41994 ( .A0(net263919), .A1(n33078), .B0(n33086), .B1(n40044), .Y(
        n15211) );
  OAI211XL U41995 ( .A0(n33086), .A1(n42939), .B0(n15187), .C0(n15188), .Y(
        n35235) );
  OA22XL U41996 ( .A0(net263919), .A1(n33070), .B0(n33078), .B1(n40043), .Y(
        n15187) );
  OAI211XL U41997 ( .A0(n33078), .A1(n42941), .B0(n15163), .C0(n15164), .Y(
        n35227) );
  OA22XL U41998 ( .A0(net262931), .A1(n33062), .B0(n33070), .B1(n40043), .Y(
        n15163) );
  OAI211XL U41999 ( .A0(n33070), .A1(n42942), .B0(n15139), .C0(n15140), .Y(
        n35219) );
  OA22XL U42000 ( .A0(net218442), .A1(n33054), .B0(n33062), .B1(n40072), .Y(
        n15139) );
  OAI211XL U42001 ( .A0(n33062), .A1(n42943), .B0(n15115), .C0(n15116), .Y(
        n35211) );
  OA22XL U42002 ( .A0(net263957), .A1(n33046), .B0(n33054), .B1(n40062), .Y(
        n15115) );
  OAI211XL U42003 ( .A0(n33054), .A1(n42976), .B0(n15091), .C0(n15092), .Y(
        n35203) );
  OA22XL U42004 ( .A0(net263957), .A1(n33038), .B0(n33046), .B1(n40042), .Y(
        n15091) );
  OAI211XL U42005 ( .A0(n33046), .A1(n42977), .B0(n15067), .C0(n15068), .Y(
        n35195) );
  OA22XL U42006 ( .A0(net263976), .A1(n33030), .B0(n33038), .B1(n40042), .Y(
        n15067) );
  OAI211XL U42007 ( .A0(n33038), .A1(n42979), .B0(n15043), .C0(n15044), .Y(
        n35187) );
  OA22XL U42008 ( .A0(net263976), .A1(n33022), .B0(n33030), .B1(n40041), .Y(
        n15043) );
  OAI211XL U42009 ( .A0(n33030), .A1(n42980), .B0(n15019), .C0(n15020), .Y(
        n35179) );
  OA22XL U42010 ( .A0(net263976), .A1(n33014), .B0(n33022), .B1(n40041), .Y(
        n15019) );
  OAI211XL U42011 ( .A0(n33022), .A1(n42981), .B0(n14995), .C0(n14996), .Y(
        n35171) );
  OA22XL U42012 ( .A0(net263995), .A1(n33006), .B0(n33014), .B1(n40040), .Y(
        n14995) );
  OAI211XL U42013 ( .A0(n33014), .A1(n42982), .B0(n14971), .C0(n14972), .Y(
        n35163) );
  OA22XL U42014 ( .A0(net263995), .A1(n32998), .B0(n33006), .B1(n40040), .Y(
        n14971) );
  OAI211XL U42015 ( .A0(n33006), .A1(n42983), .B0(n14947), .C0(n14948), .Y(
        n35155) );
  OA22XL U42016 ( .A0(net263748), .A1(n32990), .B0(n32998), .B1(n40054), .Y(
        n14947) );
  OAI211XL U42017 ( .A0(n32998), .A1(n42984), .B0(n14923), .C0(n14924), .Y(
        n35147) );
  OA22XL U42018 ( .A0(net263748), .A1(n32982), .B0(n32990), .B1(n40054), .Y(
        n14923) );
  OA22XL U42019 ( .A0(net263748), .A1(n32974), .B0(n32982), .B1(n40053), .Y(
        n14899) );
  OA22XL U42020 ( .A0(net263767), .A1(n32966), .B0(n32974), .B1(n40053), .Y(
        n14875) );
  OA22XL U42021 ( .A0(net263292), .A1(net219310), .B0(n32406), .B1(n40079),
        .Y(n13171) );
  OA22XL U42022 ( .A0(net263292), .A1(n42620), .B0(net219310), .B1(n40078),
        .Y(n13147) );
  OAI211XL U42023 ( .A0(n34064), .A1(n42799), .B0(n18121), .C0(n18122), .Y(
        n36213) );
  OA22XL U42024 ( .A0(net262893), .A1(n34048), .B0(n34056), .B1(n40124), .Y(
        n18121) );
  OAI211XL U42025 ( .A0(n34056), .A1(n42801), .B0(n18097), .C0(n18098), .Y(
        n36205) );
  OA22XL U42026 ( .A0(net262893), .A1(n34040), .B0(n34048), .B1(n40131), .Y(
        n18097) );
  OAI211XL U42027 ( .A0(n34048), .A1(n42802), .B0(n18073), .C0(n18074), .Y(
        n36197) );
  OA22XL U42028 ( .A0(net262912), .A1(n34032), .B0(n34040), .B1(n40101), .Y(
        n18073) );
  OAI211XL U42029 ( .A0(n34040), .A1(n42803), .B0(n18049), .C0(n18050), .Y(
        n36189) );
  OA22XL U42030 ( .A0(net262912), .A1(n34024), .B0(n34032), .B1(n40101), .Y(
        n18049) );
  OAI211XL U42031 ( .A0(n34032), .A1(n42804), .B0(n18025), .C0(n18026), .Y(
        n36181) );
  OA22XL U42032 ( .A0(net262722), .A1(n34016), .B0(n34024), .B1(n40092), .Y(
        n18025) );
  OAI211XL U42033 ( .A0(n34024), .A1(n42805), .B0(n18001), .C0(n18002), .Y(
        n36173) );
  OA22XL U42034 ( .A0(net262665), .A1(n34008), .B0(n34016), .B1(n40072), .Y(
        n18001) );
  OAI211XL U42035 ( .A0(n34016), .A1(n42806), .B0(n17977), .C0(n17978), .Y(
        n36165) );
  OA22XL U42036 ( .A0(net262665), .A1(n34000), .B0(n34008), .B1(n40111), .Y(
        n17977) );
  OAI211XL U42037 ( .A0(n34008), .A1(n42808), .B0(n17953), .C0(n17954), .Y(
        n36157) );
  OA22XL U42038 ( .A0(net218304), .A1(n33992), .B0(n34000), .B1(n40111), .Y(
        n17953) );
  OAI211XL U42039 ( .A0(n34000), .A1(n42809), .B0(n17929), .C0(n17930), .Y(
        n36149) );
  OA22XL U42040 ( .A0(net218400), .A1(n33984), .B0(n33992), .B1(n40110), .Y(
        n17929) );
  OAI211XL U42041 ( .A0(n33728), .A1(n42751), .B0(n17113), .C0(n17114), .Y(
        n35877) );
  OA22XL U42042 ( .A0(net261886), .A1(n33712), .B0(n33720), .B1(n40149), .Y(
        n17113) );
  OAI211XL U42043 ( .A0(n33720), .A1(n42752), .B0(n17089), .C0(n17090), .Y(
        n35869) );
  OA22XL U42044 ( .A0(net261905), .A1(n33704), .B0(n33712), .B1(n40149), .Y(
        n17089) );
  OAI211XL U42045 ( .A0(n33712), .A1(n42753), .B0(n17065), .C0(n17066), .Y(
        n35861) );
  OA22XL U42046 ( .A0(net261905), .A1(n33696), .B0(n33704), .B1(n40148), .Y(
        n17065) );
  OAI211XL U42047 ( .A0(n33704), .A1(n42754), .B0(n17041), .C0(n17042), .Y(
        n35853) );
  OA22XL U42048 ( .A0(net261924), .A1(n33688), .B0(n33696), .B1(n40148), .Y(
        n17041) );
  OAI211XL U42049 ( .A0(n33696), .A1(n42755), .B0(n17017), .C0(n17018), .Y(
        n35845) );
  OA22XL U42050 ( .A0(net261924), .A1(n33680), .B0(n33688), .B1(n40147), .Y(
        n17017) );
  OAI211XL U42051 ( .A0(n33688), .A1(n42756), .B0(n16993), .C0(n16994), .Y(
        n35837) );
  OA22XL U42052 ( .A0(net261943), .A1(n33672), .B0(n33680), .B1(n40147), .Y(
        n16993) );
  OAI211XL U42053 ( .A0(n33680), .A1(n42758), .B0(n16969), .C0(n16970), .Y(
        n35829) );
  OA22XL U42054 ( .A0(net261943), .A1(n33664), .B0(n33672), .B1(n40146), .Y(
        n16969) );
  OAI211XL U42055 ( .A0(n33672), .A1(n42759), .B0(n16945), .C0(n16946), .Y(
        n35821) );
  OA22XL U42056 ( .A0(net218578), .A1(n33656), .B0(n33664), .B1(n40146), .Y(
        n16945) );
  OAI211XL U42057 ( .A0(n33664), .A1(n42760), .B0(n16921), .C0(n16922), .Y(
        n35813) );
  OA22XL U42058 ( .A0(net218500), .A1(n33648), .B0(n33656), .B1(n40145), .Y(
        n16921) );
  OAI211XL U42059 ( .A0(n33656), .A1(n42761), .B0(n16897), .C0(n16898), .Y(
        n35805) );
  OA22XL U42060 ( .A0(net261981), .A1(n33640), .B0(n33648), .B1(n40145), .Y(
        n16897) );
  OAI211XL U42061 ( .A0(n33648), .A1(n42762), .B0(n16873), .C0(n16874), .Y(
        n35797) );
  OA22XL U42062 ( .A0(net262323), .A1(n33632), .B0(n33640), .B1(n40127), .Y(
        n16873) );
  OAI211XL U42063 ( .A0(n33640), .A1(n42763), .B0(n16849), .C0(n16850), .Y(
        n35789) );
  OA22XL U42064 ( .A0(net262266), .A1(n33624), .B0(n33632), .B1(n40130), .Y(
        n16849) );
  OAI211XL U42065 ( .A0(n33632), .A1(n42765), .B0(n16825), .C0(n16826), .Y(
        n35781) );
  OA22XL U42066 ( .A0(net262266), .A1(n33616), .B0(n33624), .B1(n40129), .Y(
        n16825) );
  OAI211XL U42067 ( .A0(n33624), .A1(n42766), .B0(n16801), .C0(n16802), .Y(
        n35773) );
  OA22XL U42068 ( .A0(net262266), .A1(n33608), .B0(n33616), .B1(n40129), .Y(
        n16801) );
  OAI211XL U42069 ( .A0(n33568), .A1(n42742), .B0(n16633), .C0(n16634), .Y(
        n35717) );
  OA22XL U42070 ( .A0(net262342), .A1(n33552), .B0(n33560), .B1(n40126), .Y(
        n16633) );
  OAI211XL U42071 ( .A0(n33560), .A1(n42743), .B0(n16609), .C0(n16610), .Y(
        n35709) );
  OA22XL U42072 ( .A0(net262342), .A1(n33544), .B0(n33552), .B1(n40126), .Y(
        n16609) );
  OAI211XL U42073 ( .A0(n33552), .A1(n42744), .B0(n16585), .C0(n16586), .Y(
        n35701) );
  OA22XL U42074 ( .A0(net262361), .A1(n33536), .B0(n33544), .B1(n40125), .Y(
        n16585) );
  OAI211XL U42075 ( .A0(n33544), .A1(n42745), .B0(n16561), .C0(n16562), .Y(
        n35693) );
  OA22XL U42076 ( .A0(net262361), .A1(n33528), .B0(n33536), .B1(n40125), .Y(
        n16561) );
  OAI211XL U42077 ( .A0(n33536), .A1(n42746), .B0(n16537), .C0(n16538), .Y(
        n35685) );
  OA22XL U42078 ( .A0(net262361), .A1(n33520), .B0(n33528), .B1(n40124), .Y(
        n16537) );
  OAI211XL U42079 ( .A0(n33528), .A1(n42747), .B0(n16513), .C0(n16514), .Y(
        n35677) );
  OA22XL U42080 ( .A0(net262380), .A1(n33512), .B0(n33520), .B1(n40124), .Y(
        n16513) );
  OAI211XL U42081 ( .A0(n33520), .A1(n42749), .B0(n16489), .C0(n16490), .Y(
        n35669) );
  OA22XL U42082 ( .A0(net262114), .A1(n33504), .B0(n33512), .B1(n40138), .Y(
        n16489) );
  OAI211XL U42083 ( .A0(n33512), .A1(n42750), .B0(n16465), .C0(n16466), .Y(
        n35661) );
  OA22XL U42084 ( .A0(net262133), .A1(n33496), .B0(n33504), .B1(n40138), .Y(
        n16465) );
  OAI211XL U42085 ( .A0(n33504), .A1(n42783), .B0(n16441), .C0(n16442), .Y(
        n35653) );
  OA22XL U42086 ( .A0(net262133), .A1(n33488), .B0(n33496), .B1(n40137), .Y(
        n16441) );
  OAI211XL U42087 ( .A0(n33496), .A1(n42784), .B0(n16417), .C0(n16418), .Y(
        n35645) );
  OA22XL U42088 ( .A0(net262133), .A1(n33480), .B0(n33488), .B1(n40137), .Y(
        n16417) );
  OAI211XL U42089 ( .A0(n33488), .A1(n42785), .B0(n16393), .C0(n16394), .Y(
        n35637) );
  OA22XL U42090 ( .A0(net262152), .A1(n33472), .B0(n33480), .B1(n40136), .Y(
        n16393) );
  OAI211XL U42091 ( .A0(n33480), .A1(n42786), .B0(n16369), .C0(n16370), .Y(
        n35629) );
  OA22XL U42092 ( .A0(net262152), .A1(n33464), .B0(n33472), .B1(n40136), .Y(
        n16369) );
  OAI211XL U42093 ( .A0(n33472), .A1(n42788), .B0(n16345), .C0(n16346), .Y(
        n35621) );
  OA22XL U42094 ( .A0(net262171), .A1(n33456), .B0(n33464), .B1(n40135), .Y(
        n16345) );
  OAI211XL U42095 ( .A0(n33464), .A1(n42789), .B0(n16321), .C0(n16322), .Y(
        n35613) );
  OA22XL U42096 ( .A0(net262171), .A1(n33448), .B0(n33456), .B1(n40135), .Y(
        n16321) );
  OAI211XL U42097 ( .A0(n33456), .A1(n42790), .B0(n16297), .C0(n16298), .Y(
        n35605) );
  OA22XL U42098 ( .A0(net262190), .A1(n33440), .B0(n33448), .B1(n40134), .Y(
        n16297) );
  OAI211XL U42099 ( .A0(n33448), .A1(n42791), .B0(n16273), .C0(n16274), .Y(
        n35597) );
  OA22XL U42100 ( .A0(net262190), .A1(n33432), .B0(n33440), .B1(n40134), .Y(
        n16273) );
  OAI211XL U42101 ( .A0(n33440), .A1(n42792), .B0(n16249), .C0(n16250), .Y(
        n35589) );
  OA22XL U42102 ( .A0(net262209), .A1(n33424), .B0(n33432), .B1(n40133), .Y(
        n16249) );
  OAI211XL U42103 ( .A0(n33432), .A1(n42793), .B0(n16225), .C0(n16226), .Y(
        n35581) );
  OA22XL U42104 ( .A0(net262209), .A1(n33416), .B0(n33424), .B1(n40133), .Y(
        n16225) );
  OAI211XL U42105 ( .A0(n33424), .A1(n42795), .B0(n16201), .C0(n16202), .Y(
        n35573) );
  OA22XL U42106 ( .A0(net262209), .A1(n33408), .B0(n33416), .B1(n40132), .Y(
        n16201) );
  OAI211XL U42107 ( .A0(n33416), .A1(n42796), .B0(n16177), .C0(n16178), .Y(
        n35565) );
  OA22XL U42108 ( .A0(net262228), .A1(n33400), .B0(n33408), .B1(n40132), .Y(
        n16177) );
  OAI211XL U42109 ( .A0(n33408), .A1(n42797), .B0(n16153), .C0(n16154), .Y(
        n35557) );
  OA22XL U42110 ( .A0(net262228), .A1(n33392), .B0(n33400), .B1(n40131), .Y(
        n16153) );
  OAI211XL U42111 ( .A0(n33400), .A1(n42798), .B0(n16129), .C0(n16130), .Y(
        n35549) );
  OA22XL U42112 ( .A0(net262247), .A1(n33384), .B0(n33392), .B1(n40131), .Y(
        n16129) );
  OAI211XL U42113 ( .A0(n33392), .A1(n42767), .B0(n16105), .C0(n16106), .Y(
        n35541) );
  OA22XL U42114 ( .A0(net218410), .A1(n33376), .B0(n33384), .B1(n40054), .Y(
        n16105) );
  OAI211XL U42115 ( .A0(n33384), .A1(n42768), .B0(n16081), .C0(n16082), .Y(
        n35533) );
  OA22XL U42116 ( .A0(net263615), .A1(n33368), .B0(n33376), .B1(n40061), .Y(
        n16081) );
  OAI211XL U42117 ( .A0(n33376), .A1(n42769), .B0(n16057), .C0(n16058), .Y(
        n35525) );
  OA22XL U42118 ( .A0(net263615), .A1(n33360), .B0(n33368), .B1(n40060), .Y(
        n16057) );
  OAI211XL U42119 ( .A0(n33368), .A1(n42770), .B0(n16033), .C0(n16034), .Y(
        n35517) );
  OA22XL U42120 ( .A0(net263634), .A1(n33352), .B0(n33360), .B1(n40060), .Y(
        n16033) );
  OAI211XL U42121 ( .A0(n33360), .A1(n42771), .B0(n16009), .C0(n16010), .Y(
        n35509) );
  OA22XL U42122 ( .A0(net263634), .A1(n33344), .B0(n33352), .B1(n40059), .Y(
        n16009) );
  OAI211XL U42123 ( .A0(n33352), .A1(n42773), .B0(n15985), .C0(n15986), .Y(
        n35501) );
  OA22XL U42124 ( .A0(net263634), .A1(n33336), .B0(n33344), .B1(n40059), .Y(
        n15985) );
  OAI211XL U42125 ( .A0(n33344), .A1(n42774), .B0(n15961), .C0(n15962), .Y(
        n35493) );
  OA22XL U42126 ( .A0(net263653), .A1(n33328), .B0(n33336), .B1(n40058), .Y(
        n15961) );
  OAI211XL U42127 ( .A0(n33336), .A1(n42775), .B0(n15937), .C0(n15938), .Y(
        n35485) );
  OA22XL U42128 ( .A0(net263653), .A1(n33320), .B0(n33328), .B1(n40058), .Y(
        n15937) );
  OAI211XL U42129 ( .A0(n33328), .A1(n42776), .B0(n15913), .C0(n15914), .Y(
        n35477) );
  OA22XL U42130 ( .A0(net263672), .A1(n33312), .B0(n33320), .B1(n40138), .Y(
        n15913) );
  OAI211XL U42131 ( .A0(n33320), .A1(n42777), .B0(n15889), .C0(n15890), .Y(
        n35469) );
  OA22XL U42132 ( .A0(net263672), .A1(n33304), .B0(n33312), .B1(n40137), .Y(
        n15889) );
  OAI211XL U42133 ( .A0(n33312), .A1(n42778), .B0(n15865), .C0(n15866), .Y(
        n35461) );
  OA22XL U42134 ( .A0(net263691), .A1(n33296), .B0(n33304), .B1(n40057), .Y(
        n15865) );
  OAI211XL U42135 ( .A0(n33304), .A1(n42780), .B0(n15841), .C0(n15842), .Y(
        n35453) );
  OA22XL U42136 ( .A0(net263691), .A1(n33288), .B0(n33296), .B1(n40057), .Y(
        n15841) );
  OAI211XL U42137 ( .A0(n33296), .A1(n42781), .B0(n15817), .C0(n15818), .Y(
        n35445) );
  OA22XL U42138 ( .A0(net263710), .A1(n33280), .B0(n33288), .B1(n40056), .Y(
        n15817) );
  OAI211XL U42139 ( .A0(n33288), .A1(n42782), .B0(n15793), .C0(n15794), .Y(
        n35437) );
  OA22XL U42140 ( .A0(net263710), .A1(n33272), .B0(n33280), .B1(n40056), .Y(
        n15793) );
  OAI211XL U42141 ( .A0(n33280), .A1(n42944), .B0(n15769), .C0(n15770), .Y(
        n35429) );
  OA22XL U42142 ( .A0(net263710), .A1(n33264), .B0(n33272), .B1(n40055), .Y(
        n15769) );
  OAI211XL U42143 ( .A0(n33272), .A1(n42945), .B0(n15745), .C0(n15746), .Y(
        n35421) );
  OA22XL U42144 ( .A0(net218468), .A1(n33256), .B0(n33264), .B1(n40055), .Y(
        n15745) );
  OAI211XL U42145 ( .A0(n33264), .A1(n42946), .B0(n15721), .C0(n15722), .Y(
        n35413) );
  OA22XL U42146 ( .A0(net263539), .A1(n33248), .B0(n33256), .B1(n40065), .Y(
        n15721) );
  OAI211XL U42147 ( .A0(n33256), .A1(n42947), .B0(n15697), .C0(n15698), .Y(
        n35405) );
  OA22XL U42148 ( .A0(net263159), .A1(n33240), .B0(n33248), .B1(n40069), .Y(
        n15697) );
  OAI211XL U42149 ( .A0(n33248), .A1(n42948), .B0(n15673), .C0(n15674), .Y(
        n35397) );
  OA22XL U42150 ( .A0(net218414), .A1(n33232), .B0(n33240), .B1(n40068), .Y(
        n15673) );
  OAI211XL U42151 ( .A0(n33240), .A1(n42949), .B0(n15649), .C0(n15650), .Y(
        n35389) );
  OA22XL U42152 ( .A0(net218376), .A1(n33224), .B0(n33232), .B1(n40068), .Y(
        n15649) );
  OAI211XL U42153 ( .A0(n33232), .A1(n42951), .B0(n15625), .C0(n15626), .Y(
        n35381) );
  OA22XL U42154 ( .A0(net263501), .A1(n33216), .B0(n33224), .B1(n40067), .Y(
        n15625) );
  OAI211XL U42155 ( .A0(n33224), .A1(n42952), .B0(n15601), .C0(n15602), .Y(
        n35373) );
  OA22XL U42156 ( .A0(net263501), .A1(n33208), .B0(n33216), .B1(n40067), .Y(
        n15601) );
  OAI211XL U42157 ( .A0(n33216), .A1(n42953), .B0(n15577), .C0(n15578), .Y(
        n35365) );
  OA22XL U42158 ( .A0(net218304), .A1(n33200), .B0(n33208), .B1(n40066), .Y(
        n15577) );
  OAI211XL U42159 ( .A0(n33208), .A1(n42954), .B0(n15553), .C0(n15554), .Y(
        n35357) );
  OA22XL U42160 ( .A0(net218490), .A1(n33192), .B0(n33200), .B1(n40066), .Y(
        n15553) );
  OAI211XL U42161 ( .A0(n33200), .A1(n42955), .B0(n15529), .C0(n15530), .Y(
        n35349) );
  OA22XL U42162 ( .A0(net263539), .A1(n33184), .B0(n33192), .B1(n40065), .Y(
        n15529) );
  OAI211XL U42163 ( .A0(n33192), .A1(n42956), .B0(n15505), .C0(n15506), .Y(
        n35341) );
  OA22XL U42164 ( .A0(net263539), .A1(n33176), .B0(n33184), .B1(n40065), .Y(
        n15505) );
  OAI211XL U42165 ( .A0(n33184), .A1(n42958), .B0(n15481), .C0(n15482), .Y(
        n35333) );
  OA22XL U42166 ( .A0(net263558), .A1(n33168), .B0(n33176), .B1(n40064), .Y(
        n15481) );
  OAI211XL U42167 ( .A0(n33176), .A1(n42959), .B0(n15457), .C0(n15458), .Y(
        n35325) );
  OA22XL U42168 ( .A0(net263558), .A1(n33160), .B0(n33168), .B1(n40064), .Y(
        n15457) );
  OAI211XL U42169 ( .A0(n33168), .A1(n42928), .B0(n15433), .C0(n15434), .Y(
        n35317) );
  OA22XL U42170 ( .A0(net263577), .A1(n33152), .B0(n33160), .B1(n40063), .Y(
        n15433) );
  OAI211XL U42171 ( .A0(n33160), .A1(n42929), .B0(n15409), .C0(n15410), .Y(
        n35309) );
  OA22XL U42172 ( .A0(net263577), .A1(n33144), .B0(n33152), .B1(n40063), .Y(
        n15409) );
  OAI211XL U42173 ( .A0(n33152), .A1(n42930), .B0(n15385), .C0(n15386), .Y(
        n35301) );
  OA22XL U42174 ( .A0(net263577), .A1(n33136), .B0(n33144), .B1(n40062), .Y(
        n15385) );
  OAI211XL U42175 ( .A0(n33144), .A1(n42931), .B0(n15361), .C0(n15362), .Y(
        n35293) );
  OA22XL U42176 ( .A0(net263596), .A1(n33128), .B0(n33136), .B1(n40062), .Y(
        n15361) );
  OAI211XL U42177 ( .A0(n33136), .A1(n42932), .B0(n15337), .C0(n15338), .Y(
        n35285) );
  OA22XL U42178 ( .A0(net218458), .A1(n33120), .B0(n33128), .B1(n40062), .Y(
        n15337) );
  OAI211XL U42179 ( .A0(n33128), .A1(n42933), .B0(n15313), .C0(n15314), .Y(
        n35277) );
  OA22XL U42180 ( .A0(net263881), .A1(n33112), .B0(n33120), .B1(n40046), .Y(
        n15313) );
  OAI211XL U42181 ( .A0(n33120), .A1(n42934), .B0(n15289), .C0(n15290), .Y(
        n35269) );
  OA22XL U42182 ( .A0(net263881), .A1(n33104), .B0(n33112), .B1(n40045), .Y(
        n15289) );
  OAI211XL U42183 ( .A0(n33112), .A1(n42936), .B0(n15265), .C0(n15266), .Y(
        n35261) );
  OA22XL U42184 ( .A0(net263900), .A1(n33096), .B0(n33104), .B1(n40045), .Y(
        n15265) );
  OAI211XL U42185 ( .A0(n33104), .A1(n42937), .B0(n15241), .C0(n15242), .Y(
        n35253) );
  OA22XL U42186 ( .A0(net263900), .A1(n33088), .B0(n33096), .B1(n40044), .Y(
        n15241) );
  OAI211XL U42187 ( .A0(n33096), .A1(n42938), .B0(n15217), .C0(n15218), .Y(
        n35245) );
  OA22XL U42188 ( .A0(net263919), .A1(n33080), .B0(n33088), .B1(n40044), .Y(
        n15217) );
  OAI211XL U42189 ( .A0(n33088), .A1(n42939), .B0(n15193), .C0(n15194), .Y(
        n35237) );
  OA22XL U42190 ( .A0(net263919), .A1(n33072), .B0(n33080), .B1(n40043), .Y(
        n15193) );
  OAI211XL U42191 ( .A0(n33080), .A1(n42940), .B0(n15169), .C0(n15170), .Y(
        n35229) );
  OA22XL U42192 ( .A0(net262190), .A1(n33064), .B0(n33072), .B1(n40043), .Y(
        n15169) );
  OAI211XL U42193 ( .A0(n33072), .A1(n42941), .B0(n15145), .C0(n15146), .Y(
        n35221) );
  OA22XL U42194 ( .A0(net218442), .A1(n33056), .B0(n33064), .B1(n40072), .Y(
        n15145) );
  OAI211XL U42195 ( .A0(n33064), .A1(n42943), .B0(n15121), .C0(n15122), .Y(
        n35213) );
  OA22XL U42196 ( .A0(net263957), .A1(n33048), .B0(n33056), .B1(n40062), .Y(
        n15121) );
  OAI211XL U42197 ( .A0(n33056), .A1(n42976), .B0(n15097), .C0(n15098), .Y(
        n35205) );
  OA22XL U42198 ( .A0(net263957), .A1(n33040), .B0(n33048), .B1(n40042), .Y(
        n15097) );
  OAI211XL U42199 ( .A0(n33048), .A1(n42977), .B0(n15073), .C0(n15074), .Y(
        n35197) );
  OA22XL U42200 ( .A0(net263957), .A1(n33032), .B0(n33040), .B1(n40042), .Y(
        n15073) );
  OAI211XL U42201 ( .A0(n33040), .A1(n42978), .B0(n15049), .C0(n15050), .Y(
        n35189) );
  OA22XL U42202 ( .A0(net263976), .A1(n33024), .B0(n33032), .B1(n40041), .Y(
        n15049) );
  OAI211XL U42203 ( .A0(n33032), .A1(n42979), .B0(n15025), .C0(n15026), .Y(
        n35181) );
  OA22XL U42204 ( .A0(net263976), .A1(n33016), .B0(n33024), .B1(n40041), .Y(
        n15025) );
  OAI211XL U42205 ( .A0(n33024), .A1(n42980), .B0(n15001), .C0(n15002), .Y(
        n35173) );
  OA22XL U42206 ( .A0(net263995), .A1(n33008), .B0(n33016), .B1(n40040), .Y(
        n15001) );
  OAI211XL U42207 ( .A0(n33016), .A1(n42982), .B0(n14977), .C0(n14978), .Y(
        n35165) );
  OA22XL U42208 ( .A0(net263995), .A1(n33000), .B0(n33008), .B1(n40040), .Y(
        n14977) );
  OAI211XL U42209 ( .A0(n33008), .A1(n42983), .B0(n14953), .C0(n14954), .Y(
        n35157) );
  OA22XL U42210 ( .A0(net218398), .A1(n32992), .B0(n33000), .B1(n40054), .Y(
        n14953) );
  OAI211XL U42211 ( .A0(n33000), .A1(n42984), .B0(n14929), .C0(n14930), .Y(
        n35149) );
  OA22XL U42212 ( .A0(net263748), .A1(n32984), .B0(n32992), .B1(n40054), .Y(
        n14929) );
  OA22XL U42213 ( .A0(net263767), .A1(n32968), .B0(n32976), .B1(n40053), .Y(
        n14881) );
  OA22XL U42214 ( .A0(net263292), .A1(net219468), .B0(n32408), .B1(n40079),
        .Y(n13177) );
  OA22XL U42215 ( .A0(net263292), .A1(n42592), .B0(net219434), .B1(n40079),
        .Y(n13153) );
  OAI211XL U42216 ( .A0(n34065), .A1(n42799), .B0(n18124), .C0(n18125), .Y(
        n36214) );
  OA22XL U42217 ( .A0(net262893), .A1(n34049), .B0(n34057), .B1(net218664),
        .Y(n18124) );
  OAI211XL U42218 ( .A0(n34057), .A1(n42800), .B0(n18100), .C0(n18101), .Y(
        n36206) );
  OA22XL U42219 ( .A0(net262893), .A1(n34041), .B0(n34049), .B1(net218674),
        .Y(n18100) );
  OAI211XL U42220 ( .A0(n34049), .A1(n42802), .B0(n18076), .C0(n18077), .Y(
        n36198) );
  OA22XL U42221 ( .A0(net262912), .A1(n34033), .B0(n34041), .B1(n40101), .Y(
        n18076) );
  OAI211XL U42222 ( .A0(n34041), .A1(n42803), .B0(n18052), .C0(n18053), .Y(
        n36190) );
  OA22XL U42223 ( .A0(net262912), .A1(n34025), .B0(n34033), .B1(n40101), .Y(
        n18052) );
  OAI211XL U42224 ( .A0(n34033), .A1(n42804), .B0(n18028), .C0(n18029), .Y(
        n36182) );
  OA22XL U42225 ( .A0(net262931), .A1(n34017), .B0(n34025), .B1(n40100), .Y(
        n18028) );
  OAI211XL U42226 ( .A0(n34025), .A1(n42805), .B0(n18004), .C0(n18005), .Y(
        n36174) );
  OA22XL U42227 ( .A0(net262665), .A1(n34009), .B0(n34017), .B1(n40068), .Y(
        n18004) );
  OAI211XL U42228 ( .A0(n34017), .A1(n42806), .B0(n17980), .C0(n17981), .Y(
        n36166) );
  OA22XL U42229 ( .A0(net262665), .A1(n34001), .B0(n34009), .B1(n40111), .Y(
        n17980) );
  OAI211XL U42230 ( .A0(n34009), .A1(n42807), .B0(n17956), .C0(n17957), .Y(
        n36158) );
  OA22XL U42231 ( .A0(net218476), .A1(n33993), .B0(n34001), .B1(n40111), .Y(
        n17956) );
  OAI211XL U42232 ( .A0(n34001), .A1(n42809), .B0(n17932), .C0(n17933), .Y(
        n36150) );
  OA22XL U42233 ( .A0(net218506), .A1(n33985), .B0(n33993), .B1(n40110), .Y(
        n17932) );
  OAI211XL U42234 ( .A0(n33729), .A1(n42751), .B0(n17116), .C0(n17117), .Y(
        n35878) );
  OA22XL U42235 ( .A0(net261886), .A1(n33713), .B0(n33721), .B1(n40149), .Y(
        n17116) );
  OAI211XL U42236 ( .A0(n33721), .A1(n42752), .B0(n17092), .C0(n17093), .Y(
        n35870) );
  OA22XL U42237 ( .A0(net261905), .A1(n33705), .B0(n33713), .B1(n40149), .Y(
        n17092) );
  OAI211XL U42238 ( .A0(n33713), .A1(n42753), .B0(n17068), .C0(n17069), .Y(
        n35862) );
  OA22XL U42239 ( .A0(net261905), .A1(n33697), .B0(n33705), .B1(n40148), .Y(
        n17068) );
  OAI211XL U42240 ( .A0(n33705), .A1(n42754), .B0(n17044), .C0(n17045), .Y(
        n35854) );
  OA22XL U42241 ( .A0(net261924), .A1(n33689), .B0(n33697), .B1(n40148), .Y(
        n17044) );
  OAI211XL U42242 ( .A0(n33697), .A1(n42755), .B0(n17020), .C0(n17021), .Y(
        n35846) );
  OA22XL U42243 ( .A0(net261924), .A1(n33681), .B0(n33689), .B1(n40147), .Y(
        n17020) );
  OAI211XL U42244 ( .A0(n33689), .A1(n42756), .B0(n16996), .C0(n16997), .Y(
        n35838) );
  OA22XL U42245 ( .A0(net261943), .A1(n33673), .B0(n33681), .B1(n40147), .Y(
        n16996) );
  OAI211XL U42246 ( .A0(n33681), .A1(n42757), .B0(n16972), .C0(n16973), .Y(
        n35830) );
  OA22XL U42247 ( .A0(net261943), .A1(n33665), .B0(n33673), .B1(n40146), .Y(
        n16972) );
  OAI211XL U42248 ( .A0(n33673), .A1(n42759), .B0(n16948), .C0(n16949), .Y(
        n35822) );
  OA22XL U42249 ( .A0(net218482), .A1(n33657), .B0(n33665), .B1(n40146), .Y(
        n16948) );
  OAI211XL U42250 ( .A0(n33665), .A1(n42760), .B0(n16924), .C0(n16925), .Y(
        n35814) );
  OA22XL U42251 ( .A0(net218502), .A1(n33649), .B0(n33657), .B1(n40145), .Y(
        n16924) );
  OAI211XL U42252 ( .A0(n33657), .A1(n42761), .B0(n16900), .C0(n16901), .Y(
        n35806) );
  OA22XL U42253 ( .A0(net218454), .A1(n33641), .B0(n33649), .B1(n40145), .Y(
        n16900) );
  OAI211XL U42254 ( .A0(n33649), .A1(n42762), .B0(n16876), .C0(n16877), .Y(
        n35798) );
  OA22XL U42255 ( .A0(net261981), .A1(n33633), .B0(n33641), .B1(n40144), .Y(
        n16876) );
  OAI211XL U42256 ( .A0(n33641), .A1(n42763), .B0(n16852), .C0(n16853), .Y(
        n35790) );
  OA22XL U42257 ( .A0(net262266), .A1(n33625), .B0(n33633), .B1(n40130), .Y(
        n16852) );
  OAI211XL U42258 ( .A0(n33633), .A1(n42764), .B0(n16828), .C0(n16829), .Y(
        n35782) );
  OA22XL U42259 ( .A0(net262266), .A1(n33617), .B0(n33625), .B1(n40129), .Y(
        n16828) );
  OAI211XL U42260 ( .A0(n33625), .A1(n42766), .B0(n16804), .C0(n16805), .Y(
        n35774) );
  OA22XL U42261 ( .A0(net262266), .A1(n33609), .B0(n33617), .B1(n40129), .Y(
        n16804) );
  OAI211XL U42262 ( .A0(n33569), .A1(n42741), .B0(n16636), .C0(n16637), .Y(
        n35718) );
  OA22XL U42263 ( .A0(net262342), .A1(n33553), .B0(n33561), .B1(n40126), .Y(
        n16636) );
  OAI211XL U42264 ( .A0(n33561), .A1(n42743), .B0(n16612), .C0(n16613), .Y(
        n35710) );
  OA22XL U42265 ( .A0(net262342), .A1(n33545), .B0(n33553), .B1(n40126), .Y(
        n16612) );
  OAI211XL U42266 ( .A0(n33553), .A1(n42744), .B0(n16588), .C0(n16589), .Y(
        n35702) );
  OA22XL U42267 ( .A0(net262342), .A1(n33537), .B0(n33545), .B1(n40125), .Y(
        n16588) );
  OAI211XL U42268 ( .A0(n33545), .A1(n42745), .B0(n16564), .C0(n16565), .Y(
        n35694) );
  OA22XL U42269 ( .A0(net262361), .A1(n33529), .B0(n33537), .B1(n40125), .Y(
        n16564) );
  OAI211XL U42270 ( .A0(n33537), .A1(n42746), .B0(n16540), .C0(n16541), .Y(
        n35686) );
  OA22XL U42271 ( .A0(net262361), .A1(n33521), .B0(n33529), .B1(n40124), .Y(
        n16540) );
  OAI211XL U42272 ( .A0(n33529), .A1(n42747), .B0(n16516), .C0(n16517), .Y(
        n35678) );
  OA22XL U42273 ( .A0(net262380), .A1(n33513), .B0(n33521), .B1(n40124), .Y(
        n16516) );
  OAI211XL U42274 ( .A0(n33521), .A1(n42748), .B0(n16492), .C0(n16493), .Y(
        n35670) );
  OA22XL U42275 ( .A0(net262190), .A1(n33505), .B0(n33513), .B1(n40134), .Y(
        n16492) );
  OAI211XL U42276 ( .A0(n33513), .A1(n42750), .B0(n16468), .C0(n16469), .Y(
        n35662) );
  OA22XL U42277 ( .A0(net262114), .A1(n33497), .B0(n33505), .B1(n40138), .Y(
        n16468) );
  OAI211XL U42278 ( .A0(n33505), .A1(n42783), .B0(n16444), .C0(n16445), .Y(
        n35654) );
  OA22XL U42279 ( .A0(net262133), .A1(n33489), .B0(n33497), .B1(n40137), .Y(
        n16444) );
  OAI211XL U42280 ( .A0(n33497), .A1(n42784), .B0(n16420), .C0(n16421), .Y(
        n35646) );
  OA22XL U42281 ( .A0(net262133), .A1(n33481), .B0(n33489), .B1(n40137), .Y(
        n16420) );
  OAI211XL U42282 ( .A0(n33489), .A1(n42785), .B0(n16396), .C0(n16397), .Y(
        n35638) );
  OA22XL U42283 ( .A0(net262152), .A1(n33473), .B0(n33481), .B1(n40136), .Y(
        n16396) );
  OAI211XL U42284 ( .A0(n33481), .A1(n42786), .B0(n16372), .C0(n16373), .Y(
        n35630) );
  OA22XL U42285 ( .A0(net262152), .A1(n33465), .B0(n33473), .B1(n40136), .Y(
        n16372) );
  OAI211XL U42286 ( .A0(n33473), .A1(n42787), .B0(n16348), .C0(n16349), .Y(
        n35622) );
  OA22XL U42287 ( .A0(net262171), .A1(n33457), .B0(n33465), .B1(n40135), .Y(
        n16348) );
  OAI211XL U42288 ( .A0(n33465), .A1(n42789), .B0(n16324), .C0(n16325), .Y(
        n35614) );
  OA22XL U42289 ( .A0(net262171), .A1(n33449), .B0(n33457), .B1(n40135), .Y(
        n16324) );
  OAI211XL U42290 ( .A0(n33457), .A1(n42790), .B0(n16300), .C0(n16301), .Y(
        n35606) );
  OA22XL U42291 ( .A0(net262190), .A1(n33441), .B0(n33449), .B1(n40134), .Y(
        n16300) );
  OAI211XL U42292 ( .A0(n33449), .A1(n42791), .B0(n16276), .C0(n16277), .Y(
        n35598) );
  OA22XL U42293 ( .A0(net262190), .A1(n33433), .B0(n33441), .B1(n40134), .Y(
        n16276) );
  OAI211XL U42294 ( .A0(n33441), .A1(n42792), .B0(n16252), .C0(n16253), .Y(
        n35590) );
  OA22XL U42295 ( .A0(net262209), .A1(n33425), .B0(n33433), .B1(n40133), .Y(
        n16252) );
  OAI211XL U42296 ( .A0(n33433), .A1(n42793), .B0(n16228), .C0(n16229), .Y(
        n35582) );
  OA22XL U42297 ( .A0(net262209), .A1(n33417), .B0(n33425), .B1(n40133), .Y(
        n16228) );
  OAI211XL U42298 ( .A0(n33425), .A1(n42794), .B0(n16204), .C0(n16205), .Y(
        n35574) );
  OA22XL U42299 ( .A0(net262209), .A1(n33409), .B0(n33417), .B1(n40132), .Y(
        n16204) );
  OAI211XL U42300 ( .A0(n33417), .A1(n42796), .B0(n16180), .C0(n16181), .Y(
        n35566) );
  OA22XL U42301 ( .A0(net262228), .A1(n33401), .B0(n33409), .B1(n40132), .Y(
        n16180) );
  OAI211XL U42302 ( .A0(n33409), .A1(n42797), .B0(n16156), .C0(n16157), .Y(
        n35558) );
  OA22XL U42303 ( .A0(net262228), .A1(n33393), .B0(n33401), .B1(n40131), .Y(
        n16156) );
  OAI211XL U42304 ( .A0(n33401), .A1(n42798), .B0(n16132), .C0(n16133), .Y(
        n35550) );
  OA22XL U42305 ( .A0(net262247), .A1(n33385), .B0(n33393), .B1(n40131), .Y(
        n16132) );
  OAI211XL U42306 ( .A0(n33393), .A1(n42767), .B0(n16108), .C0(n16109), .Y(
        n35542) );
  OA22XL U42307 ( .A0(net262380), .A1(n33377), .B0(n33385), .B1(n40123), .Y(
        n16108) );
  OAI211XL U42308 ( .A0(n33385), .A1(n42768), .B0(n16084), .C0(n16085), .Y(
        n35534) );
  OA22XL U42309 ( .A0(net263615), .A1(n33369), .B0(n33377), .B1(n40061), .Y(
        n16084) );
  OAI211XL U42310 ( .A0(n33377), .A1(n42769), .B0(n16060), .C0(n16061), .Y(
        n35526) );
  OA22XL U42311 ( .A0(net263615), .A1(n33361), .B0(n33369), .B1(n40060), .Y(
        n16060) );
  OAI211XL U42312 ( .A0(n33369), .A1(n42770), .B0(n16036), .C0(n16037), .Y(
        n35518) );
  OA22XL U42313 ( .A0(net263615), .A1(n33353), .B0(n33361), .B1(n40060), .Y(
        n16036) );
  OAI211XL U42314 ( .A0(n33361), .A1(n42771), .B0(n16012), .C0(n16013), .Y(
        n35510) );
  OA22XL U42315 ( .A0(net263634), .A1(n33345), .B0(n33353), .B1(n40059), .Y(
        n16012) );
  OAI211XL U42316 ( .A0(n33353), .A1(n42772), .B0(n15988), .C0(n15989), .Y(
        n35502) );
  OA22XL U42317 ( .A0(net263634), .A1(n33337), .B0(n33345), .B1(n40059), .Y(
        n15988) );
  OAI211XL U42318 ( .A0(n33345), .A1(n42774), .B0(n15964), .C0(n15965), .Y(
        n35494) );
  OA22XL U42319 ( .A0(net263653), .A1(n33329), .B0(n33337), .B1(n40058), .Y(
        n15964) );
  OAI211XL U42320 ( .A0(n33337), .A1(n42775), .B0(n15940), .C0(n15941), .Y(
        n35486) );
  OA22XL U42321 ( .A0(net263653), .A1(n33321), .B0(n33329), .B1(n40058), .Y(
        n15940) );
  OAI211XL U42322 ( .A0(n33329), .A1(n42776), .B0(n15916), .C0(n15917), .Y(
        n35478) );
  OA22XL U42323 ( .A0(net263672), .A1(n33313), .B0(n33321), .B1(net218642),
        .Y(n15916) );
  OAI211XL U42324 ( .A0(n33321), .A1(n42777), .B0(n15892), .C0(n15893), .Y(
        n35470) );
  OA22XL U42325 ( .A0(net263672), .A1(n33305), .B0(n33313), .B1(n40068), .Y(
        n15892) );
  OAI211XL U42326 ( .A0(n33313), .A1(n42778), .B0(n15868), .C0(n15869), .Y(
        n35462) );
  OA22XL U42327 ( .A0(net263691), .A1(n33297), .B0(n33305), .B1(n40057), .Y(
        n15868) );
  OAI211XL U42328 ( .A0(n33305), .A1(n42779), .B0(n15844), .C0(n15845), .Y(
        n35454) );
  OA22XL U42329 ( .A0(net263691), .A1(n33289), .B0(n33297), .B1(n40057), .Y(
        n15844) );
  OAI211XL U42330 ( .A0(n33297), .A1(n42781), .B0(n15820), .C0(n15821), .Y(
        n35446) );
  OA22XL U42331 ( .A0(net263710), .A1(n33281), .B0(n33289), .B1(n40056), .Y(
        n15820) );
  OAI211XL U42332 ( .A0(n33289), .A1(n42782), .B0(n15796), .C0(n15797), .Y(
        n35438) );
  OA22XL U42333 ( .A0(net263710), .A1(n33273), .B0(n33281), .B1(n40056), .Y(
        n15796) );
  OAI211XL U42334 ( .A0(n33281), .A1(n42952), .B0(n15772), .C0(n15773), .Y(
        n35430) );
  OA22XL U42335 ( .A0(net263710), .A1(n33265), .B0(n33273), .B1(n40055), .Y(
        n15772) );
  OAI211XL U42336 ( .A0(n33273), .A1(n42945), .B0(n15748), .C0(n15749), .Y(
        n35422) );
  OA22XL U42337 ( .A0(net218370), .A1(n33257), .B0(n33265), .B1(n40055), .Y(
        n15748) );
  OAI211XL U42338 ( .A0(n33265), .A1(n42946), .B0(n15724), .C0(n15725), .Y(
        n35414) );
  OA22XL U42339 ( .A0(net218392), .A1(n33249), .B0(n33257), .B1(n40054), .Y(
        n15724) );
  OAI211XL U42340 ( .A0(n33257), .A1(n42947), .B0(n15700), .C0(n15701), .Y(
        n35406) );
  OA22XL U42341 ( .A0(net218428), .A1(n33241), .B0(n33249), .B1(n40069), .Y(
        n15700) );
  OAI211XL U42342 ( .A0(n33249), .A1(n42948), .B0(n15676), .C0(n15677), .Y(
        n35398) );
  OA22XL U42343 ( .A0(net263045), .A1(n33233), .B0(n33241), .B1(n40068), .Y(
        n15676) );
  OAI211XL U42344 ( .A0(n33241), .A1(n42949), .B0(n15652), .C0(n15653), .Y(
        n35390) );
  OA22XL U42345 ( .A0(net218430), .A1(n33225), .B0(n33233), .B1(n40068), .Y(
        n15652) );
  OAI211XL U42346 ( .A0(n33233), .A1(n42950), .B0(n15628), .C0(n15629), .Y(
        n35382) );
  OA22XL U42347 ( .A0(net263501), .A1(n33217), .B0(n33225), .B1(n40067), .Y(
        n15628) );
  OAI211XL U42348 ( .A0(n33225), .A1(n42952), .B0(n15604), .C0(n15605), .Y(
        n35374) );
  OA22XL U42349 ( .A0(net263501), .A1(n33209), .B0(n33217), .B1(n40067), .Y(
        n15604) );
  OAI211XL U42350 ( .A0(n33217), .A1(n42953), .B0(n15580), .C0(n15581), .Y(
        n35366) );
  OA22XL U42351 ( .A0(net218424), .A1(n33201), .B0(n33209), .B1(n40066), .Y(
        n15580) );
  OAI211XL U42352 ( .A0(n33209), .A1(n42954), .B0(n15556), .C0(n15557), .Y(
        n35358) );
  OA22XL U42353 ( .A0(net218434), .A1(n33193), .B0(n33201), .B1(n40066), .Y(
        n15556) );
  OAI211XL U42354 ( .A0(n33201), .A1(n42955), .B0(n15532), .C0(n15533), .Y(
        n35350) );
  OA22XL U42355 ( .A0(net263539), .A1(n33185), .B0(n33193), .B1(n40065), .Y(
        n15532) );
  OAI211XL U42356 ( .A0(n33193), .A1(n42956), .B0(n15508), .C0(n15509), .Y(
        n35342) );
  OA22XL U42357 ( .A0(net263539), .A1(n33177), .B0(n33185), .B1(n40065), .Y(
        n15508) );
  OAI211XL U42358 ( .A0(n33185), .A1(n42957), .B0(n15484), .C0(n15485), .Y(
        n35334) );
  OA22XL U42359 ( .A0(net263558), .A1(n33169), .B0(n33177), .B1(n40064), .Y(
        n15484) );
  OAI211XL U42360 ( .A0(n33177), .A1(n42959), .B0(n15460), .C0(n15461), .Y(
        n35326) );
  OA22XL U42361 ( .A0(net263558), .A1(n33161), .B0(n33169), .B1(n40064), .Y(
        n15460) );
  OAI211XL U42362 ( .A0(n33169), .A1(n42935), .B0(n15436), .C0(n15437), .Y(
        n35318) );
  OA22XL U42363 ( .A0(net263558), .A1(n33153), .B0(n33161), .B1(n40063), .Y(
        n15436) );
  OAI211XL U42364 ( .A0(n33161), .A1(n42929), .B0(n15412), .C0(n15413), .Y(
        n35310) );
  OA22XL U42365 ( .A0(net263577), .A1(n33145), .B0(n33153), .B1(n40063), .Y(
        n15412) );
  OAI211XL U42366 ( .A0(n33153), .A1(n42930), .B0(n15388), .C0(n15389), .Y(
        n35302) );
  OA22XL U42367 ( .A0(net263577), .A1(n33137), .B0(n33145), .B1(n40062), .Y(
        n15388) );
  OAI211XL U42368 ( .A0(n33145), .A1(n42931), .B0(n15364), .C0(n15365), .Y(
        n35294) );
  OA22XL U42369 ( .A0(net263596), .A1(n33129), .B0(n33137), .B1(n40062), .Y(
        n15364) );
  OAI211XL U42370 ( .A0(n33137), .A1(n42932), .B0(n15340), .C0(n15341), .Y(
        n35286) );
  OA22XL U42371 ( .A0(net263596), .A1(n33121), .B0(n33129), .B1(n40061), .Y(
        n15340) );
  OAI211XL U42372 ( .A0(n33129), .A1(n42933), .B0(n15316), .C0(n15317), .Y(
        n35278) );
  OA22XL U42373 ( .A0(net263881), .A1(n33113), .B0(n33121), .B1(n40046), .Y(
        n15316) );
  OAI211XL U42374 ( .A0(n33121), .A1(n42934), .B0(n15292), .C0(n15293), .Y(
        n35270) );
  OA22XL U42375 ( .A0(net263881), .A1(n33105), .B0(n33113), .B1(n40045), .Y(
        n15292) );
  OAI211XL U42376 ( .A0(n33113), .A1(n42936), .B0(n15268), .C0(n15269), .Y(
        n35262) );
  OA22XL U42377 ( .A0(net263900), .A1(n33097), .B0(n33105), .B1(n40045), .Y(
        n15268) );
  OAI211XL U42378 ( .A0(n33105), .A1(n42937), .B0(n15244), .C0(n15245), .Y(
        n35254) );
  OA22XL U42379 ( .A0(net263900), .A1(n33089), .B0(n33097), .B1(n40044), .Y(
        n15244) );
  OAI211XL U42380 ( .A0(n33097), .A1(n42938), .B0(n15220), .C0(n15221), .Y(
        n35246) );
  OA22XL U42381 ( .A0(net263919), .A1(n33081), .B0(n33089), .B1(n40044), .Y(
        n15220) );
  OAI211XL U42382 ( .A0(n33089), .A1(n42939), .B0(n15196), .C0(n15197), .Y(
        n35238) );
  OA22XL U42383 ( .A0(net263919), .A1(n33073), .B0(n33081), .B1(n40043), .Y(
        n15196) );
  OAI211XL U42384 ( .A0(n33081), .A1(n42940), .B0(n15172), .C0(n15173), .Y(
        n35230) );
  OA22XL U42385 ( .A0(net218414), .A1(n33065), .B0(n33073), .B1(n40043), .Y(
        n15172) );
  OAI211XL U42386 ( .A0(n33073), .A1(n42941), .B0(n15148), .C0(n15149), .Y(
        n35222) );
  OA22XL U42387 ( .A0(net218456), .A1(n33057), .B0(n33065), .B1(net218670),
        .Y(n15148) );
  OAI211XL U42388 ( .A0(n33065), .A1(n42942), .B0(n15124), .C0(n15125), .Y(
        n35214) );
  OA22XL U42389 ( .A0(net218504), .A1(n33049), .B0(n33057), .B1(net218870),
        .Y(n15124) );
  OAI211XL U42390 ( .A0(n33057), .A1(n42944), .B0(n15100), .C0(n15101), .Y(
        n35206) );
  OA22XL U42391 ( .A0(net263957), .A1(n33041), .B0(n33049), .B1(n40042), .Y(
        n15100) );
  OAI211XL U42392 ( .A0(n33049), .A1(n42977), .B0(n15076), .C0(n15077), .Y(
        n35198) );
  OA22XL U42393 ( .A0(net263957), .A1(n33033), .B0(n33041), .B1(n40042), .Y(
        n15076) );
  OAI211XL U42394 ( .A0(n33041), .A1(n42978), .B0(n15052), .C0(n15053), .Y(
        n35190) );
  OA22XL U42395 ( .A0(net263976), .A1(n33025), .B0(n33033), .B1(n40041), .Y(
        n15052) );
  OAI211XL U42396 ( .A0(n33033), .A1(n42979), .B0(n15028), .C0(n15029), .Y(
        n35182) );
  OA22XL U42397 ( .A0(net263976), .A1(n33017), .B0(n33025), .B1(n40041), .Y(
        n15028) );
  OAI211XL U42398 ( .A0(n33025), .A1(n42980), .B0(n15004), .C0(n15005), .Y(
        n35174) );
  OA22XL U42399 ( .A0(net263995), .A1(n33009), .B0(n33017), .B1(n40040), .Y(
        n15004) );
  OAI211XL U42400 ( .A0(n33017), .A1(n42981), .B0(n14980), .C0(n14981), .Y(
        n35166) );
  OA22XL U42401 ( .A0(net263995), .A1(n33001), .B0(n33009), .B1(n40040), .Y(
        n14980) );
  OAI211XL U42402 ( .A0(n33009), .A1(n42983), .B0(n14956), .C0(n14957), .Y(
        n35158) );
  OA22XL U42403 ( .A0(net263805), .A1(n32993), .B0(n33001), .B1(n40050), .Y(
        n14956) );
  OAI211XL U42404 ( .A0(n33001), .A1(n42984), .B0(n14932), .C0(n14933), .Y(
        n35150) );
  OA22XL U42405 ( .A0(net263748), .A1(n32985), .B0(n32993), .B1(n40054), .Y(
        n14932) );
  OAI211XL U42406 ( .A0(n32993), .A1(n42985), .B0(n14908), .C0(n14909), .Y(
        n35142) );
  OA22XL U42407 ( .A0(net263748), .A1(n32977), .B0(n32985), .B1(n40053), .Y(
        n14908) );
  OAI211XL U42408 ( .A0(n32985), .A1(n42986), .B0(n14884), .C0(n14885), .Y(
        n35134) );
  OAI211XL U42409 ( .A0(n32977), .A1(n42987), .B0(n14860), .C0(n14861), .Y(
        n35126) );
  OAI211XL U42410 ( .A0(n32969), .A1(n42988), .B0(n14836), .C0(n14837), .Y(
        n35118) );
  OAI211XL U42411 ( .A0(n32961), .A1(n42989), .B0(n14812), .C0(n14813), .Y(
        n35110) );
  OA22XL U42412 ( .A0(net263292), .A1(n42725), .B0(n32401), .B1(n40079), .Y(
        n13156) );
  OA22XL U42413 ( .A0(net263292), .A1(n41380), .B0(n42725), .B1(n40078), .Y(
        n13132) );
  OAI211XL U42414 ( .A0(n34092), .A1(n42828), .B0(n18205), .C0(n18206), .Y(
        n36241) );
  OA22XL U42415 ( .A0(net262855), .A1(n34076), .B0(n34084), .B1(n40103), .Y(
        n18205) );
  OAI211XL U42416 ( .A0(n34084), .A1(n42829), .B0(n18181), .C0(n18182), .Y(
        n36233) );
  OA22XL U42417 ( .A0(net262874), .A1(n34068), .B0(n34076), .B1(n40103), .Y(
        n18181) );
  OAI211XL U42418 ( .A0(n34076), .A1(n42830), .B0(n18157), .C0(n18158), .Y(
        n36225) );
  OA22XL U42419 ( .A0(net262874), .A1(n34060), .B0(n34068), .B1(n40102), .Y(
        n18157) );
  OAI211XL U42420 ( .A0(n33988), .A1(n42810), .B0(n17893), .C0(n17894), .Y(
        n36137) );
  OA22XL U42421 ( .A0(net262703), .A1(n33972), .B0(n33980), .B1(n40110), .Y(
        n17893) );
  OAI211XL U42422 ( .A0(n33980), .A1(n42812), .B0(n17869), .C0(n17870), .Y(
        n36129) );
  OA22XL U42423 ( .A0(net262703), .A1(n33964), .B0(n33972), .B1(n40109), .Y(
        n17869) );
  OAI211XL U42424 ( .A0(n33972), .A1(n42813), .B0(n17845), .C0(n17846), .Y(
        n36121) );
  OA22XL U42425 ( .A0(net262722), .A1(n33956), .B0(n33964), .B1(n40109), .Y(
        n17845) );
  OAI211XL U42426 ( .A0(n33900), .A1(n42855), .B0(n17629), .C0(n17630), .Y(
        n36049) );
  OA22XL U42427 ( .A0(net261981), .A1(n33884), .B0(n33892), .B1(n40144), .Y(
        n17629) );
  OAI211XL U42428 ( .A0(n33892), .A1(n42856), .B0(n17605), .C0(n17606), .Y(
        n36041) );
  OA22XL U42429 ( .A0(net262000), .A1(n33876), .B0(n33884), .B1(n40144), .Y(
        n17605) );
  OAI211XL U42430 ( .A0(n33884), .A1(n42858), .B0(n17581), .C0(n17582), .Y(
        n36033) );
  OA22XL U42431 ( .A0(net262000), .A1(n33868), .B0(n33876), .B1(n40143), .Y(
        n17581) );
  OAI211XL U42432 ( .A0(n33876), .A1(n42859), .B0(n17557), .C0(n17558), .Y(
        n36025) );
  OA22XL U42433 ( .A0(net262000), .A1(n33860), .B0(n33868), .B1(n40143), .Y(
        n17557) );
  OAI211XL U42434 ( .A0(n33868), .A1(n42860), .B0(n17533), .C0(n17534), .Y(
        n36017) );
  OA22XL U42435 ( .A0(net262019), .A1(n33852), .B0(n33860), .B1(net218836),
        .Y(n17533) );
  OAI211XL U42436 ( .A0(n33860), .A1(n42861), .B0(n17509), .C0(n17510), .Y(
        n36009) );
  OA22XL U42437 ( .A0(net262019), .A1(n33844), .B0(n33852), .B1(n40053), .Y(
        n17509) );
  OAI211XL U42438 ( .A0(n33852), .A1(n42862), .B0(n17485), .C0(n17486), .Y(
        n36001) );
  OA22XL U42439 ( .A0(net262038), .A1(n33836), .B0(n33844), .B1(n40142), .Y(
        n17485) );
  OAI211XL U42440 ( .A0(n33844), .A1(n42831), .B0(n17461), .C0(n17462), .Y(
        n35993) );
  OA22XL U42441 ( .A0(net262038), .A1(n33828), .B0(n33836), .B1(n40142), .Y(
        n17461) );
  OAI211XL U42442 ( .A0(n33836), .A1(n42832), .B0(n17437), .C0(n17438), .Y(
        n35985) );
  OA22XL U42443 ( .A0(net262057), .A1(n33820), .B0(n33828), .B1(n40141), .Y(
        n17437) );
  OAI211XL U42444 ( .A0(n33828), .A1(n42833), .B0(n17413), .C0(n17414), .Y(
        n35977) );
  OA22XL U42445 ( .A0(net262057), .A1(n33812), .B0(n33820), .B1(n40141), .Y(
        n17413) );
  OAI211XL U42446 ( .A0(n33820), .A1(n42834), .B0(n17389), .C0(n17390), .Y(
        n35969) );
  OA22XL U42447 ( .A0(net263235), .A1(n33804), .B0(n33812), .B1(n40140), .Y(
        n17389) );
  OAI211XL U42448 ( .A0(n33812), .A1(n42836), .B0(n17365), .C0(n17366), .Y(
        n35961) );
  OA22XL U42449 ( .A0(net263463), .A1(n33796), .B0(n33804), .B1(n40140), .Y(
        n17365) );
  OAI211XL U42450 ( .A0(n33804), .A1(n42837), .B0(n17341), .C0(n17342), .Y(
        n35953) );
  OA22XL U42451 ( .A0(net218474), .A1(n33788), .B0(n33796), .B1(net218844),
        .Y(n17341) );
  OAI211XL U42452 ( .A0(n33772), .A1(n42841), .B0(n17245), .C0(n17246), .Y(
        n35921) );
  OA22XL U42453 ( .A0(net218294), .A1(n33756), .B0(n33764), .B1(net218610),
        .Y(n17245) );
  OAI211XL U42454 ( .A0(n33764), .A1(n42843), .B0(n17221), .C0(n17222), .Y(
        n35913) );
  OA22XL U42455 ( .A0(net218294), .A1(n33748), .B0(n33756), .B1(net218610),
        .Y(n17221) );
  OAI211XL U42456 ( .A0(n33756), .A1(n42844), .B0(n17197), .C0(n17198), .Y(
        n35905) );
  OA22XL U42457 ( .A0(net261867), .A1(n33740), .B0(n33748), .B1(n40151), .Y(
        n17197) );
  OAI211XL U42458 ( .A0(n33748), .A1(n42845), .B0(n17173), .C0(n17174), .Y(
        n35897) );
  OA22XL U42459 ( .A0(net261867), .A1(n33732), .B0(n33740), .B1(n40151), .Y(
        n17173) );
  OAI211XL U42460 ( .A0(n33740), .A1(n42846), .B0(n17149), .C0(n17150), .Y(
        n35889) );
  OA22XL U42461 ( .A0(net261886), .A1(n33724), .B0(n33732), .B1(n40150), .Y(
        n17149) );
  OAI211XL U42462 ( .A0(n34093), .A1(n42827), .B0(n18208), .C0(n18209), .Y(
        n36242) );
  OA22XL U42463 ( .A0(net262855), .A1(n34077), .B0(n34085), .B1(n40103), .Y(
        n18208) );
  OAI211XL U42464 ( .A0(n34085), .A1(n42829), .B0(n18184), .C0(n18185), .Y(
        n36234) );
  OA22XL U42465 ( .A0(net262874), .A1(n34069), .B0(n34077), .B1(n40103), .Y(
        n18184) );
  OAI211XL U42466 ( .A0(n34077), .A1(n42830), .B0(n18160), .C0(n18161), .Y(
        n36226) );
  OA22XL U42467 ( .A0(net262874), .A1(n34061), .B0(n34069), .B1(n40102), .Y(
        n18160) );
  OAI211XL U42468 ( .A0(n33989), .A1(n42810), .B0(n17896), .C0(n17897), .Y(
        n36138) );
  OA22XL U42469 ( .A0(net262703), .A1(n33973), .B0(n33981), .B1(n40110), .Y(
        n17896) );
  OAI211XL U42470 ( .A0(n33981), .A1(n42811), .B0(n17872), .C0(n17873), .Y(
        n36130) );
  OA22XL U42471 ( .A0(net262703), .A1(n33965), .B0(n33973), .B1(n40109), .Y(
        n17872) );
  OAI211XL U42472 ( .A0(n33973), .A1(n42813), .B0(n17848), .C0(n17849), .Y(
        n36122) );
  OA22XL U42473 ( .A0(net262722), .A1(n33957), .B0(n33965), .B1(n40109), .Y(
        n17848) );
  OAI211XL U42474 ( .A0(n33965), .A1(n42814), .B0(n17824), .C0(n17825), .Y(
        n36114) );
  OA22XL U42475 ( .A0(net262722), .A1(n33949), .B0(n33957), .B1(n40130), .Y(
        n17824) );
  OAI211XL U42476 ( .A0(n33957), .A1(n42847), .B0(n17800), .C0(n17801), .Y(
        n36106) );
  OA22XL U42477 ( .A0(net262741), .A1(n33941), .B0(n33949), .B1(n40058), .Y(
        n17800) );
  OAI211XL U42478 ( .A0(n33949), .A1(n42848), .B0(n17776), .C0(n17777), .Y(
        n36098) );
  OA22XL U42479 ( .A0(net262741), .A1(n33933), .B0(n33941), .B1(n40108), .Y(
        n17776) );
  OAI211XL U42480 ( .A0(n33941), .A1(n42849), .B0(n17752), .C0(n17753), .Y(
        n36090) );
  OA22XL U42481 ( .A0(net218504), .A1(n33925), .B0(n33933), .B1(n40108), .Y(
        n17752) );
  OAI211XL U42482 ( .A0(n33933), .A1(n42850), .B0(n17728), .C0(n17729), .Y(
        n36082) );
  OA22XL U42483 ( .A0(net218456), .A1(n33917), .B0(n33925), .B1(n40051), .Y(
        n17728) );
  OAI211XL U42484 ( .A0(n33925), .A1(n42852), .B0(n17704), .C0(n17705), .Y(
        n36074) );
  OA22XL U42485 ( .A0(net218452), .A1(n33909), .B0(n33917), .B1(net218632),
        .Y(n17704) );
  OAI211XL U42486 ( .A0(n33917), .A1(n42853), .B0(n17680), .C0(n17681), .Y(
        n36066) );
  OA22XL U42487 ( .A0(net262779), .A1(n33901), .B0(n33909), .B1(n40107), .Y(
        n17680) );
  OAI211XL U42488 ( .A0(n33909), .A1(n42854), .B0(n17656), .C0(n17657), .Y(
        n36058) );
  OA22XL U42489 ( .A0(net262779), .A1(n33893), .B0(n33901), .B1(n40107), .Y(
        n17656) );
  OAI211XL U42490 ( .A0(n33901), .A1(n42855), .B0(n17632), .C0(n17633), .Y(
        n36050) );
  OA22XL U42491 ( .A0(net261981), .A1(n33885), .B0(n33893), .B1(n40144), .Y(
        n17632) );
  OAI211XL U42492 ( .A0(n33893), .A1(n42856), .B0(n17608), .C0(n17609), .Y(
        n36042) );
  OA22XL U42493 ( .A0(net261981), .A1(n33877), .B0(n33885), .B1(n40144), .Y(
        n17608) );
  OAI211XL U42494 ( .A0(n33885), .A1(n42857), .B0(n17584), .C0(n17585), .Y(
        n36034) );
  OA22XL U42495 ( .A0(net262000), .A1(n33869), .B0(n33877), .B1(n40143), .Y(
        n17584) );
  OAI211XL U42496 ( .A0(n33877), .A1(n42859), .B0(n17560), .C0(n17561), .Y(
        n36026) );
  OA22XL U42497 ( .A0(net262000), .A1(n33861), .B0(n33869), .B1(n40143), .Y(
        n17560) );
  OAI211XL U42498 ( .A0(n33869), .A1(n42860), .B0(n17536), .C0(n17537), .Y(
        n36018) );
  OA22XL U42499 ( .A0(net262019), .A1(n33853), .B0(n33861), .B1(n40059), .Y(
        n17536) );
  OAI211XL U42500 ( .A0(n33861), .A1(n42861), .B0(n17512), .C0(n17513), .Y(
        n36010) );
  OA22XL U42501 ( .A0(net262019), .A1(n33845), .B0(n33853), .B1(n40046), .Y(
        n17512) );
  OAI211XL U42502 ( .A0(n33853), .A1(n42862), .B0(n17488), .C0(n17489), .Y(
        n36002) );
  OA22XL U42503 ( .A0(net262038), .A1(n33837), .B0(n33845), .B1(n40142), .Y(
        n17488) );
  OAI211XL U42504 ( .A0(n33845), .A1(n42831), .B0(n17464), .C0(n17465), .Y(
        n35994) );
  OA22XL U42505 ( .A0(net262038), .A1(n33829), .B0(n33837), .B1(n40142), .Y(
        n17464) );
  OAI211XL U42506 ( .A0(n33837), .A1(n42832), .B0(n17440), .C0(n17441), .Y(
        n35986) );
  OA22XL U42507 ( .A0(net262057), .A1(n33821), .B0(n33829), .B1(n40141), .Y(
        n17440) );
  OAI211XL U42508 ( .A0(n33829), .A1(n42833), .B0(n17416), .C0(n17417), .Y(
        n35978) );
  OA22XL U42509 ( .A0(net262057), .A1(n33813), .B0(n33821), .B1(n40141), .Y(
        n17416) );
  OAI211XL U42510 ( .A0(n33821), .A1(n42834), .B0(n17392), .C0(n17393), .Y(
        n35970) );
  OA22XL U42511 ( .A0(net263292), .A1(n33805), .B0(n33813), .B1(n40140), .Y(
        n17392) );
  OAI211XL U42512 ( .A0(n33813), .A1(n42835), .B0(n17368), .C0(n17369), .Y(
        n35962) );
  OA22XL U42513 ( .A0(net263235), .A1(n33797), .B0(n33805), .B1(n40140), .Y(
        n17368) );
  OAI211XL U42514 ( .A0(n33805), .A1(n42837), .B0(n17344), .C0(n17345), .Y(
        n35954) );
  OA22XL U42515 ( .A0(net263235), .A1(n33789), .B0(n33797), .B1(n40087), .Y(
        n17344) );
  OAI211XL U42516 ( .A0(n33797), .A1(n42838), .B0(n17320), .C0(n17321), .Y(
        n35946) );
  OA22XL U42517 ( .A0(net262095), .A1(n33781), .B0(n33789), .B1(n40087), .Y(
        n17320) );
  OAI211XL U42518 ( .A0(n33789), .A1(n42839), .B0(n17296), .C0(n17297), .Y(
        n35938) );
  OA22XL U42519 ( .A0(net262095), .A1(n33773), .B0(n33781), .B1(n40139), .Y(
        n17296) );
  OAI211XL U42520 ( .A0(n33781), .A1(n42840), .B0(n17272), .C0(n17273), .Y(
        n35930) );
  OA22XL U42521 ( .A0(net262114), .A1(n33765), .B0(n33773), .B1(n40139), .Y(
        n17272) );
  OAI211XL U42522 ( .A0(n33773), .A1(n42841), .B0(n17248), .C0(n17249), .Y(
        n35922) );
  OA22XL U42523 ( .A0(net218294), .A1(n33757), .B0(n33765), .B1(net218610),
        .Y(n17248) );
  OAI211XL U42524 ( .A0(n33765), .A1(n42842), .B0(n17224), .C0(n17225), .Y(
        n35914) );
  OA22XL U42525 ( .A0(net218294), .A1(n33749), .B0(n33757), .B1(net218610),
        .Y(n17224) );
  OAI211XL U42526 ( .A0(n33757), .A1(n42844), .B0(n17200), .C0(n17201), .Y(
        n35906) );
  OA22XL U42527 ( .A0(net261867), .A1(n33741), .B0(n33749), .B1(n40151), .Y(
        n17200) );
  OAI211XL U42528 ( .A0(n33749), .A1(n42845), .B0(n17176), .C0(n17177), .Y(
        n35898) );
  OA22XL U42529 ( .A0(net261867), .A1(n33733), .B0(n33741), .B1(n40151), .Y(
        n17176) );
  OAI211XL U42530 ( .A0(n33741), .A1(n42846), .B0(n17152), .C0(n17153), .Y(
        n35890) );
  OA22XL U42531 ( .A0(net261886), .A1(n33725), .B0(n33733), .B1(n40150), .Y(
        n17152) );
  OAI211XL U42532 ( .A0(n34094), .A1(n42827), .B0(n18211), .C0(n18212), .Y(
        n36243) );
  OA22XL U42533 ( .A0(net262855), .A1(n34078), .B0(n34086), .B1(n40103), .Y(
        n18211) );
  OAI211XL U42534 ( .A0(n34086), .A1(n42828), .B0(n18187), .C0(n18188), .Y(
        n36235) );
  OA22XL U42535 ( .A0(net262874), .A1(n34070), .B0(n34078), .B1(n40103), .Y(
        n18187) );
  OAI211XL U42536 ( .A0(n34078), .A1(n42830), .B0(n18163), .C0(n18164), .Y(
        n36227) );
  OA22XL U42537 ( .A0(net262874), .A1(n34062), .B0(n34070), .B1(n40102), .Y(
        n18163) );
  OAI211XL U42538 ( .A0(n33990), .A1(n42810), .B0(n17899), .C0(n17900), .Y(
        n36139) );
  OA22XL U42539 ( .A0(net262703), .A1(n33974), .B0(n33982), .B1(n40110), .Y(
        n17899) );
  OAI211XL U42540 ( .A0(n33982), .A1(n42811), .B0(n17875), .C0(n17876), .Y(
        n36131) );
  OA22XL U42541 ( .A0(net262703), .A1(n33966), .B0(n33974), .B1(n40109), .Y(
        n17875) );
  OAI211XL U42542 ( .A0(n33974), .A1(n42812), .B0(n17851), .C0(n17852), .Y(
        n36123) );
  OA22XL U42543 ( .A0(net262722), .A1(n33958), .B0(n33966), .B1(n40109), .Y(
        n17851) );
  OAI211XL U42544 ( .A0(n33966), .A1(n42814), .B0(n17827), .C0(n17828), .Y(
        n36115) );
  OA22XL U42545 ( .A0(net262722), .A1(n33950), .B0(n33958), .B1(n40130), .Y(
        n17827) );
  OAI211XL U42546 ( .A0(n33958), .A1(n42855), .B0(n17803), .C0(n17804), .Y(
        n36107) );
  OA22XL U42547 ( .A0(net262741), .A1(n33942), .B0(n33950), .B1(n40130), .Y(
        n17803) );
  OAI211XL U42548 ( .A0(n33950), .A1(n42848), .B0(n17779), .C0(n17780), .Y(
        n36099) );
  OA22XL U42549 ( .A0(net262741), .A1(n33934), .B0(n33942), .B1(n40108), .Y(
        n17779) );
  OAI211XL U42550 ( .A0(n33942), .A1(n42849), .B0(n17755), .C0(n17756), .Y(
        n36091) );
  OA22XL U42551 ( .A0(net218504), .A1(n33926), .B0(n33934), .B1(n40108), .Y(
        n17755) );
  OAI211XL U42552 ( .A0(n33934), .A1(n42850), .B0(n17731), .C0(n17732), .Y(
        n36083) );
  OA22XL U42553 ( .A0(net218506), .A1(n33918), .B0(n33926), .B1(n40068), .Y(
        n17731) );
  OAI211XL U42554 ( .A0(n33926), .A1(n42851), .B0(n17707), .C0(n17708), .Y(
        n36075) );
  OA22XL U42555 ( .A0(net218312), .A1(n33910), .B0(n33918), .B1(n40068), .Y(
        n17707) );
  OAI211XL U42556 ( .A0(n33918), .A1(n42853), .B0(n17683), .C0(n17684), .Y(
        n36067) );
  OA22XL U42557 ( .A0(net262779), .A1(n33902), .B0(n33910), .B1(n40107), .Y(
        n17683) );
  OAI211XL U42558 ( .A0(n33910), .A1(n42854), .B0(n17659), .C0(n17660), .Y(
        n36059) );
  OA22XL U42559 ( .A0(net262779), .A1(n33894), .B0(n33902), .B1(n40107), .Y(
        n17659) );
  OAI211XL U42560 ( .A0(n33902), .A1(n42855), .B0(n17635), .C0(n17636), .Y(
        n36051) );
  OA22XL U42561 ( .A0(net261981), .A1(n33886), .B0(n33894), .B1(n40144), .Y(
        n17635) );
  OAI211XL U42562 ( .A0(n33894), .A1(n42856), .B0(n17611), .C0(n17612), .Y(
        n36043) );
  OA22XL U42563 ( .A0(net261981), .A1(n33878), .B0(n33886), .B1(n40144), .Y(
        n17611) );
  OAI211XL U42564 ( .A0(n33886), .A1(n42857), .B0(n17587), .C0(n17588), .Y(
        n36035) );
  OA22XL U42565 ( .A0(net262000), .A1(n33870), .B0(n33878), .B1(n40143), .Y(
        n17587) );
  OAI211XL U42566 ( .A0(n33878), .A1(n42858), .B0(n17563), .C0(n17564), .Y(
        n36027) );
  OA22XL U42567 ( .A0(net262000), .A1(n33862), .B0(n33870), .B1(n40143), .Y(
        n17563) );
  OAI211XL U42568 ( .A0(n33870), .A1(n42860), .B0(n17539), .C0(n17540), .Y(
        n36019) );
  OA22XL U42569 ( .A0(net262019), .A1(n33854), .B0(n33862), .B1(n40060), .Y(
        n17539) );
  OAI211XL U42570 ( .A0(n33862), .A1(n42861), .B0(n17515), .C0(n17516), .Y(
        n36011) );
  OA22XL U42571 ( .A0(net262019), .A1(n33846), .B0(n33854), .B1(n40040), .Y(
        n17515) );
  OAI211XL U42572 ( .A0(n33854), .A1(n42862), .B0(n17491), .C0(n17492), .Y(
        n36003) );
  OA22XL U42573 ( .A0(net262038), .A1(n33838), .B0(n33846), .B1(n40142), .Y(
        n17491) );
  OAI211XL U42574 ( .A0(n33846), .A1(n42839), .B0(n17467), .C0(n17468), .Y(
        n35995) );
  OA22XL U42575 ( .A0(net262038), .A1(n33830), .B0(n33838), .B1(n40142), .Y(
        n17467) );
  OAI211XL U42576 ( .A0(n33838), .A1(n42832), .B0(n17443), .C0(n17444), .Y(
        n35987) );
  OA22XL U42577 ( .A0(net262057), .A1(n33822), .B0(n33830), .B1(n40141), .Y(
        n17443) );
  OAI211XL U42578 ( .A0(n33830), .A1(n42833), .B0(n17419), .C0(n17420), .Y(
        n35979) );
  OA22XL U42579 ( .A0(net262057), .A1(n33814), .B0(n33822), .B1(n40141), .Y(
        n17419) );
  OAI211XL U42580 ( .A0(n33822), .A1(n42834), .B0(n17395), .C0(n17396), .Y(
        n35971) );
  OA22XL U42581 ( .A0(net262057), .A1(n33806), .B0(n33814), .B1(n40140), .Y(
        n17395) );
  OAI211XL U42582 ( .A0(n33814), .A1(n42835), .B0(n17371), .C0(n17372), .Y(
        n35963) );
  OA22XL U42583 ( .A0(net263216), .A1(n33798), .B0(n33806), .B1(n40140), .Y(
        n17371) );
  OAI211XL U42584 ( .A0(n33806), .A1(n42836), .B0(n17347), .C0(n17348), .Y(
        n35955) );
  OA22XL U42585 ( .A0(net263292), .A1(n33790), .B0(n33798), .B1(n40088), .Y(
        n17347) );
  OAI211XL U42586 ( .A0(n33798), .A1(n42838), .B0(n17323), .C0(n17324), .Y(
        n35947) );
  OA22XL U42587 ( .A0(net262095), .A1(n33782), .B0(n33790), .B1(n40042), .Y(
        n17323) );
  OAI211XL U42588 ( .A0(n33790), .A1(n42839), .B0(n17299), .C0(n17300), .Y(
        n35939) );
  OA22XL U42589 ( .A0(net262095), .A1(n33774), .B0(n33782), .B1(n40139), .Y(
        n17299) );
  OAI211XL U42590 ( .A0(n33782), .A1(n42840), .B0(n17275), .C0(n17276), .Y(
        n35931) );
  OA22XL U42591 ( .A0(net262114), .A1(n33766), .B0(n33774), .B1(n40139), .Y(
        n17275) );
  OAI211XL U42592 ( .A0(n33774), .A1(n42841), .B0(n17251), .C0(n17252), .Y(
        n35923) );
  OA22XL U42593 ( .A0(net218294), .A1(n33758), .B0(n33766), .B1(net218610),
        .Y(n17251) );
  OAI211XL U42594 ( .A0(n33766), .A1(n42842), .B0(n17227), .C0(n17228), .Y(
        n35915) );
  OA22XL U42595 ( .A0(net218294), .A1(n33750), .B0(n33758), .B1(net218610),
        .Y(n17227) );
  OAI211XL U42596 ( .A0(n33758), .A1(n42843), .B0(n17203), .C0(n17204), .Y(
        n35907) );
  OA22XL U42597 ( .A0(net261867), .A1(n33742), .B0(n33750), .B1(n40151), .Y(
        n17203) );
  OAI211XL U42598 ( .A0(n33750), .A1(n42845), .B0(n17179), .C0(n17180), .Y(
        n35899) );
  OA22XL U42599 ( .A0(net261867), .A1(n33734), .B0(n33742), .B1(n40151), .Y(
        n17179) );
  OAI211XL U42600 ( .A0(n33742), .A1(n42846), .B0(n17155), .C0(n17156), .Y(
        n35891) );
  OA22XL U42601 ( .A0(net261886), .A1(n33726), .B0(n33734), .B1(n40150), .Y(
        n17155) );
  OAI211XL U42602 ( .A0(n33734), .A1(n42847), .B0(n17131), .C0(n17132), .Y(
        n35883) );
  OA22XL U42603 ( .A0(net261886), .A1(n33718), .B0(n33726), .B1(n40150), .Y(
        n17131) );
  OAI211XL U42604 ( .A0(n34096), .A1(n42827), .B0(n18217), .C0(n18218), .Y(
        n36245) );
  OA22XL U42605 ( .A0(net262855), .A1(n34080), .B0(n34088), .B1(n40103), .Y(
        n18217) );
  OAI211XL U42606 ( .A0(n34088), .A1(n42828), .B0(n18193), .C0(n18194), .Y(
        n36237) );
  OA22XL U42607 ( .A0(net262874), .A1(n34072), .B0(n34080), .B1(n40103), .Y(
        n18193) );
  OAI211XL U42608 ( .A0(n34080), .A1(n42829), .B0(n18169), .C0(n18170), .Y(
        n36229) );
  OA22XL U42609 ( .A0(net262874), .A1(n34064), .B0(n34072), .B1(n40102), .Y(
        n18169) );
  OAI211XL U42610 ( .A0(n34072), .A1(n42830), .B0(n18145), .C0(n18146), .Y(
        n36221) );
  OA22XL U42611 ( .A0(net262874), .A1(n34056), .B0(n34064), .B1(n40102), .Y(
        n18145) );
  OAI211XL U42612 ( .A0(n33992), .A1(n42810), .B0(n17905), .C0(n17906), .Y(
        n36141) );
  OA22XL U42613 ( .A0(net262703), .A1(n33976), .B0(n33984), .B1(n40110), .Y(
        n17905) );
  OAI211XL U42614 ( .A0(n33984), .A1(n42811), .B0(n17881), .C0(n17882), .Y(
        n36133) );
  OA22XL U42615 ( .A0(net262703), .A1(n33968), .B0(n33976), .B1(n40109), .Y(
        n17881) );
  OAI211XL U42616 ( .A0(n33976), .A1(n42812), .B0(n17857), .C0(n17858), .Y(
        n36125) );
  OA22XL U42617 ( .A0(net262722), .A1(n33960), .B0(n33968), .B1(n40109), .Y(
        n17857) );
  OAI211XL U42618 ( .A0(n33968), .A1(n42813), .B0(n17833), .C0(n17834), .Y(
        n36117) );
  OA22XL U42619 ( .A0(net262722), .A1(n33952), .B0(n33960), .B1(n40094), .Y(
        n17833) );
  OAI211XL U42620 ( .A0(n33960), .A1(n42814), .B0(n17809), .C0(n17810), .Y(
        n36109) );
  OA22XL U42621 ( .A0(net262741), .A1(n33944), .B0(n33952), .B1(n40051), .Y(
        n17809) );
  OAI211XL U42622 ( .A0(n33952), .A1(n42848), .B0(n17785), .C0(n17786), .Y(
        n36101) );
  OA22XL U42623 ( .A0(net262741), .A1(n33936), .B0(n33944), .B1(n40108), .Y(
        n17785) );
  OAI211XL U42624 ( .A0(n33944), .A1(n42849), .B0(n17761), .C0(n17762), .Y(
        n36093) );
  OA22XL U42625 ( .A0(net262741), .A1(n33928), .B0(n33936), .B1(n40108), .Y(
        n17761) );
  OAI211XL U42626 ( .A0(n33936), .A1(n42850), .B0(n17737), .C0(n17738), .Y(
        n36085) );
  OA22XL U42627 ( .A0(net218442), .A1(n33920), .B0(n33928), .B1(n40052), .Y(
        n17737) );
  OAI211XL U42628 ( .A0(n33928), .A1(n42851), .B0(n17713), .C0(n17714), .Y(
        n36077) );
  OA22XL U42629 ( .A0(net218452), .A1(n33912), .B0(n33920), .B1(n40057), .Y(
        n17713) );
  OAI211XL U42630 ( .A0(n33920), .A1(n42852), .B0(n17689), .C0(n17690), .Y(
        n36069) );
  OA22XL U42631 ( .A0(net262779), .A1(n33904), .B0(n33912), .B1(n40107), .Y(
        n17689) );
  OAI211XL U42632 ( .A0(n33912), .A1(n42853), .B0(n17665), .C0(n17666), .Y(
        n36061) );
  OA22XL U42633 ( .A0(net262779), .A1(n33896), .B0(n33904), .B1(n40107), .Y(
        n17665) );
  OAI211XL U42634 ( .A0(n33904), .A1(n42855), .B0(n17641), .C0(n17642), .Y(
        n36053) );
  OA22XL U42635 ( .A0(net262114), .A1(n33888), .B0(n33896), .B1(n40138), .Y(
        n17641) );
  OAI211XL U42636 ( .A0(n33896), .A1(n42856), .B0(n17617), .C0(n17618), .Y(
        n36045) );
  OA22XL U42637 ( .A0(net261981), .A1(n33880), .B0(n33888), .B1(n40144), .Y(
        n17617) );
  OAI211XL U42638 ( .A0(n33888), .A1(n42857), .B0(n17593), .C0(n17594), .Y(
        n36037) );
  OA22XL U42639 ( .A0(net262000), .A1(n33872), .B0(n33880), .B1(n40143), .Y(
        n17593) );
  OAI211XL U42640 ( .A0(n33880), .A1(n42858), .B0(n17569), .C0(n17570), .Y(
        n36029) );
  OA22XL U42641 ( .A0(net262000), .A1(n33864), .B0(n33872), .B1(n40143), .Y(
        n17569) );
  OAI211XL U42642 ( .A0(n33872), .A1(n42859), .B0(n17545), .C0(n17546), .Y(
        n36021) );
  OA22XL U42643 ( .A0(net262019), .A1(n33856), .B0(n33864), .B1(n40041), .Y(
        n17545) );
  OAI211XL U42644 ( .A0(n33864), .A1(n42860), .B0(n17521), .C0(n17522), .Y(
        n36013) );
  OA22XL U42645 ( .A0(net262019), .A1(n33848), .B0(n33856), .B1(n40058), .Y(
        n17521) );
  OAI211XL U42646 ( .A0(n33856), .A1(n42862), .B0(n17497), .C0(n17498), .Y(
        n36005) );
  OA22XL U42647 ( .A0(net262038), .A1(n33840), .B0(n33848), .B1(n40142), .Y(
        n17497) );
  OAI211XL U42648 ( .A0(n33848), .A1(n42863), .B0(n17473), .C0(n17474), .Y(
        n35997) );
  OA22XL U42649 ( .A0(net262038), .A1(n33832), .B0(n33840), .B1(n40142), .Y(
        n17473) );
  OAI211XL U42650 ( .A0(n33840), .A1(n42832), .B0(n17449), .C0(n17450), .Y(
        n35989) );
  OA22XL U42651 ( .A0(net262038), .A1(n33824), .B0(n33832), .B1(n40141), .Y(
        n17449) );
  OAI211XL U42652 ( .A0(n33832), .A1(n42833), .B0(n17425), .C0(n17426), .Y(
        n35981) );
  OA22XL U42653 ( .A0(net262057), .A1(n33816), .B0(n33824), .B1(n40141), .Y(
        n17425) );
  OAI211XL U42654 ( .A0(n33824), .A1(n42834), .B0(n17401), .C0(n17402), .Y(
        n35973) );
  OA22XL U42655 ( .A0(net262057), .A1(n33808), .B0(n33816), .B1(n40140), .Y(
        n17401) );
  OAI211XL U42656 ( .A0(n33816), .A1(n42835), .B0(n17377), .C0(n17378), .Y(
        n35965) );
  OA22XL U42657 ( .A0(net263292), .A1(n33800), .B0(n33808), .B1(n40140), .Y(
        n17377) );
  OAI211XL U42658 ( .A0(n33808), .A1(n42836), .B0(n17353), .C0(n17354), .Y(
        n35957) );
  OA22XL U42659 ( .A0(net263292), .A1(n33792), .B0(n33800), .B1(n40047), .Y(
        n17353) );
  OAI211XL U42660 ( .A0(n33800), .A1(n42837), .B0(n17329), .C0(n17330), .Y(
        n35949) );
  OA22XL U42661 ( .A0(net262095), .A1(n33784), .B0(n33792), .B1(n40049), .Y(
        n17329) );
  OAI211XL U42662 ( .A0(n33792), .A1(n42838), .B0(n17305), .C0(n17306), .Y(
        n35941) );
  OA22XL U42663 ( .A0(net262095), .A1(n33776), .B0(n33784), .B1(n40139), .Y(
        n17305) );
  OAI211XL U42664 ( .A0(n33784), .A1(n42840), .B0(n17281), .C0(n17282), .Y(
        n35933) );
  OA22XL U42665 ( .A0(net262114), .A1(n33768), .B0(n33776), .B1(n40139), .Y(
        n17281) );
  OAI211XL U42666 ( .A0(n33776), .A1(n42841), .B0(n17257), .C0(n17258), .Y(
        n35925) );
  OA22XL U42667 ( .A0(net261905), .A1(n33760), .B0(n33768), .B1(n40148), .Y(
        n17257) );
  OAI211XL U42668 ( .A0(n33768), .A1(n42842), .B0(n17233), .C0(n17234), .Y(
        n35917) );
  OA22XL U42669 ( .A0(net218294), .A1(n33752), .B0(n33760), .B1(net218610),
        .Y(n17233) );
  OAI211XL U42670 ( .A0(n33760), .A1(n42843), .B0(n17209), .C0(n17210), .Y(
        n35909) );
  OA22XL U42671 ( .A0(net261867), .A1(n33744), .B0(n33752), .B1(n40151), .Y(
        n17209) );
  OAI211XL U42672 ( .A0(n33752), .A1(n42844), .B0(n17185), .C0(n17186), .Y(
        n35901) );
  OA22XL U42673 ( .A0(net261867), .A1(n33736), .B0(n33744), .B1(n40151), .Y(
        n17185) );
  OAI211XL U42674 ( .A0(n33744), .A1(n42845), .B0(n17161), .C0(n17162), .Y(
        n35893) );
  OA22XL U42675 ( .A0(net261886), .A1(n33728), .B0(n33736), .B1(n40150), .Y(
        n17161) );
  OAI211XL U42676 ( .A0(n33736), .A1(n42847), .B0(n17137), .C0(n17138), .Y(
        n35885) );
  OA22XL U42677 ( .A0(net261886), .A1(n33720), .B0(n33728), .B1(n40150), .Y(
        n17137) );
  OAI211XL U42678 ( .A0(n34081), .A1(n42829), .B0(n18172), .C0(n18173), .Y(
        n36230) );
  OA22XL U42679 ( .A0(net262874), .A1(n34065), .B0(n34073), .B1(n40102), .Y(
        n18172) );
  OAI211XL U42680 ( .A0(n34073), .A1(n42830), .B0(n18148), .C0(n18149), .Y(
        n36222) );
  OA22XL U42681 ( .A0(net262874), .A1(n34057), .B0(n34065), .B1(n40102), .Y(
        n18148) );
  OAI211XL U42682 ( .A0(n33993), .A1(n42810), .B0(n17908), .C0(n17909), .Y(
        n36142) );
  OA22XL U42683 ( .A0(net262703), .A1(n33977), .B0(n33985), .B1(n40110), .Y(
        n17908) );
  OAI211XL U42684 ( .A0(n33985), .A1(n42811), .B0(n17884), .C0(n17885), .Y(
        n36134) );
  OA22XL U42685 ( .A0(net262703), .A1(n33969), .B0(n33977), .B1(n40109), .Y(
        n17884) );
  OAI211XL U42686 ( .A0(n33977), .A1(n42812), .B0(n17860), .C0(n17861), .Y(
        n36126) );
  OA22XL U42687 ( .A0(net262722), .A1(n33961), .B0(n33969), .B1(n40109), .Y(
        n17860) );
  OAI211XL U42688 ( .A0(n33969), .A1(n42813), .B0(n17836), .C0(n17837), .Y(
        n36118) );
  OA22XL U42689 ( .A0(net262722), .A1(n33953), .B0(n33961), .B1(net218866),
        .Y(n17836) );
  OAI211XL U42690 ( .A0(n33961), .A1(n42814), .B0(n17812), .C0(n17813), .Y(
        n36110) );
  OA22XL U42691 ( .A0(net262722), .A1(n33945), .B0(n33953), .B1(n40052), .Y(
        n17812) );
  OAI211XL U42692 ( .A0(n33953), .A1(n42848), .B0(n17788), .C0(n17789), .Y(
        n36102) );
  OA22XL U42693 ( .A0(net262741), .A1(n33937), .B0(n33945), .B1(n40108), .Y(
        n17788) );
  OAI211XL U42694 ( .A0(n33945), .A1(n42849), .B0(n17764), .C0(n17765), .Y(
        n36094) );
  OA22XL U42695 ( .A0(net262741), .A1(n33929), .B0(n33937), .B1(n40108), .Y(
        n17764) );
  OAI211XL U42696 ( .A0(n33937), .A1(n42850), .B0(n17740), .C0(n17741), .Y(
        n36086) );
  OA22XL U42697 ( .A0(net218462), .A1(n33921), .B0(n33929), .B1(n40068), .Y(
        n17740) );
  OAI211XL U42698 ( .A0(n33929), .A1(n42851), .B0(n17716), .C0(n17717), .Y(
        n36078) );
  OA22XL U42699 ( .A0(net218462), .A1(n33913), .B0(n33921), .B1(n40068), .Y(
        n17716) );
  OAI211XL U42700 ( .A0(n33921), .A1(n42852), .B0(n17692), .C0(n17693), .Y(
        n36070) );
  OA22XL U42701 ( .A0(net262779), .A1(n33905), .B0(n33913), .B1(n40107), .Y(
        n17692) );
  OAI211XL U42702 ( .A0(n33913), .A1(n42853), .B0(n17668), .C0(n17669), .Y(
        n36062) );
  OA22XL U42703 ( .A0(net262779), .A1(n33897), .B0(n33905), .B1(n40107), .Y(
        n17668) );
  OAI211XL U42704 ( .A0(n33905), .A1(n42854), .B0(n17644), .C0(n17645), .Y(
        n36054) );
  OA22XL U42705 ( .A0(net262798), .A1(n33889), .B0(n33897), .B1(n40106), .Y(
        n17644) );
  OAI211XL U42706 ( .A0(n33897), .A1(n42856), .B0(n17620), .C0(n17621), .Y(
        n36046) );
  OA22XL U42707 ( .A0(net261981), .A1(n33881), .B0(n33889), .B1(n40144), .Y(
        n17620) );
  OAI211XL U42708 ( .A0(n33889), .A1(n42857), .B0(n17596), .C0(n17597), .Y(
        n36038) );
  OA22XL U42709 ( .A0(net262000), .A1(n33873), .B0(n33881), .B1(n40143), .Y(
        n17596) );
  OAI211XL U42710 ( .A0(n33881), .A1(n42858), .B0(n17572), .C0(n17573), .Y(
        n36030) );
  OA22XL U42711 ( .A0(net262000), .A1(n33865), .B0(n33873), .B1(n40143), .Y(
        n17572) );
  OAI211XL U42712 ( .A0(n33873), .A1(n42859), .B0(n17548), .C0(n17549), .Y(
        n36022) );
  OA22XL U42713 ( .A0(net262019), .A1(n33857), .B0(n33865), .B1(net218864),
        .Y(n17548) );
  OAI211XL U42714 ( .A0(n33865), .A1(n42860), .B0(n17524), .C0(n17525), .Y(
        n36014) );
  OA22XL U42715 ( .A0(net262019), .A1(n33849), .B0(n33857), .B1(net218860),
        .Y(n17524) );
  OAI211XL U42716 ( .A0(n33857), .A1(n42861), .B0(n17500), .C0(n17501), .Y(
        n36006) );
  OA22XL U42717 ( .A0(net262019), .A1(n33841), .B0(n33849), .B1(n40142), .Y(
        n17500) );
  OAI211XL U42718 ( .A0(n33849), .A1(n42863), .B0(n17476), .C0(n17477), .Y(
        n35998) );
  OA22XL U42719 ( .A0(net262038), .A1(n33833), .B0(n33841), .B1(n40142), .Y(
        n17476) );
  OAI211XL U42720 ( .A0(n33841), .A1(n42831), .B0(n17452), .C0(n17453), .Y(
        n35990) );
  OA22XL U42721 ( .A0(net262038), .A1(n33825), .B0(n33833), .B1(n40141), .Y(
        n17452) );
  OAI211XL U42722 ( .A0(n33833), .A1(n42833), .B0(n17428), .C0(n17429), .Y(
        n35982) );
  OA22XL U42723 ( .A0(net262057), .A1(n33817), .B0(n33825), .B1(n40141), .Y(
        n17428) );
  OAI211XL U42724 ( .A0(n33825), .A1(n42834), .B0(n17404), .C0(n17405), .Y(
        n35974) );
  OA22XL U42725 ( .A0(net262057), .A1(n33809), .B0(n33817), .B1(n40140), .Y(
        n17404) );
  OAI211XL U42726 ( .A0(n33817), .A1(n42835), .B0(n17380), .C0(n17381), .Y(
        n35966) );
  OA22XL U42727 ( .A0(net218302), .A1(n33801), .B0(n33809), .B1(n40140), .Y(
        n17380) );
  OAI211XL U42728 ( .A0(n33809), .A1(n42836), .B0(n17356), .C0(n17357), .Y(
        n35958) );
  OA22XL U42729 ( .A0(net218298), .A1(n33793), .B0(n33801), .B1(net218852),
        .Y(n17356) );
  OAI211XL U42730 ( .A0(n33801), .A1(n42837), .B0(n17332), .C0(n17333), .Y(
        n35950) );
  OA22XL U42731 ( .A0(net262095), .A1(n33785), .B0(n33793), .B1(net218854),
        .Y(n17332) );
  OAI211XL U42732 ( .A0(n33793), .A1(n42838), .B0(n17308), .C0(n17309), .Y(
        n35942) );
  OA22XL U42733 ( .A0(net262095), .A1(n33777), .B0(n33785), .B1(n40139), .Y(
        n17308) );
  OAI211XL U42734 ( .A0(n33785), .A1(n42840), .B0(n17284), .C0(n17285), .Y(
        n35934) );
  OA22XL U42735 ( .A0(net262114), .A1(n33769), .B0(n33777), .B1(n40139), .Y(
        n17284) );
  OAI211XL U42736 ( .A0(n33777), .A1(n42841), .B0(n17260), .C0(n17261), .Y(
        n35926) );
  OA22XL U42737 ( .A0(net262114), .A1(n33761), .B0(n33769), .B1(n40138), .Y(
        n17260) );
  OAI211XL U42738 ( .A0(n33769), .A1(n42842), .B0(n17236), .C0(n17237), .Y(
        n35918) );
  OA22XL U42739 ( .A0(net218294), .A1(n33753), .B0(n33761), .B1(net218610),
        .Y(n17236) );
  OAI211XL U42740 ( .A0(n33761), .A1(n42843), .B0(n17212), .C0(n17213), .Y(
        n35910) );
  OA22XL U42741 ( .A0(net261867), .A1(n33745), .B0(n33753), .B1(n40151), .Y(
        n17212) );
  OAI211XL U42742 ( .A0(n33753), .A1(n42844), .B0(n17188), .C0(n17189), .Y(
        n35902) );
  OA22XL U42743 ( .A0(net261867), .A1(n33737), .B0(n33745), .B1(n40151), .Y(
        n17188) );
  OAI211XL U42744 ( .A0(n33745), .A1(n42845), .B0(n17164), .C0(n17165), .Y(
        n35894) );
  OA22XL U42745 ( .A0(net261886), .A1(n33729), .B0(n33737), .B1(n40150), .Y(
        n17164) );
  OAI211XL U42746 ( .A0(n33737), .A1(n42846), .B0(n17140), .C0(n17141), .Y(
        n35886) );
  OA22XL U42747 ( .A0(net261886), .A1(n33721), .B0(n33729), .B1(n40150), .Y(
        n17140) );
  OAI211XL U42748 ( .A0(n33612), .A1(n42736), .B0(n16765), .C0(n16766), .Y(
        n35761) );
  OA22XL U42749 ( .A0(net262285), .A1(n33596), .B0(n33604), .B1(n40090), .Y(
        n16765) );
  OAI211XL U42750 ( .A0(n33596), .A1(n42738), .B0(n16717), .C0(n16718), .Y(
        n35745) );
  OA22XL U42751 ( .A0(net262304), .A1(n33580), .B0(n33588), .B1(n40128), .Y(
        n16717) );
  OAI211XL U42752 ( .A0(n33588), .A1(n42739), .B0(n16693), .C0(n16694), .Y(
        n35737) );
  OA22XL U42753 ( .A0(net262304), .A1(n33572), .B0(n33580), .B1(n40128), .Y(
        n16693) );
  OAI211XL U42754 ( .A0(n33613), .A1(n42736), .B0(n16768), .C0(n16769), .Y(
        n35762) );
  OA22XL U42755 ( .A0(net262285), .A1(n33597), .B0(n33605), .B1(net218780),
        .Y(n16768) );
  OAI211XL U42756 ( .A0(n33589), .A1(n42739), .B0(n16696), .C0(n16697), .Y(
        n35738) );
  OA22XL U42757 ( .A0(net262304), .A1(n33573), .B0(n33581), .B1(n40128), .Y(
        n16696) );
  OAI211XL U42758 ( .A0(n33614), .A1(n42736), .B0(n16771), .C0(n16772), .Y(
        n35763) );
  OA22XL U42759 ( .A0(net262285), .A1(n33598), .B0(n33606), .B1(net218786),
        .Y(n16771) );
  OAI211XL U42760 ( .A0(n33590), .A1(n42738), .B0(n16699), .C0(n16700), .Y(
        n35739) );
  OA22XL U42761 ( .A0(net262304), .A1(n33574), .B0(n33582), .B1(n40128), .Y(
        n16699) );
  OAI211XL U42762 ( .A0(n33616), .A1(n42736), .B0(n16777), .C0(n16778), .Y(
        n35765) );
  OA22XL U42763 ( .A0(net262285), .A1(n33600), .B0(n33608), .B1(net218760),
        .Y(n16777) );
  OAI211XL U42764 ( .A0(n33592), .A1(n42738), .B0(n16705), .C0(n16706), .Y(
        n35741) );
  OA22XL U42765 ( .A0(net262304), .A1(n33576), .B0(n33584), .B1(n40128), .Y(
        n16705) );
  OAI211XL U42766 ( .A0(n33584), .A1(n42739), .B0(n16681), .C0(n16682), .Y(
        n35733) );
  OA22XL U42767 ( .A0(net262323), .A1(n33568), .B0(n33576), .B1(n40127), .Y(
        n16681) );
  OAI211XL U42768 ( .A0(n33617), .A1(n42736), .B0(n16780), .C0(n16781), .Y(
        n35766) );
  OA22XL U42769 ( .A0(net262285), .A1(n33601), .B0(n33609), .B1(n40078), .Y(
        n16780) );
  OAI211XL U42770 ( .A0(n33593), .A1(n42738), .B0(n16708), .C0(n16709), .Y(
        n35742) );
  OA22XL U42771 ( .A0(net262304), .A1(n33577), .B0(n33585), .B1(n40128), .Y(
        n16708) );
  OAI211XL U42772 ( .A0(n33585), .A1(n42739), .B0(n16684), .C0(n16685), .Y(
        n35734) );
  OA22XL U42773 ( .A0(net262323), .A1(n33569), .B0(n33577), .B1(n40127), .Y(
        n16684) );
  OAI211XL U42774 ( .A0(n33604), .A1(n42737), .B0(n16741), .C0(n16742), .Y(
        n35753) );
  OA22XL U42775 ( .A0(net262304), .A1(n33588), .B0(n33596), .B1(net218762),
        .Y(n16741) );
  OAI211XL U42776 ( .A0(n33580), .A1(n42740), .B0(n16669), .C0(n16670), .Y(
        n35729) );
  OA22XL U42777 ( .A0(net262323), .A1(n33564), .B0(n33572), .B1(n40127), .Y(
        n16669) );
  OAI211XL U42778 ( .A0(n33605), .A1(n42737), .B0(n16744), .C0(n16745), .Y(
        n35754) );
  OA22XL U42779 ( .A0(net262304), .A1(n33589), .B0(n33597), .B1(n40093), .Y(
        n16744) );
  OAI211XL U42780 ( .A0(n33597), .A1(n42834), .B0(n16720), .C0(n16721), .Y(
        n35746) );
  OA22XL U42781 ( .A0(net262304), .A1(n33581), .B0(n33589), .B1(n40128), .Y(
        n16720) );
  OAI211XL U42782 ( .A0(n33581), .A1(n42740), .B0(n16672), .C0(n16673), .Y(
        n35730) );
  OA22XL U42783 ( .A0(net262323), .A1(n33565), .B0(n33573), .B1(n40127), .Y(
        n16672) );
  OAI211XL U42784 ( .A0(n33606), .A1(n42737), .B0(n16747), .C0(n16748), .Y(
        n35755) );
  OA22XL U42785 ( .A0(net262285), .A1(n33590), .B0(n33598), .B1(net218748),
        .Y(n16747) );
  OAI211XL U42786 ( .A0(n33598), .A1(n42849), .B0(n16723), .C0(n16724), .Y(
        n35747) );
  OA22XL U42787 ( .A0(net262304), .A1(n33582), .B0(n33590), .B1(n40128), .Y(
        n16723) );
  OAI211XL U42788 ( .A0(n33582), .A1(n42740), .B0(n16675), .C0(n16676), .Y(
        n35731) );
  OA22XL U42789 ( .A0(net262323), .A1(n33566), .B0(n33574), .B1(n40127), .Y(
        n16675) );
  OAI211XL U42790 ( .A0(n33608), .A1(n42737), .B0(n16753), .C0(n16754), .Y(
        n35757) );
  OA22XL U42791 ( .A0(net262285), .A1(n33592), .B0(n33600), .B1(net218780),
        .Y(n16753) );
  OAI211XL U42792 ( .A0(n33600), .A1(n42864), .B0(n16729), .C0(n16730), .Y(
        n35749) );
  OA22XL U42793 ( .A0(net262304), .A1(n33584), .B0(n33592), .B1(n40128), .Y(
        n16729) );
  OAI211XL U42794 ( .A0(n33576), .A1(n42740), .B0(n16657), .C0(n16658), .Y(
        n35725) );
  OA22XL U42795 ( .A0(net262323), .A1(n33560), .B0(n33568), .B1(n40127), .Y(
        n16657) );
  OAI211XL U42796 ( .A0(n33609), .A1(n42737), .B0(n16756), .C0(n16757), .Y(
        n35758) );
  OA22XL U42797 ( .A0(net262285), .A1(n33593), .B0(n33601), .B1(net218786),
        .Y(n16756) );
  OAI211XL U42798 ( .A0(n33601), .A1(n42838), .B0(n16732), .C0(n16733), .Y(
        n35750) );
  OA22XL U42799 ( .A0(net262304), .A1(n33585), .B0(n33593), .B1(n40128), .Y(
        n16732) );
  OAI211XL U42800 ( .A0(n33577), .A1(n42740), .B0(n16660), .C0(n16661), .Y(
        n35726) );
  OA22XL U42801 ( .A0(net262323), .A1(n33561), .B0(n33569), .B1(n40127), .Y(
        n16660) );
  OAI211XL U42802 ( .A0(n32948), .A1(n42991), .B0(n14773), .C0(n14774), .Y(
        n35097) );
  OAI211XL U42803 ( .A0(n32945), .A1(n42991), .B0(n14764), .C0(n14765), .Y(
        n35094) );
  XOR2XL U42804 ( .A(n36768), .B(n32873), .Y(n46626) );
  XOR2XL U42805 ( .A(n36773), .B(n32881), .Y(n46624) );
  XOR2XL U42806 ( .A(n32841), .B(n36780), .Y(n45573) );
  XOR2XL U42807 ( .A(n36764), .B(n32889), .Y(n46623) );
  XOR2XL U42808 ( .A(n32993), .B(n36780), .Y(n46076) );
  XOR2XL U42809 ( .A(n32948), .B(n36827), .Y(n43462) );
  XOR2XL U42810 ( .A(n41300), .B(n32932), .Y(n46087) );
  XOR2XL U42811 ( .A(n41303), .B(n32916), .Y(n46086) );
  XOR2XL U42812 ( .A(n41304), .B(n32948), .Y(n46085) );
  NOR2XL U42813 ( .A(n10903), .B(n46858), .Y(net211773) );
  XOR2XL U42814 ( .A(n36740), .B(n32940), .Y(n46858) );
  XOR2XL U42815 ( .A(n32956), .B(n36824), .Y(n43463) );
  XOR2XL U42816 ( .A(n32852), .B(n36827), .Y(n43495) );
  XOR2XL U42817 ( .A(n32916), .B(n36823), .Y(n43437) );
  XOR2XL U42818 ( .A(n36743), .B(n32948), .Y(n46856) );
  XOR2XL U42819 ( .A(n32908), .B(n36831), .Y(n43477) );
  XOR2XL U42820 ( .A(n32972), .B(n36825), .Y(n43457) );
  XOR2XL U42821 ( .A(n32980), .B(n36827), .Y(n43418) );
  XOR2XL U42822 ( .A(n36764), .B(n32833), .Y(n46634) );
  XOR2XL U42823 ( .A(n32969), .B(n36778), .Y(n46079) );
  XOR2XL U42824 ( .A(n36748), .B(n32964), .Y(n46849) );
  XOR2XL U42825 ( .A(n32996), .B(n36823), .Y(n43409) );
  XOR2XL U42826 ( .A(n32849), .B(n36779), .Y(n46628) );
  XOR2XL U42827 ( .A(n32860), .B(n36824), .Y(n46627) );
  XOR2XL U42828 ( .A(n33004), .B(n36831), .Y(n43428) );
  XOR2XL U42829 ( .A(n41302), .B(n32956), .Y(n46078) );
  XOR2XL U42830 ( .A(n41302), .B(n32924), .Y(n47753) );
  XOR2XL U42831 ( .A(n36740), .B(n32956), .Y(n46855) );
  XOR2XL U42832 ( .A(n32889), .B(n36778), .Y(n45585) );
  XOR2XL U42833 ( .A(n32932), .B(n36827), .Y(n43448) );
  XOR2XL U42834 ( .A(n36741), .B(n32916), .Y(n47758) );
  XOR2XL U42835 ( .A(n32985), .B(n36776), .Y(n47792) );
  XOR2XL U42836 ( .A(n32900), .B(n36831), .Y(n43486) );
  XOR2XL U42837 ( .A(n32849), .B(n36770), .Y(n46615) );
  XOR2XL U42838 ( .A(n36773), .B(n32977), .Y(n47797) );
  XOR2XL U42839 ( .A(n36767), .B(n32897), .Y(n46618) );
  XOR2XL U42840 ( .A(n32940), .B(n36824), .Y(n43447) );
  XOR2XL U42841 ( .A(n32884), .B(n36825), .Y(n43487) );
  XOR2XL U42842 ( .A(n36740), .B(n32932), .Y(n46859) );
  XOR2XL U42843 ( .A(n36773), .B(n32865), .Y(n46625) );
  XOR2XL U42844 ( .A(n41302), .B(n32964), .Y(n46077) );
  XOR2XL U42845 ( .A(n41301), .B(n32908), .Y(n45582) );
  XOR2XL U42846 ( .A(n32964), .B(n36825), .Y(n43468) );
  XOR2XL U42847 ( .A(n32988), .B(n36822), .Y(n43423) );
  XOR2XL U42848 ( .A(n32924), .B(n36831), .Y(n43442) );
  XOR2XL U42849 ( .A(n41303), .B(n32940), .Y(n46080) );
  NOR2XL U42850 ( .A(n10807), .B(n46854), .Y(net211793) );
  XOR2XL U42851 ( .A(n36768), .B(n32969), .Y(n46854) );
  XOR2XL U42852 ( .A(n36742), .B(n32908), .Y(n46617) );
  NOR2XL U42853 ( .A(n10808), .B(n46699), .Y(n46703) );
  XOR2XL U42854 ( .A(n32985), .B(n36773), .Y(n46699) );
  XOR2XL U42855 ( .A(n32892), .B(n36829), .Y(n43492) );
  XOR2XL U42856 ( .A(n32857), .B(n36786), .Y(n46610) );
  XOR2XL U42857 ( .A(n36741), .B(n32924), .Y(n46857) );
  NAND2XL U42858 ( .A(n9875), .B(n9986), .Y(n48554) );
  NOR2XL U42859 ( .A(n9677), .B(net266151), .Y(n47950) );
  AOI2BB2XL U42860 ( .B0(net264652), .B1(n48568), .A0N(net217184), .A1N(n34388), .Y(n48569) );
  OA22XL U42861 ( .A0(net262551), .A1(n34364), .B0(n34372), .B1(n40117), .Y(
        n19069) );
  AOI2BB2XL U42862 ( .B0(net264652), .B1(n41387), .A0N(net217212), .A1N(n34380), .Y(n48572) );
  OA22XL U42863 ( .A0(net262570), .A1(n34356), .B0(n34364), .B1(n40117), .Y(
        n19045) );
  AOI2BB2XL U42864 ( .B0(net265245), .B1(n48575), .A0N(n40290), .A1N(n34372),
        .Y(n48576) );
  OA22XL U42865 ( .A0(net262570), .A1(n34348), .B0(n34356), .B1(n40116), .Y(
        n19021) );
  AOI2BB2XL U42866 ( .B0(net265378), .B1(n48579), .A0N(n40314), .A1N(n34364),
        .Y(n48580) );
  OA22XL U42867 ( .A0(net262589), .A1(n34340), .B0(n34348), .B1(n40116), .Y(
        n18997) );
  AOI2BB2XL U42868 ( .B0(net221802), .B1(n48583), .A0N(n40280), .A1N(n34356),
        .Y(n48584) );
  OA22XL U42869 ( .A0(net262589), .A1(n34332), .B0(n34340), .B1(n40115), .Y(
        n18973) );
  AOI2BB2XL U42870 ( .B0(net265188), .B1(n41270), .A0N(n40280), .A1N(n34348),
        .Y(n48587) );
  OA22XL U42871 ( .A0(net262608), .A1(n34324), .B0(n34332), .B1(n40115), .Y(
        n18949) );
  AOI2BB2XL U42872 ( .B0(net265169), .B1(n48590), .A0N(n40280), .A1N(n34340),
        .Y(n48591) );
  OA22XL U42873 ( .A0(net262608), .A1(n34316), .B0(n34324), .B1(n40114), .Y(
        n18925) );
  AOI2BB2XL U42874 ( .B0(net265169), .B1(n48594), .A0N(n40280), .A1N(n34332),
        .Y(n48595) );
  OA22XL U42875 ( .A0(net262608), .A1(n34308), .B0(n34316), .B1(n40114), .Y(
        n18901) );
  AOI2BB2XL U42876 ( .B0(net264979), .B1(n48598), .A0N(n40280), .A1N(n34324),
        .Y(n48599) );
  OA22XL U42877 ( .A0(net262627), .A1(n34300), .B0(n34308), .B1(n40113), .Y(
        n18877) );
  AOI2BB2XL U42878 ( .B0(net265112), .B1(n48602), .A0N(n40280), .A1N(n34316),
        .Y(n48603) );
  OA22XL U42879 ( .A0(net262627), .A1(n34292), .B0(n34300), .B1(n40113), .Y(
        n18853) );
  AOI2BB2XL U42880 ( .B0(net265378), .B1(n48614), .A0N(n40280), .A1N(n34292),
        .Y(n48615) );
  OA22XL U42881 ( .A0(net262380), .A1(n34268), .B0(n34276), .B1(n40123), .Y(
        n18781) );
  AOI2BB2XL U42882 ( .B0(net265245), .B1(n48618), .A0N(n40280), .A1N(n34284),
        .Y(n48619) );
  OA22XL U42883 ( .A0(net262399), .A1(n34260), .B0(n34268), .B1(n40123), .Y(
        n18757) );
  AOI2BB2XL U42884 ( .B0(net264682), .B1(n48630), .A0N(n40280), .A1N(n34260),
        .Y(n48631) );
  OA22XL U42885 ( .A0(net262418), .A1(n34236), .B0(n34244), .B1(n40121), .Y(
        n18685) );
  AOI2BB2XL U42886 ( .B0(net264682), .B1(n48634), .A0N(n40280), .A1N(n34252),
        .Y(n48635) );
  OA22XL U42887 ( .A0(net262437), .A1(n34228), .B0(n34236), .B1(n40121), .Y(
        n18661) );
  AOI2BB2XL U42888 ( .B0(net265682), .B1(n48884), .A0N(n40284), .A1N(n34390),
        .Y(n48885) );
  OA22XL U42889 ( .A0(net262551), .A1(n34366), .B0(n34374), .B1(n40117), .Y(
        n19075) );
  AOI2BB2XL U42890 ( .B0(net264903), .B1(n49062), .A0N(n40278), .A1N(n34336),
        .Y(n49063) );
  OA22XL U42891 ( .A0(net262608), .A1(n34312), .B0(n34320), .B1(n40114), .Y(
        n18913) );
  AOI2BB2XL U42892 ( .B0(net264903), .B1(n49082), .A0N(n40278), .A1N(n34296),
        .Y(n49083) );
  OA22XL U42893 ( .A0(net262646), .A1(n34272), .B0(n34280), .B1(n40086), .Y(
        n18793) );
  AOI2BB2XL U42894 ( .B0(net264846), .B1(n49086), .A0N(n40278), .A1N(n34288),
        .Y(n49087) );
  OA22XL U42895 ( .A0(net262399), .A1(n34264), .B0(n34272), .B1(n40123), .Y(
        n18769) );
  AOI2BB2XL U42896 ( .B0(net264846), .B1(n49098), .A0N(n40278), .A1N(n34264),
        .Y(n49099) );
  OA22XL U42897 ( .A0(net262418), .A1(n34240), .B0(n34248), .B1(n40121), .Y(
        n18697) );
  AOI2BB2XL U42898 ( .B0(net264903), .B1(n49102), .A0N(n40278), .A1N(n34256),
        .Y(n49103) );
  OA22XL U42899 ( .A0(net262418), .A1(n34232), .B0(n34240), .B1(n40121), .Y(
        n18673) );
  AOI2BB2XL U42900 ( .B0(net264577), .B1(n49192), .A0N(n40287), .A1N(n34385),
        .Y(n49193) );
  OA22XL U42901 ( .A0(net262551), .A1(n34361), .B0(n34369), .B1(n40117), .Y(
        n19060) );
  AOI2BB2XL U42902 ( .B0(net265549), .B1(n49347), .A0N(n40279), .A1N(n34386),
        .Y(n49348) );
  OA22XL U42903 ( .A0(net262551), .A1(n34362), .B0(n34370), .B1(n40117), .Y(
        n19063) );
  AOI2BB2XL U42904 ( .B0(net264846), .B1(n41349), .A0N(n40287), .A1N(n34352),
        .Y(n49055) );
  OA22XL U42905 ( .A0(net262589), .A1(n34328), .B0(n34336), .B1(n40115), .Y(
        n18961) );
  NAND2XL U42906 ( .A(n43009), .B(n49070), .Y(n49060) );
  AOI2BB2XL U42907 ( .B0(net264846), .B1(n49058), .A0N(net217218), .A1N(n34344), .Y(n49059) );
  OA22XL U42908 ( .A0(net262608), .A1(n34320), .B0(n34328), .B1(n40114), .Y(
        n18937) );
  AOI2BB2XL U42909 ( .B0(net264903), .B1(n49066), .A0N(n40289), .A1N(n34328),
        .Y(n49067) );
  OA22XL U42910 ( .A0(net262627), .A1(n34304), .B0(n34312), .B1(n40113), .Y(
        n18889) );
  AOI2BB2XL U42911 ( .B0(net264846), .B1(n49070), .A0N(n40310), .A1N(n34320),
        .Y(n49071) );
  OA22XL U42912 ( .A0(net262627), .A1(n34296), .B0(n34304), .B1(n40113), .Y(
        n18865) );
  NAND2XL U42913 ( .A(n43009), .B(n49047), .Y(n49037) );
  AOI2BB2XL U42914 ( .B0(net264532), .B1(n41234), .A0N(n40306), .A1N(n34392),
        .Y(n49036) );
  OA22XL U42915 ( .A0(net262551), .A1(n34368), .B0(n34376), .B1(n40117), .Y(
        n19081) );
  NAND2XL U42916 ( .A(n43009), .B(n49051), .Y(n49041) );
  AOI2BB2XL U42917 ( .B0(net264532), .B1(n49039), .A0N(n40309), .A1N(n34384),
        .Y(n49040) );
  OA22XL U42918 ( .A0(net262551), .A1(n34360), .B0(n34368), .B1(n40117), .Y(
        n19057) );
  NAND2XL U42919 ( .A(n43009), .B(n41349), .Y(n49045) );
  AOI2BB2XL U42920 ( .B0(net264532), .B1(n49043), .A0N(n40306), .A1N(n34376),
        .Y(n49044) );
  OA22XL U42921 ( .A0(net262570), .A1(n34352), .B0(n34360), .B1(n40116), .Y(
        n19033) );
  NAND2XL U42922 ( .A(n43009), .B(n49058), .Y(n49049) );
  AOI2BB2XL U42923 ( .B0(net264532), .B1(n49047), .A0N(n40292), .A1N(n34368),
        .Y(n49048) );
  OA22XL U42924 ( .A0(net262570), .A1(n34344), .B0(n34352), .B1(n40116), .Y(
        n19009) );
  NAND2XL U42925 ( .A(n43009), .B(n49062), .Y(n49053) );
  AOI2BB2XL U42926 ( .B0(net264532), .B1(n49051), .A0N(n40287), .A1N(n34360),
        .Y(n49052) );
  OA22XL U42927 ( .A0(net262589), .A1(n34336), .B0(n34344), .B1(n40115), .Y(
        n18985) );
  AOI2BB2XL U42928 ( .B0(net264742), .B1(n48802), .A0N(n40282), .A1N(n34237),
        .Y(n48803) );
  OA22XL U42929 ( .A0(net262437), .A1(n34213), .B0(n34221), .B1(n40120), .Y(
        n18616) );
  AOI2BB2XL U42930 ( .B0(net264742), .B1(n48806), .A0N(n40283), .A1N(n34229),
        .Y(n48807) );
  OA22XL U42931 ( .A0(net262456), .A1(n34205), .B0(n34213), .B1(n40046), .Y(
        n18592) );
  AOI2BB2XL U42932 ( .B0(net264712), .B1(n48810), .A0N(n40283), .A1N(n34221),
        .Y(n48811) );
  OA22XL U42933 ( .A0(net262456), .A1(n34197), .B0(n34205), .B1(n40053), .Y(
        n18568) );
  AOI2BB2XL U42934 ( .B0(net264742), .B1(n48814), .A0N(n40283), .A1N(n34213),
        .Y(n48815) );
  OA22XL U42935 ( .A0(net262475), .A1(n34189), .B0(n34197), .B1(n40119), .Y(
        n18544) );
  AOI2BB2XL U42936 ( .B0(net264712), .B1(n48818), .A0N(n40283), .A1N(n34205),
        .Y(n48819) );
  OA22XL U42937 ( .A0(net262475), .A1(n34181), .B0(n34189), .B1(n40119), .Y(
        n18520) );
  AOI2BB2XL U42938 ( .B0(net264712), .B1(n48822), .A0N(n40283), .A1N(n34197),
        .Y(n48823) );
  OA22XL U42939 ( .A0(net263596), .A1(n34173), .B0(n34181), .B1(n40055), .Y(
        n18496) );
  AOI2BB2XL U42940 ( .B0(net264742), .B1(n48830), .A0N(n40283), .A1N(n34181),
        .Y(n48831) );
  OA22XL U42941 ( .A0(net262513), .A1(n34157), .B0(n34165), .B1(n40118), .Y(
        n18448) );
  AOI2BB2XL U42942 ( .B0(net221718), .B1(n48834), .A0N(n40283), .A1N(n34173),
        .Y(n48835) );
  OA22XL U42943 ( .A0(net262513), .A1(n34149), .B0(n34157), .B1(n40118), .Y(
        n18424) );
  AOI2BB2XL U42944 ( .B0(net264712), .B1(n48838), .A0N(n40283), .A1N(n34165),
        .Y(n48839) );
  OA22XL U42945 ( .A0(net262798), .A1(n41801), .B0(n34149), .B1(n40106), .Y(
        n18400) );
  AOI2BB2XL U42946 ( .B0(net264712), .B1(n48846), .A0N(n40283), .A1N(n34149),
        .Y(n48847) );
  OA22XL U42947 ( .A0(net262817), .A1(n34125), .B0(n41802), .B1(n40105), .Y(
        n18352) );
  AOI2BB2XL U42948 ( .B0(net264742), .B1(n48854), .A0N(n40283), .A1N(n41802),
        .Y(n48855) );
  OA22XL U42949 ( .A0(net262817), .A1(n34109), .B0(n34117), .B1(n40074), .Y(
        n18304) );
  AOI2BB2XL U42950 ( .B0(net264652), .B1(n48561), .A0N(net217272), .A1N(n34404), .Y(n48562) );
  OA22XL U42951 ( .A0(net262532), .A1(n34380), .B0(n34388), .B1(n40079), .Y(
        n19117) );
  AOI2BB2XL U42952 ( .B0(net264979), .B1(n48606), .A0N(n40280), .A1N(n34308),
        .Y(n48607) );
  OA22XL U42953 ( .A0(net262646), .A1(n34284), .B0(n34292), .B1(n40112), .Y(
        n18829) );
  AOI2BB2XL U42954 ( .B0(net265226), .B1(n48610), .A0N(n40280), .A1N(n34300),
        .Y(n48611) );
  OA22XL U42955 ( .A0(net262646), .A1(n34276), .B0(n34284), .B1(n40112), .Y(
        n18805) );
  AOI2BB2XL U42956 ( .B0(net265150), .B1(n48622), .A0N(n40280), .A1N(n34276),
        .Y(n48623) );
  OA22XL U42957 ( .A0(net262399), .A1(n34252), .B0(n34260), .B1(n40122), .Y(
        n18733) );
  AOI2BB2XL U42958 ( .B0(net221810), .B1(n48626), .A0N(n40280), .A1N(n34268),
        .Y(n48627) );
  OA22XL U42959 ( .A0(net262418), .A1(n34244), .B0(n34252), .B1(n40122), .Y(
        n18709) );
  AOI2BB2XL U42960 ( .B0(net264682), .B1(n48638), .A0N(n40280), .A1N(n34244),
        .Y(n48639) );
  OA22XL U42961 ( .A0(net262437), .A1(n34220), .B0(n34228), .B1(n40120), .Y(
        n18637) );
  AOI2BB2XL U42962 ( .B0(net264682), .B1(n48642), .A0N(n40280), .A1N(n34236),
        .Y(n48643) );
  OA22XL U42963 ( .A0(net262456), .A1(n34212), .B0(n34220), .B1(n40120), .Y(
        n18613) );
  AOI2BB2XL U42964 ( .B0(net264682), .B1(n48646), .A0N(n40280), .A1N(n34228),
        .Y(n48647) );
  OA22XL U42965 ( .A0(net262456), .A1(n34204), .B0(n34212), .B1(n40054), .Y(
        n18589) );
  AOI2BB2XL U42966 ( .B0(net264682), .B1(n48650), .A0N(n40280), .A1N(n34220),
        .Y(n48651) );
  OA22XL U42967 ( .A0(net262456), .A1(n34196), .B0(n34204), .B1(n40042), .Y(
        n18565) );
  AOI2BB2XL U42968 ( .B0(net264682), .B1(n48654), .A0N(n40280), .A1N(n34212),
        .Y(n48655) );
  OA22XL U42969 ( .A0(net262475), .A1(n34188), .B0(n34196), .B1(n40119), .Y(
        n18541) );
  AOI2BB2XL U42970 ( .B0(net264682), .B1(n48658), .A0N(n40281), .A1N(n34204),
        .Y(n48659) );
  OA22XL U42971 ( .A0(net262475), .A1(n34180), .B0(n34188), .B1(n40119), .Y(
        n18517) );
  AOI2BB2XL U42972 ( .B0(net264682), .B1(n48662), .A0N(n40281), .A1N(n34196),
        .Y(n48663) );
  OA22XL U42973 ( .A0(net263596), .A1(n34172), .B0(n34180), .B1(n40055), .Y(
        n18493) );
  AOI2BB2XL U42974 ( .B0(net264682), .B1(n48666), .A0N(n40281), .A1N(n34188),
        .Y(n48667) );
  OA22XL U42975 ( .A0(net263406), .A1(n34164), .B0(n34172), .B1(n40128), .Y(
        n18469) );
  AOI2BB2XL U42976 ( .B0(net264682), .B1(n48670), .A0N(n40281), .A1N(n34180),
        .Y(n48671) );
  OA22XL U42977 ( .A0(net262513), .A1(n34156), .B0(n34164), .B1(n40118), .Y(
        n18445) );
  AOI2BB2XL U42978 ( .B0(net264682), .B1(n48674), .A0N(n40281), .A1N(n34172),
        .Y(n48675) );
  OA22XL U42979 ( .A0(net262513), .A1(n34148), .B0(n34156), .B1(n40118), .Y(
        n18421) );
  AOI2BB2XL U42980 ( .B0(net264682), .B1(n48678), .A0N(n40281), .A1N(n34164),
        .Y(n48679) );
  OA22XL U42981 ( .A0(net262798), .A1(n34140), .B0(n34148), .B1(n40106), .Y(
        n18397) );
  AOI2BB2XL U42982 ( .B0(net264682), .B1(n48682), .A0N(n40281), .A1N(n34156),
        .Y(n48683) );
  OA22XL U42983 ( .A0(net262798), .A1(n41799), .B0(n34140), .B1(n40106), .Y(
        n18373) );
  AOI2BB2XL U42984 ( .B0(net265530), .B1(n48686), .A0N(n40281), .A1N(n34148),
        .Y(n48687) );
  OA22XL U42985 ( .A0(net262817), .A1(n34124), .B0(n41799), .B1(n40105), .Y(
        n18349) );
  AOI2BB2XL U42986 ( .B0(net265150), .B1(n48690), .A0N(n40281), .A1N(n34140),
        .Y(n48691) );
  OA22XL U42987 ( .A0(net262817), .A1(n34116), .B0(n34124), .B1(n40105), .Y(
        n18325) );
  AOI2BB2XL U42988 ( .B0(net265226), .B1(n48694), .A0N(n40281), .A1N(n41799),
        .Y(n48695) );
  OA22XL U42989 ( .A0(net262836), .A1(n34108), .B0(n34116), .B1(n40082), .Y(
        n18301) );
  AOI2BB2XL U42990 ( .B0(net265416), .B1(n48698), .A0N(n40281), .A1N(n34124),
        .Y(n48699) );
  OA22XL U42991 ( .A0(net262836), .A1(n34100), .B0(n34108), .B1(n40073), .Y(
        n18277) );
  OA22XL U42992 ( .A0(net262855), .A1(n34084), .B0(n34092), .B1(n40104), .Y(
        n18229) );
  AOI2BB2XL U42993 ( .B0(net265511), .B1(n41643), .A0N(n40281), .A1N(n34405),
        .Y(n48720) );
  OA22XL U42994 ( .A0(net262532), .A1(n34381), .B0(n34389), .B1(n40070), .Y(
        n19120) );
  AOI2BB2XL U42995 ( .B0(net265169), .B1(n48726), .A0N(n40281), .A1N(n34389),
        .Y(n48727) );
  OA22XL U42996 ( .A0(net262551), .A1(n34365), .B0(n34373), .B1(n40117), .Y(
        n19072) );
  AOI2BB2XL U42997 ( .B0(net265378), .B1(n48730), .A0N(n40281), .A1N(n34381),
        .Y(n48731) );
  OA22XL U42998 ( .A0(net262570), .A1(n34357), .B0(n34365), .B1(n40117), .Y(
        n19048) );
  AOI2BB2XL U42999 ( .B0(net265492), .B1(n48734), .A0N(n40282), .A1N(n34373),
        .Y(n48735) );
  OA22XL U43000 ( .A0(net262570), .A1(n34349), .B0(n34357), .B1(n40116), .Y(
        n19024) );
  AOI2BB2XL U43001 ( .B0(net265511), .B1(n48738), .A0N(n40282), .A1N(n34365),
        .Y(n48739) );
  OA22XL U43002 ( .A0(net262589), .A1(n34341), .B0(n34349), .B1(n40116), .Y(
        n19000) );
  AOI2BB2XL U43003 ( .B0(net265188), .B1(n48742), .A0N(n40282), .A1N(n34357),
        .Y(n48743) );
  OA22XL U43004 ( .A0(net262589), .A1(n34333), .B0(n34341), .B1(n40115), .Y(
        n18976) );
  AOI2BB2XL U43005 ( .B0(net264712), .B1(n48746), .A0N(n40282), .A1N(n34349),
        .Y(n48747) );
  OA22XL U43006 ( .A0(net262589), .A1(n34325), .B0(n34333), .B1(n40115), .Y(
        n18952) );
  AOI2BB2XL U43007 ( .B0(net264712), .B1(n48750), .A0N(n40282), .A1N(n34341),
        .Y(n48751) );
  OA22XL U43008 ( .A0(net262608), .A1(n34317), .B0(n34325), .B1(n40114), .Y(
        n18928) );
  AOI2BB2XL U43009 ( .B0(net264712), .B1(n48754), .A0N(n40282), .A1N(n34333),
        .Y(n48755) );
  OA22XL U43010 ( .A0(net262608), .A1(n34309), .B0(n34317), .B1(n40114), .Y(
        n18904) );
  AOI2BB2XL U43011 ( .B0(net264712), .B1(n48758), .A0N(n40282), .A1N(n34325),
        .Y(n48759) );
  OA22XL U43012 ( .A0(net262627), .A1(n34301), .B0(n34309), .B1(n40113), .Y(
        n18880) );
  AOI2BB2XL U43013 ( .B0(net264712), .B1(n48762), .A0N(n40282), .A1N(n34317),
        .Y(n48763) );
  OA22XL U43014 ( .A0(net262627), .A1(n34293), .B0(n34301), .B1(n40113), .Y(
        n18856) );
  AOI2BB2XL U43015 ( .B0(net264712), .B1(n48766), .A0N(n40282), .A1N(n34309),
        .Y(n48767) );
  OA22XL U43016 ( .A0(net262646), .A1(n34285), .B0(n34293), .B1(n40112), .Y(
        n18832) );
  AOI2BB2XL U43017 ( .B0(net264712), .B1(n48770), .A0N(n40282), .A1N(n34301),
        .Y(n48771) );
  OA22XL U43018 ( .A0(net262646), .A1(n34277), .B0(n34285), .B1(n40112), .Y(
        n18808) );
  AOI2BB2XL U43019 ( .B0(net264712), .B1(n48774), .A0N(n40282), .A1N(n34293),
        .Y(n48775) );
  OA22XL U43020 ( .A0(net262380), .A1(n34269), .B0(n34277), .B1(n40123), .Y(
        n18784) );
  AOI2BB2XL U43021 ( .B0(net264712), .B1(n48778), .A0N(n40282), .A1N(n34285),
        .Y(n48779) );
  OA22XL U43022 ( .A0(net262399), .A1(n34261), .B0(n34269), .B1(n40123), .Y(
        n18760) );
  AOI2BB2XL U43023 ( .B0(net264712), .B1(n48782), .A0N(n40282), .A1N(n34277),
        .Y(n48783) );
  OA22XL U43024 ( .A0(net262399), .A1(n34253), .B0(n34261), .B1(n40122), .Y(
        n18736) );
  AOI2BB2XL U43025 ( .B0(net264712), .B1(n48786), .A0N(n40282), .A1N(n34269),
        .Y(n48787) );
  OA22XL U43026 ( .A0(net262418), .A1(n34245), .B0(n34253), .B1(n40122), .Y(
        n18712) );
  AOI2BB2XL U43027 ( .B0(net264712), .B1(n48790), .A0N(n40282), .A1N(n34261),
        .Y(n48791) );
  OA22XL U43028 ( .A0(net262418), .A1(n34237), .B0(n34245), .B1(n40121), .Y(
        n18688) );
  AOI2BB2XL U43029 ( .B0(net264712), .B1(n48794), .A0N(n40282), .A1N(n34253),
        .Y(n48795) );
  OA22XL U43030 ( .A0(net262437), .A1(n34229), .B0(n34237), .B1(n40121), .Y(
        n18664) );
  AOI2BB2XL U43031 ( .B0(net264712), .B1(n48798), .A0N(n40282), .A1N(n34245),
        .Y(n48799) );
  OA22XL U43032 ( .A0(net262437), .A1(n34221), .B0(n34229), .B1(n40120), .Y(
        n18640) );
  AOI2BB2XL U43033 ( .B0(net265739), .B1(n48826), .A0N(n40283), .A1N(n34189),
        .Y(n48827) );
  OA22XL U43034 ( .A0(net262798), .A1(n34165), .B0(n34173), .B1(n40093), .Y(
        n18472) );
  AOI2BB2XL U43035 ( .B0(net265796), .B1(n48842), .A0N(n40283), .A1N(n34157),
        .Y(n48843) );
  OA22XL U43036 ( .A0(net262798), .A1(n41802), .B0(n41801), .B1(n40106), .Y(
        n18376) );
  AOI2BB2XL U43037 ( .B0(net265644), .B1(n48850), .A0N(n40283), .A1N(n41801),
        .Y(n48851) );
  OA22XL U43038 ( .A0(net262817), .A1(n34117), .B0(n34125), .B1(n40105), .Y(
        n18328) );
  AOI2BB2XL U43039 ( .B0(net265777), .B1(n48864), .A0N(n40283), .A1N(n34109),
        .Y(n48865) );
  OA22XL U43040 ( .A0(net262855), .A1(n34085), .B0(n34093), .B1(n40104), .Y(
        n18232) );
  AOI2BB2XL U43041 ( .B0(net265644), .B1(n41345), .A0N(n40284), .A1N(n34406),
        .Y(n48878) );
  OA22XL U43042 ( .A0(net262532), .A1(n34382), .B0(n34390), .B1(n40093), .Y(
        n19123) );
  AOI2BB2XL U43043 ( .B0(net264979), .B1(n41367), .A0N(n40284), .A1N(n34382),
        .Y(n48888) );
  OA22XL U43044 ( .A0(net262570), .A1(n34358), .B0(n34366), .B1(n40117), .Y(
        n19051) );
  AOI2BB2XL U43045 ( .B0(net265625), .B1(n48891), .A0N(n40284), .A1N(n34374),
        .Y(n48892) );
  OA22XL U43046 ( .A0(net262570), .A1(n34350), .B0(n34358), .B1(n40116), .Y(
        n19027) );
  AOI2BB2XL U43047 ( .B0(net265739), .B1(n48895), .A0N(n40284), .A1N(n34366),
        .Y(n48896) );
  OA22XL U43048 ( .A0(net262570), .A1(n34342), .B0(n34350), .B1(n40116), .Y(
        n19003) );
  AOI2BB2XL U43049 ( .B0(net265682), .B1(n41655), .A0N(n40284), .A1N(n34358),
        .Y(n48899) );
  OA22XL U43050 ( .A0(net262589), .A1(n34334), .B0(n34342), .B1(n40115), .Y(
        n18979) );
  AOI2BB2XL U43051 ( .B0(net264742), .B1(n48902), .A0N(n40284), .A1N(n34350),
        .Y(n48903) );
  OA22XL U43052 ( .A0(net262589), .A1(n34326), .B0(n34334), .B1(n40115), .Y(
        n18955) );
  AOI2BB2XL U43053 ( .B0(net264742), .B1(n48906), .A0N(n40284), .A1N(n34342),
        .Y(n48907) );
  OA22XL U43054 ( .A0(net262608), .A1(n34318), .B0(n34326), .B1(n40114), .Y(
        n18931) );
  AOI2BB2XL U43055 ( .B0(net264742), .B1(n48910), .A0N(n40284), .A1N(n34334),
        .Y(n48911) );
  OA22XL U43056 ( .A0(net262608), .A1(n34310), .B0(n34318), .B1(n40114), .Y(
        n18907) );
  AOI2BB2XL U43057 ( .B0(net264742), .B1(n48914), .A0N(n40284), .A1N(n34326),
        .Y(n48915) );
  OA22XL U43058 ( .A0(net262627), .A1(n34302), .B0(n34310), .B1(n40113), .Y(
        n18883) );
  AOI2BB2XL U43059 ( .B0(net264742), .B1(n48918), .A0N(n40284), .A1N(n34318),
        .Y(n48919) );
  OA22XL U43060 ( .A0(net262627), .A1(n34294), .B0(n34302), .B1(n40113), .Y(
        n18859) );
  AOI2BB2XL U43061 ( .B0(net264742), .B1(n48922), .A0N(n40284), .A1N(n34310),
        .Y(n48923) );
  OA22XL U43062 ( .A0(net262646), .A1(n34286), .B0(n34294), .B1(n40112), .Y(
        n18835) );
  AOI2BB2XL U43063 ( .B0(net264742), .B1(n48926), .A0N(n40284), .A1N(n34302),
        .Y(n48927) );
  OA22XL U43064 ( .A0(net262646), .A1(n34278), .B0(n34286), .B1(n40112), .Y(
        n18811) );
  AOI2BB2XL U43065 ( .B0(net264742), .B1(n48930), .A0N(n40284), .A1N(n34294),
        .Y(n48931) );
  OA22XL U43066 ( .A0(net262380), .A1(n34270), .B0(n34278), .B1(n40123), .Y(
        n18787) );
  AOI2BB2XL U43067 ( .B0(net264742), .B1(n48934), .A0N(n40284), .A1N(n34286),
        .Y(n48935) );
  OA22XL U43068 ( .A0(net262399), .A1(n34262), .B0(n34270), .B1(n40123), .Y(
        n18763) );
  AOI2BB2XL U43069 ( .B0(net265245), .B1(n48938), .A0N(n40284), .A1N(n34278),
        .Y(n48939) );
  OA22XL U43070 ( .A0(net262399), .A1(n34254), .B0(n34262), .B1(n40122), .Y(
        n18739) );
  AOI2BB2XL U43071 ( .B0(net264742), .B1(n48942), .A0N(n40284), .A1N(n34270),
        .Y(n48943) );
  OA22XL U43072 ( .A0(net262418), .A1(n34246), .B0(n34254), .B1(n40122), .Y(
        n18715) );
  AOI2BB2XL U43073 ( .B0(net264742), .B1(n48946), .A0N(n40284), .A1N(n34262),
        .Y(n48947) );
  OA22XL U43074 ( .A0(net262418), .A1(n34238), .B0(n34246), .B1(n40121), .Y(
        n18691) );
  AOI2BB2XL U43075 ( .B0(net264742), .B1(n48950), .A0N(n40285), .A1N(n34254),
        .Y(n48951) );
  OA22XL U43076 ( .A0(net262437), .A1(n34230), .B0(n34238), .B1(n40121), .Y(
        n18667) );
  AOI2BB2XL U43077 ( .B0(net264742), .B1(n48954), .A0N(n40285), .A1N(n34246),
        .Y(n48955) );
  OA22XL U43078 ( .A0(net262437), .A1(n34222), .B0(n34230), .B1(n40120), .Y(
        n18643) );
  AOI2BB2XL U43079 ( .B0(net264742), .B1(n48958), .A0N(n40285), .A1N(n34238),
        .Y(n48959) );
  OA22XL U43080 ( .A0(net262437), .A1(n34214), .B0(n34222), .B1(n40120), .Y(
        n18619) );
  AOI2BB2XL U43081 ( .B0(net264577), .B1(n48962), .A0N(n40285), .A1N(n34230),
        .Y(n48963) );
  OA22XL U43082 ( .A0(net262456), .A1(n34206), .B0(n34214), .B1(n40127), .Y(
        n18595) );
  AOI2BB2XL U43083 ( .B0(net264607), .B1(n48966), .A0N(n40285), .A1N(n34222),
        .Y(n48967) );
  OA22XL U43084 ( .A0(net262456), .A1(n34198), .B0(n34206), .B1(n40042), .Y(
        n18571) );
  AOI2BB2XL U43085 ( .B0(net264652), .B1(n48970), .A0N(n40285), .A1N(n34214),
        .Y(n48971) );
  OA22XL U43086 ( .A0(net262475), .A1(n34190), .B0(n34198), .B1(n40119), .Y(
        n18547) );
  AOI2BB2XL U43087 ( .B0(net264652), .B1(n48974), .A0N(n40285), .A1N(n34206),
        .Y(n48975) );
  OA22XL U43088 ( .A0(net262475), .A1(n34182), .B0(n34190), .B1(n40119), .Y(
        n18523) );
  AOI2BB2XL U43089 ( .B0(net264607), .B1(n48978), .A0N(n40285), .A1N(n34198),
        .Y(n48979) );
  OA22XL U43090 ( .A0(net263387), .A1(n34174), .B0(n34182), .B1(n40058), .Y(
        n18499) );
  AOI2BB2XL U43091 ( .B0(net264652), .B1(n48982), .A0N(n40285), .A1N(n34190),
        .Y(n48983) );
  OA22XL U43092 ( .A0(net263843), .A1(n34166), .B0(n34174), .B1(n40049), .Y(
        n18475) );
  AOI2BB2XL U43093 ( .B0(net221892), .B1(n48986), .A0N(n40285), .A1N(n34182),
        .Y(n48987) );
  OA22XL U43094 ( .A0(net262513), .A1(n34158), .B0(n34166), .B1(n40118), .Y(
        n18451) );
  AOI2BB2XL U43095 ( .B0(net221892), .B1(n48990), .A0N(n40285), .A1N(n34174),
        .Y(n48991) );
  OA22XL U43096 ( .A0(net262513), .A1(n34150), .B0(n34158), .B1(n40118), .Y(
        n18427) );
  AOI2BB2XL U43097 ( .B0(net264607), .B1(n48994), .A0N(n40285), .A1N(n34166),
        .Y(n48995) );
  OA22XL U43098 ( .A0(net262798), .A1(n41804), .B0(n34150), .B1(n40106), .Y(
        n18403) );
  AOI2BB2XL U43099 ( .B0(net264577), .B1(n48998), .A0N(n40285), .A1N(n34158),
        .Y(n48999) );
  OA22XL U43100 ( .A0(net262798), .A1(n41805), .B0(n41804), .B1(n40106), .Y(
        n18379) );
  AOI2BB2XL U43101 ( .B0(net221892), .B1(n49002), .A0N(n40285), .A1N(n34150),
        .Y(n49003) );
  OA22XL U43102 ( .A0(net262817), .A1(n34126), .B0(n41805), .B1(n40105), .Y(
        n18355) );
  AOI2BB2XL U43103 ( .B0(net264592), .B1(n49006), .A0N(n40285), .A1N(n41804),
        .Y(n49007) );
  OA22XL U43104 ( .A0(net262817), .A1(n34118), .B0(n34126), .B1(n40105), .Y(
        n18331) );
  NAND2XL U43105 ( .A(n42992), .B(n49515), .Y(n49012) );
  AOI2BB2XL U43106 ( .B0(net264577), .B1(n49010), .A0N(n40285), .A1N(n41805),
        .Y(n49011) );
  OA22XL U43107 ( .A0(net262817), .A1(n34110), .B0(n34118), .B1(n40076), .Y(
        n18307) );
  AOI2BB2XL U43108 ( .B0(net264846), .B1(n49078), .A0N(n40278), .A1N(n34304),
        .Y(n49079) );
  OA22XL U43109 ( .A0(net262646), .A1(n34280), .B0(n34288), .B1(n40112), .Y(
        n18817) );
  AOI2BB2XL U43110 ( .B0(net264903), .B1(n49090), .A0N(n40278), .A1N(n34280),
        .Y(n49091) );
  OA22XL U43111 ( .A0(net262399), .A1(n34256), .B0(n34264), .B1(n40122), .Y(
        n18745) );
  AOI2BB2XL U43112 ( .B0(net264903), .B1(n49094), .A0N(n40278), .A1N(n34272),
        .Y(n49095) );
  OA22XL U43113 ( .A0(net262418), .A1(n34248), .B0(n34256), .B1(n40122), .Y(
        n18721) );
  AOI2BB2XL U43114 ( .B0(net264846), .B1(n49106), .A0N(n40278), .A1N(n34248),
        .Y(n49107) );
  OA22XL U43115 ( .A0(net262437), .A1(n34224), .B0(n34232), .B1(n40120), .Y(
        n18649) );
  AOI2BB2XL U43116 ( .B0(net264682), .B1(n49110), .A0N(n40278), .A1N(n34240),
        .Y(n49111) );
  OA22XL U43117 ( .A0(net262437), .A1(n34216), .B0(n34224), .B1(n40120), .Y(
        n18625) );
  AOI2BB2XL U43118 ( .B0(net221720), .B1(n49114), .A0N(n40278), .A1N(n34232),
        .Y(n49115) );
  OA22XL U43119 ( .A0(net262456), .A1(n34208), .B0(n34216), .B1(n40053), .Y(
        n18601) );
  AOI2BB2XL U43120 ( .B0(net221720), .B1(n49118), .A0N(n40278), .A1N(n34224),
        .Y(n49119) );
  OA22XL U43121 ( .A0(net262456), .A1(n34200), .B0(n34208), .B1(n40054), .Y(
        n18577) );
  AOI2BB2XL U43122 ( .B0(net264682), .B1(n49122), .A0N(n40278), .A1N(n34216),
        .Y(n49123) );
  OA22XL U43123 ( .A0(net262475), .A1(n34192), .B0(n34200), .B1(n40119), .Y(
        n18553) );
  AOI2BB2XL U43124 ( .B0(net264682), .B1(n49126), .A0N(n40278), .A1N(n34208),
        .Y(n49127) );
  OA22XL U43125 ( .A0(net262475), .A1(n34184), .B0(n34192), .B1(n40119), .Y(
        n18529) );
  AOI2BB2XL U43126 ( .B0(net221736), .B1(n49130), .A0N(n40278), .A1N(n34200),
        .Y(n49131) );
  OA22XL U43127 ( .A0(net263843), .A1(n34176), .B0(n34184), .B1(n40070), .Y(
        n18505) );
  AOI2BB2XL U43128 ( .B0(net221736), .B1(n41231), .A0N(n40278), .A1N(n34192),
        .Y(n49134) );
  OA22XL U43129 ( .A0(net262798), .A1(n34168), .B0(n34176), .B1(n40050), .Y(
        n18481) );
  AOI2BB2XL U43130 ( .B0(net221720), .B1(n49137), .A0N(n40278), .A1N(n34184),
        .Y(n49138) );
  OA22XL U43131 ( .A0(net262798), .A1(n34160), .B0(n34168), .B1(n40118), .Y(
        n18457) );
  AOI2BB2XL U43132 ( .B0(net264682), .B1(n49141), .A0N(net217202), .A1N(n34176), .Y(n49142) );
  OA22XL U43133 ( .A0(net262513), .A1(n34152), .B0(n34160), .B1(n40118), .Y(
        n18433) );
  AOI2BB2XL U43134 ( .B0(net221720), .B1(n41259), .A0N(n40278), .A1N(n34168),
        .Y(n49145) );
  OA22XL U43135 ( .A0(net262513), .A1(n34144), .B0(n34152), .B1(n40092), .Y(
        n18409) );
  AOI2BB2XL U43136 ( .B0(net221720), .B1(n49148), .A0N(n40278), .A1N(n34160),
        .Y(n49149) );
  OA22XL U43137 ( .A0(net262798), .A1(n42058), .B0(n34144), .B1(n40106), .Y(
        n18385) );
  AOI2BB2XL U43138 ( .B0(net264682), .B1(n49152), .A0N(net217196), .A1N(n34152), .Y(n49153) );
  OA22XL U43139 ( .A0(net262798), .A1(n34128), .B0(n42058), .B1(n40105), .Y(
        n18361) );
  AOI2BB2XL U43140 ( .B0(net264682), .B1(n49156), .A0N(net217276), .A1N(n34144), .Y(n49157) );
  OA22XL U43141 ( .A0(net262817), .A1(n34120), .B0(n34128), .B1(n40105), .Y(
        n18337) );
  AOI2BB2XL U43142 ( .B0(net221720), .B1(n49160), .A0N(n40306), .A1N(n42058),
        .Y(n49161) );
  OA22XL U43143 ( .A0(net262817), .A1(n34112), .B0(n34120), .B1(n40080), .Y(
        n18313) );
  NAND2XL U43144 ( .A(n43006), .B(n49513), .Y(n49166) );
  AOI2BB2XL U43145 ( .B0(net264577), .B1(n49164), .A0N(n40306), .A1N(n34128),
        .Y(n49165) );
  OA22XL U43146 ( .A0(net262836), .A1(n34104), .B0(n34112), .B1(n40081), .Y(
        n18289) );
  AOI2BB2XL U43147 ( .B0(net264577), .B1(n49171), .A0N(n40306), .A1N(n34112),
        .Y(n49172) );
  OA22XL U43148 ( .A0(net262855), .A1(n34088), .B0(n34096), .B1(n40104), .Y(
        n18241) );
  AOI2BB2XL U43149 ( .B0(net264577), .B1(n49185), .A0N(net217188), .A1N(n34401), .Y(n49186) );
  OA22XL U43150 ( .A0(net262551), .A1(n34377), .B0(n34385), .B1(n40048), .Y(
        n19108) );
  AOI2BB2XL U43151 ( .B0(net264577), .B1(n49196), .A0N(n40289), .A1N(n34377),
        .Y(n49197) );
  OA22XL U43152 ( .A0(net262570), .A1(n34353), .B0(n34361), .B1(n40116), .Y(
        n19036) );
  AOI2BB2XL U43153 ( .B0(net264577), .B1(n49200), .A0N(n40287), .A1N(n34369),
        .Y(n49201) );
  OA22XL U43154 ( .A0(net262570), .A1(n34345), .B0(n34353), .B1(n40116), .Y(
        n19012) );
  AOI2BB2XL U43155 ( .B0(net264577), .B1(n49204), .A0N(n40287), .A1N(n34361),
        .Y(n49205) );
  OA22XL U43156 ( .A0(net262589), .A1(n34337), .B0(n34345), .B1(n40115), .Y(
        n18988) );
  AOI2BB2XL U43157 ( .B0(net264577), .B1(n49208), .A0N(n40289), .A1N(n34353),
        .Y(n49209) );
  OA22XL U43158 ( .A0(net262589), .A1(n34329), .B0(n34337), .B1(n40115), .Y(
        n18964) );
  AOI2BB2XL U43159 ( .B0(net264577), .B1(n49212), .A0N(net217182), .A1N(n34345), .Y(n49213) );
  OA22XL U43160 ( .A0(net262608), .A1(n34321), .B0(n34329), .B1(n40114), .Y(
        n18940) );
  AOI2BB2XL U43161 ( .B0(net264577), .B1(n49216), .A0N(n40306), .A1N(n34337),
        .Y(n49217) );
  OA22XL U43162 ( .A0(net262608), .A1(n34313), .B0(n34321), .B1(n40114), .Y(
        n18916) );
  AOI2BB2XL U43163 ( .B0(net264577), .B1(n49220), .A0N(net217206), .A1N(n34329), .Y(n49221) );
  OA22XL U43164 ( .A0(net262627), .A1(n34305), .B0(n34313), .B1(n40113), .Y(
        n18892) );
  AOI2BB2XL U43165 ( .B0(net264592), .B1(n49224), .A0N(net217178), .A1N(n34321), .Y(n49225) );
  OA22XL U43166 ( .A0(net262627), .A1(n34297), .B0(n34305), .B1(n40113), .Y(
        n18868) );
  AOI2BB2XL U43167 ( .B0(net264592), .B1(n49228), .A0N(net217188), .A1N(n34313), .Y(n49229) );
  OA22XL U43168 ( .A0(net262627), .A1(n34289), .B0(n34297), .B1(n40112), .Y(
        n18844) );
  AOI2BB2XL U43169 ( .B0(net264592), .B1(n49232), .A0N(net217178), .A1N(n34305), .Y(n49233) );
  OA22XL U43170 ( .A0(net262646), .A1(n34281), .B0(n34289), .B1(n40112), .Y(
        n18820) );
  AOI2BB2XL U43171 ( .B0(net264592), .B1(n49236), .A0N(net217182), .A1N(n34297), .Y(n49237) );
  OA22XL U43172 ( .A0(net262646), .A1(n34273), .B0(n34281), .B1(n40095), .Y(
        n18796) );
  AOI2BB2XL U43173 ( .B0(net264592), .B1(n49240), .A0N(net217178), .A1N(n34289), .Y(n49241) );
  OA22XL U43174 ( .A0(net262399), .A1(n34265), .B0(n34273), .B1(n40123), .Y(
        n18772) );
  AOI2BB2XL U43175 ( .B0(net264592), .B1(n49244), .A0N(net217178), .A1N(n34281), .Y(n49245) );
  OA22XL U43176 ( .A0(net262399), .A1(n34257), .B0(n34265), .B1(n40122), .Y(
        n18748) );
  AOI2BB2XL U43177 ( .B0(net264592), .B1(n49248), .A0N(net217178), .A1N(n34273), .Y(n49249) );
  OA22XL U43178 ( .A0(net262399), .A1(n34249), .B0(n34257), .B1(n40122), .Y(
        n18724) );
  AOI2BB2XL U43179 ( .B0(net264592), .B1(n49252), .A0N(net217178), .A1N(n34265), .Y(n49253) );
  OA22XL U43180 ( .A0(net262418), .A1(n34241), .B0(n34249), .B1(n40121), .Y(
        n18700) );
  AOI2BB2XL U43181 ( .B0(net264592), .B1(n49256), .A0N(net217178), .A1N(n34257), .Y(n49257) );
  OA22XL U43182 ( .A0(net262418), .A1(n34233), .B0(n34241), .B1(n40121), .Y(
        n18676) );
  AOI2BB2XL U43183 ( .B0(net264592), .B1(n49260), .A0N(net217272), .A1N(n34249), .Y(n49261) );
  OA22XL U43184 ( .A0(net262437), .A1(n34225), .B0(n34233), .B1(n40120), .Y(
        n18652) );
  AOI2BB2XL U43185 ( .B0(net264592), .B1(n49264), .A0N(net217190), .A1N(n34241), .Y(n49265) );
  OA22XL U43186 ( .A0(net262437), .A1(n34217), .B0(n34225), .B1(n40120), .Y(
        n18628) );
  AOI2BB2XL U43187 ( .B0(net264592), .B1(n49268), .A0N(net217178), .A1N(n34233), .Y(n49269) );
  OA22XL U43188 ( .A0(net262456), .A1(n34209), .B0(n34217), .B1(n40127), .Y(
        n18604) );
  AOI2BB2XL U43189 ( .B0(net264592), .B1(n49272), .A0N(net217196), .A1N(n34225), .Y(n49273) );
  OA22XL U43190 ( .A0(net262456), .A1(n34201), .B0(n34209), .B1(n40056), .Y(
        n18580) );
  AOI2BB2XL U43191 ( .B0(net264607), .B1(n49276), .A0N(net217272), .A1N(n34217), .Y(n49277) );
  OA22XL U43192 ( .A0(net262475), .A1(n34193), .B0(n34201), .B1(n40119), .Y(
        n18556) );
  AOI2BB2XL U43193 ( .B0(net264607), .B1(n49280), .A0N(net217206), .A1N(n34209), .Y(n49281) );
  OA22XL U43194 ( .A0(net262475), .A1(n34185), .B0(n34193), .B1(n40119), .Y(
        n18532) );
  AOI2BB2XL U43195 ( .B0(net264607), .B1(n49284), .A0N(net217196), .A1N(n34201), .Y(n49285) );
  OA22XL U43196 ( .A0(net262798), .A1(n34177), .B0(n34185), .B1(n40092), .Y(
        n18508) );
  AOI2BB2XL U43197 ( .B0(net264607), .B1(n49288), .A0N(net217190), .A1N(n34193), .Y(n49289) );
  OA22XL U43198 ( .A0(net263406), .A1(n34169), .B0(n34177), .B1(n40092), .Y(
        n18484) );
  AOI2BB2XL U43199 ( .B0(net264607), .B1(n41227), .A0N(n40279), .A1N(n34185),
        .Y(n49292) );
  OA22XL U43200 ( .A0(net262703), .A1(n34161), .B0(n34169), .B1(n40118), .Y(
        n18460) );
  AOI2BB2XL U43201 ( .B0(net264607), .B1(n49295), .A0N(n40279), .A1N(n34177),
        .Y(n49296) );
  OA22XL U43202 ( .A0(net262513), .A1(n34153), .B0(n34161), .B1(n40118), .Y(
        n18436) );
  AOI2BB2XL U43203 ( .B0(net264607), .B1(n49299), .A0N(n40279), .A1N(n34169),
        .Y(n49300) );
  OA22XL U43204 ( .A0(net262513), .A1(n34145), .B0(n34153), .B1(n40085), .Y(
        n18412) );
  AOI2BB2XL U43205 ( .B0(net264607), .B1(n49303), .A0N(n40279), .A1N(n34161),
        .Y(n49304) );
  OA22XL U43206 ( .A0(net262798), .A1(n42060), .B0(n34145), .B1(n40106), .Y(
        n18388) );
  AOI2BB2XL U43207 ( .B0(net264607), .B1(n49307), .A0N(n40279), .A1N(n34153),
        .Y(n49308) );
  OA22XL U43208 ( .A0(net262798), .A1(n42061), .B0(n42060), .B1(n40105), .Y(
        n18364) );
  AOI2BB2XL U43209 ( .B0(net264607), .B1(n49311), .A0N(n40279), .A1N(n34145),
        .Y(n49312) );
  OA22XL U43210 ( .A0(net262817), .A1(n34121), .B0(n42061), .B1(n40105), .Y(
        n18340) );
  AOI2BB2XL U43211 ( .B0(net264607), .B1(n49315), .A0N(n40279), .A1N(n42060),
        .Y(n49316) );
  OA22XL U43212 ( .A0(net262817), .A1(n34113), .B0(n34121), .B1(n40129), .Y(
        n18316) );
  NAND2XL U43213 ( .A(n43003), .B(n49512), .Y(n49321) );
  AOI2BB2XL U43214 ( .B0(net264607), .B1(n49319), .A0N(n40279), .A1N(n42061),
        .Y(n49320) );
  OA22XL U43215 ( .A0(net262836), .A1(n34105), .B0(n34113), .B1(n40075), .Y(
        n18292) );
  AOI2BB2XL U43216 ( .B0(net221892), .B1(n49340), .A0N(n40279), .A1N(n34402),
        .Y(n49341) );
  OA22XL U43217 ( .A0(net262532), .A1(n34378), .B0(n34386), .B1(n40086), .Y(
        n19111) );
  AOI2BB2XL U43218 ( .B0(net221892), .B1(n49351), .A0N(n40279), .A1N(n34378),
        .Y(n49352) );
  OA22XL U43219 ( .A0(net262570), .A1(n34354), .B0(n34362), .B1(n40117), .Y(
        n19039) );
  AOI2BB2XL U43220 ( .B0(net221892), .B1(n49355), .A0N(n40279), .A1N(n34370),
        .Y(n49356) );
  OA22XL U43221 ( .A0(net262570), .A1(n34346), .B0(n34354), .B1(n40116), .Y(
        n19015) );
  AOI2BB2XL U43222 ( .B0(net221892), .B1(n49359), .A0N(n40279), .A1N(n34362),
        .Y(n49360) );
  OA22XL U43223 ( .A0(net262589), .A1(n34338), .B0(n34346), .B1(n40116), .Y(
        n18991) );
  AOI2BB2XL U43224 ( .B0(net265606), .B1(n49363), .A0N(n40302), .A1N(n34354),
        .Y(n49364) );
  OA22XL U43225 ( .A0(net262589), .A1(n34330), .B0(n34338), .B1(n40115), .Y(
        n18967) );
  AOI2BB2XL U43226 ( .B0(net221892), .B1(n49367), .A0N(net217196), .A1N(n34346), .Y(n49368) );
  OA22XL U43227 ( .A0(net262608), .A1(n34322), .B0(n34330), .B1(n40114), .Y(
        n18943) );
  AOI2BB2XL U43228 ( .B0(net265378), .B1(n49371), .A0N(n40310), .A1N(n34338),
        .Y(n49372) );
  OA22XL U43229 ( .A0(net262608), .A1(n34314), .B0(n34322), .B1(n40114), .Y(
        n18919) );
  AOI2BB2XL U43230 ( .B0(net221892), .B1(n49375), .A0N(net217210), .A1N(n34330), .Y(n49376) );
  OA22XL U43231 ( .A0(net262627), .A1(n34306), .B0(n34314), .B1(n40113), .Y(
        n18895) );
  AOI2BB2XL U43232 ( .B0(net221892), .B1(n49379), .A0N(n40287), .A1N(n34322),
        .Y(n49380) );
  OA22XL U43233 ( .A0(net262627), .A1(n34298), .B0(n34306), .B1(n40113), .Y(
        n18871) );
  AOI2BB2XL U43234 ( .B0(net221892), .B1(n49383), .A0N(net217210), .A1N(n34314), .Y(n49384) );
  OA22XL U43235 ( .A0(net262627), .A1(n34290), .B0(n34298), .B1(n40112), .Y(
        n18847) );
  AOI2BB2XL U43236 ( .B0(net221804), .B1(n49387), .A0N(n40309), .A1N(n34306),
        .Y(n49388) );
  OA22XL U43237 ( .A0(net262646), .A1(n34282), .B0(n34290), .B1(n40112), .Y(
        n18823) );
  AOI2BB2XL U43238 ( .B0(net221788), .B1(n49391), .A0N(n40300), .A1N(n34298),
        .Y(n49392) );
  OA22XL U43239 ( .A0(net262646), .A1(n34274), .B0(n34282), .B1(n40089), .Y(
        n18799) );
  AOI2BB2XL U43240 ( .B0(net265150), .B1(n49395), .A0N(n40292), .A1N(n34290),
        .Y(n49396) );
  OA22XL U43241 ( .A0(net262399), .A1(n34266), .B0(n34274), .B1(n40123), .Y(
        n18775) );
  AOI2BB2XL U43242 ( .B0(net265150), .B1(n49399), .A0N(n40287), .A1N(n34282),
        .Y(n49400) );
  OA22XL U43243 ( .A0(net262399), .A1(n34258), .B0(n34266), .B1(n40122), .Y(
        n18751) );
  AOI2BB2XL U43244 ( .B0(net221788), .B1(n49403), .A0N(n40287), .A1N(n34274),
        .Y(n49404) );
  OA22XL U43245 ( .A0(net262399), .A1(n34250), .B0(n34258), .B1(n40122), .Y(
        n18727) );
  AOI2BB2XL U43246 ( .B0(net265150), .B1(n49407), .A0N(n40298), .A1N(n34266),
        .Y(n49408) );
  OA22XL U43247 ( .A0(net262418), .A1(n34242), .B0(n34250), .B1(n40121), .Y(
        n18703) );
  AOI2BB2XL U43248 ( .B0(net221788), .B1(n49411), .A0N(n40303), .A1N(n34258),
        .Y(n49412) );
  OA22XL U43249 ( .A0(net262418), .A1(n34234), .B0(n34242), .B1(n40121), .Y(
        n18679) );
  AOI2BB2XL U43250 ( .B0(net221788), .B1(n49415), .A0N(n40287), .A1N(n34250),
        .Y(n49416) );
  OA22XL U43251 ( .A0(net262437), .A1(n34226), .B0(n34234), .B1(n40120), .Y(
        n18655) );
  AOI2BB2XL U43252 ( .B0(net265150), .B1(n49419), .A0N(n40292), .A1N(n34242),
        .Y(n49420) );
  OA22XL U43253 ( .A0(net262437), .A1(n34218), .B0(n34226), .B1(n40120), .Y(
        n18631) );
  AOI2BB2XL U43254 ( .B0(net221788), .B1(n49423), .A0N(n40292), .A1N(n34234),
        .Y(n49424) );
  OA22XL U43255 ( .A0(net262456), .A1(n34210), .B0(n34218), .B1(n40040), .Y(
        n18607) );
  AOI2BB2XL U43256 ( .B0(net265150), .B1(n41221), .A0N(n40287), .A1N(n34226),
        .Y(n49427) );
  OA22XL U43257 ( .A0(net262456), .A1(n34202), .B0(n34210), .B1(n40046), .Y(
        n18583) );
  AOI2BB2XL U43258 ( .B0(net265150), .B1(n49430), .A0N(n40296), .A1N(n34218),
        .Y(n49431) );
  OA22XL U43259 ( .A0(net262475), .A1(n34194), .B0(n34202), .B1(n40119), .Y(
        n18559) );
  AOI2BB2XL U43260 ( .B0(net221788), .B1(n49434), .A0N(n40287), .A1N(n34210),
        .Y(n49435) );
  OA22XL U43261 ( .A0(net262475), .A1(n34186), .B0(n34194), .B1(n40119), .Y(
        n18535) );
  AOI2BB2XL U43262 ( .B0(net265150), .B1(n49438), .A0N(n40314), .A1N(n34202),
        .Y(n49439) );
  OA22XL U43263 ( .A0(net262475), .A1(n34178), .B0(n34186), .B1(n40058), .Y(
        n18511) );
  AOI2BB2XL U43264 ( .B0(net221788), .B1(n49442), .A0N(n40289), .A1N(n34194),
        .Y(n49443) );
  OA22XL U43265 ( .A0(net263634), .A1(n34170), .B0(n34178), .B1(n40092), .Y(
        n18487) );
  AOI2BB2XL U43266 ( .B0(net264652), .B1(n49446), .A0N(net217212), .A1N(n34186), .Y(n49447) );
  OA22XL U43267 ( .A0(net262722), .A1(n34162), .B0(n34170), .B1(n40118), .Y(
        n18463) );
  AOI2BB2XL U43268 ( .B0(net264652), .B1(n49450), .A0N(n40314), .A1N(n34178),
        .Y(n49451) );
  OA22XL U43269 ( .A0(net262513), .A1(n34154), .B0(n34162), .B1(n40118), .Y(
        n18439) );
  AOI2BB2XL U43270 ( .B0(net264652), .B1(n49454), .A0N(net217196), .A1N(n34170), .Y(n49455) );
  OA22XL U43271 ( .A0(net262513), .A1(n34146), .B0(n34154), .B1(n40084), .Y(
        n18415) );
  AOI2BB2XL U43272 ( .B0(net264652), .B1(n49458), .A0N(n40314), .A1N(n34162),
        .Y(n49459) );
  OA22XL U43273 ( .A0(net262798), .A1(n34138), .B0(n34146), .B1(n40106), .Y(
        n18391) );
  AOI2BB2XL U43274 ( .B0(net264652), .B1(n49462), .A0N(net217212), .A1N(n34154), .Y(n49463) );
  OA22XL U43275 ( .A0(net262798), .A1(n42063), .B0(n34138), .B1(n40105), .Y(
        n18367) );
  AOI2BB2XL U43276 ( .B0(net264652), .B1(n49466), .A0N(n40314), .A1N(n34146),
        .Y(n49467) );
  OA22XL U43277 ( .A0(net262817), .A1(n34122), .B0(n42063), .B1(n40105), .Y(
        n18343) );
  AOI2BB2XL U43278 ( .B0(net264652), .B1(n49470), .A0N(n40314), .A1N(n34138),
        .Y(n49471) );
  OA22XL U43279 ( .A0(net262817), .A1(n34114), .B0(n34122), .B1(n40076), .Y(
        n18319) );
  NAND2XL U43280 ( .A(n43000), .B(n49510), .Y(n49476) );
  AOI2BB2XL U43281 ( .B0(net264652), .B1(n49474), .A0N(net217196), .A1N(n42063), .Y(n49475) );
  OA22XL U43282 ( .A0(net262836), .A1(n34106), .B0(n34114), .B1(n40143), .Y(
        n18295) );
  AOI2BB2XL U43283 ( .B0(net264652), .B1(n49478), .A0N(n40314), .A1N(n34122),
        .Y(n49479) );
  OA22XL U43284 ( .A0(net262836), .A1(n34098), .B0(n34106), .B1(n40104), .Y(
        n18271) );
  AOI2BB2XL U43285 ( .B0(net264903), .B1(n49074), .A0N(n40287), .A1N(n34312),
        .Y(n49075) );
  OA22XL U43286 ( .A0(net262646), .A1(n34288), .B0(n34296), .B1(n40112), .Y(
        n18841) );
  NAND2XL U43287 ( .A(n43009), .B(n49039), .Y(n49031) );
  AOI2BB2XL U43288 ( .B0(net264532), .B1(n49029), .A0N(n40291), .A1N(n34408),
        .Y(n49030) );
  OA22XL U43289 ( .A0(net262532), .A1(n34384), .B0(n34392), .B1(n40077), .Y(
        n19129) );
  AOI2BB2XL U43290 ( .B0(net221730), .B1(n37546), .A0N(n40283), .A1N(n34117),
        .Y(n48861) );
  OA22XL U43291 ( .A0(net262836), .A1(n34093), .B0(n34101), .B1(n40104), .Y(
        n18256) );
  AOI2BB2XL U43292 ( .B0(net264652), .B1(n48557), .A0N(net217186), .A1N(n41798), .Y(n48558) );
  OA22XL U43293 ( .A0(net262532), .A1(n34388), .B0(n34396), .B1(n40086), .Y(
        n19141) );
  AOI2BB2XL U43294 ( .B0(net264652), .B1(n37554), .A0N(net217212), .A1N(n34396), .Y(n48565) );
  OA22XL U43295 ( .A0(net262551), .A1(n34372), .B0(n34380), .B1(n40079), .Y(
        n19093) );
  AOI2BB2XL U43296 ( .B0(net265492), .B1(n37544), .A0N(n40281), .A1N(n34116),
        .Y(n48702) );
  OA22XL U43297 ( .A0(net262836), .A1(n34092), .B0(n34100), .B1(n40104), .Y(
        n18253) );
  AOI2BB2XL U43298 ( .B0(net265112), .B1(n48716), .A0N(n40281), .A1N(n41800),
        .Y(n48717) );
  OA22XL U43299 ( .A0(net262532), .A1(n34389), .B0(n34397), .B1(n40071), .Y(
        n19144) );
  AOI2BB2XL U43300 ( .B0(net265416), .B1(n37549), .A0N(n40281), .A1N(n34397),
        .Y(n48723) );
  OA22XL U43301 ( .A0(net262551), .A1(n34373), .B0(n34381), .B1(n40070), .Y(
        n19096) );
  NAND2XL U43302 ( .A(n42995), .B(n49516), .Y(n48859) );
  AOI2BB2XL U43303 ( .B0(net265796), .B1(n37545), .A0N(n40283), .A1N(n34125),
        .Y(n48858) );
  OA22XL U43304 ( .A0(net262836), .A1(n34101), .B0(n34109), .B1(n40074), .Y(
        n18280) );
  AOI2BB2XL U43305 ( .B0(net265625), .B1(n48874), .A0N(n40283), .A1N(n41803),
        .Y(n48875) );
  OA22XL U43306 ( .A0(net262532), .A1(n34390), .B0(n34398), .B1(n40070), .Y(
        n19147) );
  AOI2BB2XL U43307 ( .B0(net265777), .B1(n37550), .A0N(n40284), .A1N(n34398),
        .Y(n48881) );
  OA22XL U43308 ( .A0(net262551), .A1(n34374), .B0(n34382), .B1(n40086), .Y(
        n19099) );
  NAND2XL U43309 ( .A(n42992), .B(n49514), .Y(n49015) );
  AOI2BB2XL U43310 ( .B0(net264592), .B1(n37547), .A0N(n40285), .A1N(n34126),
        .Y(n49014) );
  OA22XL U43311 ( .A0(net262836), .A1(n34102), .B0(n34110), .B1(n40080), .Y(
        n18283) );
  AOI2BB2XL U43312 ( .B0(net264592), .B1(n37548), .A0N(n40285), .A1N(n34118),
        .Y(n49017) );
  OA22XL U43313 ( .A0(net262836), .A1(n34094), .B0(n34102), .B1(n40104), .Y(
        n18259) );
  AOI2BB2XL U43314 ( .B0(net264577), .B1(n37541), .A0N(n40289), .A1N(n34120),
        .Y(n49168) );
  OA22XL U43315 ( .A0(net262836), .A1(n34096), .B0(n34104), .B1(n40104), .Y(
        n18265) );
  AOI2BB2XL U43316 ( .B0(net264577), .B1(n49181), .A0N(n40289), .A1N(n42059),
        .Y(n49182) );
  OA22XL U43317 ( .A0(net262532), .A1(n34385), .B0(n34393), .B1(n40077), .Y(
        n19132) );
  AOI2BB2XL U43318 ( .B0(net264577), .B1(n37552), .A0N(n40306), .A1N(n34393),
        .Y(n49189) );
  OA22XL U43319 ( .A0(net262551), .A1(n34369), .B0(n34377), .B1(n40117), .Y(
        n19084) );
  NAND2XL U43320 ( .A(n43003), .B(n49511), .Y(n49324) );
  AOI2BB2XL U43321 ( .B0(net264607), .B1(n37542), .A0N(n40279), .A1N(n34121),
        .Y(n49323) );
  OA22XL U43322 ( .A0(net262836), .A1(n34097), .B0(n34105), .B1(n40104), .Y(
        n18268) );
  AOI2BB2XL U43323 ( .B0(net264607), .B1(n37543), .A0N(n40279), .A1N(n34113),
        .Y(n49327) );
  OA22XL U43324 ( .A0(net262855), .A1(n34089), .B0(n34097), .B1(n40104), .Y(
        n18244) );
  AOI2BB2XL U43325 ( .B0(net221892), .B1(n49336), .A0N(n40279), .A1N(n42062),
        .Y(n49337) );
  OA22XL U43326 ( .A0(net262532), .A1(n34386), .B0(n34394), .B1(net218866),
        .Y(n19135) );
  AOI2BB2XL U43327 ( .B0(net221892), .B1(n37553), .A0N(n40279), .A1N(n34394),
        .Y(n49344) );
  OA22XL U43328 ( .A0(net262551), .A1(n34370), .B0(n34378), .B1(n40093), .Y(
        n19087) );
  AOI2BB2XL U43329 ( .B0(net264532), .B1(n37195), .A0N(n40314), .A1N(n34114),
        .Y(n49482) );
  OA22XL U43330 ( .A0(net262855), .A1(n34090), .B0(n34098), .B1(n40104), .Y(
        n18247) );
  NAND2XL U43331 ( .A(n43009), .B(n41234), .Y(n49027) );
  AOI2BB2XL U43332 ( .B0(net264532), .B1(n49025), .A0N(n40300), .A1N(n42057),
        .Y(n49026) );
  OA22XL U43333 ( .A0(net262532), .A1(n34392), .B0(n34400), .B1(n40090), .Y(
        n19153) );
  NAND2XL U43334 ( .A(n43009), .B(n49043), .Y(n49034) );
  AOI2BB2XL U43335 ( .B0(net264532), .B1(n37551), .A0N(net217202), .A1N(n34400), .Y(n49033) );
  OA22XL U43336 ( .A0(net262551), .A1(n34376), .B0(n34384), .B1(n40062), .Y(
        n19105) );
  XNOR2XL U43337 ( .A(n32818), .B(n42568), .Y(net216311) );
  XNOR2XL U43338 ( .A(n32762), .B(n42558), .Y(net216239) );
  XNOR2XL U43339 ( .A(n36839), .B(n32730), .Y(net213473) );
  XNOR2XL U43340 ( .A(n32698), .B(n42558), .Y(net216176) );
  XNOR2XL U43341 ( .A(n32634), .B(n42563), .Y(net215070) );
  XNOR2XL U43342 ( .A(n32794), .B(n42568), .Y(net216257) );
  XNOR2XL U43343 ( .A(n32802), .B(n42558), .Y(net216266) );
  XNOR2XL U43344 ( .A(n32754), .B(n42558), .Y(net216230) );
  XNOR2XL U43345 ( .A(n32658), .B(n41630), .Y(n44613) );
  XNOR2XL U43346 ( .A(n32690), .B(n42564), .Y(net216167) );
  XNOR2XL U43347 ( .A(n32730), .B(n42558), .Y(net216203) );
  XNOR2XL U43348 ( .A(n32626), .B(n42563), .Y(net215061) );
  XNOR2XL U43349 ( .A(n32786), .B(n42558), .Y(net216248) );
  XNOR2XL U43350 ( .A(n32810), .B(n42568), .Y(net216275) );
  XNOR2XL U43351 ( .A(n32642), .B(n42563), .Y(net215079) );
  XNOR2XL U43352 ( .A(n32706), .B(n42558), .Y(net216185) );
  XNOR2XL U43353 ( .A(n32834), .B(n42563), .Y(net216284) );
  XNOR2XL U43354 ( .A(n32770), .B(n42558), .Y(net216212) );
  XNOR2XL U43355 ( .A(n32682), .B(n42558), .Y(net216158) );
  XNOR2XL U43356 ( .A(n32826), .B(n42568), .Y(net216302) );
  OAI221XL U43357 ( .A0(n32398), .A1(n9727), .B0(n9728), .B1(n50087), .C0(
        n9729), .Y(nxt_data_num[2]) );
  XNOR2XL U43358 ( .A(n32650), .B(n42563), .Y(n44366) );
  XNOR2XL U43359 ( .A(n32714), .B(n42558), .Y(n43532) );
  XNOR2XL U43360 ( .A(n32842), .B(n42568), .Y(n43505) );
  XNOR2XL U43361 ( .A(n32778), .B(n42558), .Y(n43525) );
  XNOR2XL U43362 ( .A(n32602), .B(n42564), .Y(net215043) );
  XNOR2XL U43363 ( .A(n36847), .B(n32762), .Y(net212023) );
  XNOR2XL U43364 ( .A(n36844), .B(n32690), .Y(net212079) );
  XNOR2XL U43365 ( .A(n36843), .B(n32754), .Y(net212049) );
  XNOR2XL U43366 ( .A(n36736), .B(n32842), .Y(net212145) );
  XNOR2XL U43367 ( .A(n36736), .B(n32826), .Y(net212135) );
  NAND4X1 U43368 ( .A(n46648), .B(n46647), .C(n46646), .D(n46645), .Y(n10206)
         );
  XNOR2XL U43369 ( .A(n36844), .B(n32698), .Y(n46647) );
  NAND4X1 U43370 ( .A(n45616), .B(n45615), .C(n45614), .D(n45613), .Y(n10205)
         );
  XNOR2XL U43371 ( .A(n36840), .B(n32706), .Y(n45615) );
  XNOR2XL U43372 ( .A(n36734), .B(n32770), .Y(n46670) );
  XNOR2XL U43373 ( .A(n36734), .B(n32858), .Y(net212190) );
  XNOR2XL U43374 ( .A(n36840), .B(n32778), .Y(n45601) );
  XNOR2XL U43375 ( .A(n36734), .B(n32794), .Y(n47915) );
  XNOR2XL U43376 ( .A(n36735), .B(n32786), .Y(n47910) );
  XNOR2XL U43377 ( .A(n36733), .B(n32626), .Y(n47863) );
  XOR2XL U43378 ( .A(n36768), .B(n32809), .Y(n46642) );
  XOR2XL U43379 ( .A(n32676), .B(n36824), .Y(n44620) );
  XOR2XL U43380 ( .A(n41304), .B(n32700), .Y(n46644) );
  XOR2XL U43381 ( .A(n41299), .B(n32708), .Y(n45612) );
  XOR2XL U43382 ( .A(n36740), .B(n32660), .Y(n46651) );
  XOR2XL U43383 ( .A(n32740), .B(n36827), .Y(n44621) );
  XOR2XL U43384 ( .A(n32756), .B(n36823), .Y(n43521) );
  XOR2XL U43385 ( .A(n32660), .B(n36821), .Y(n44610) );
  XOR2XL U43386 ( .A(n32809), .B(n36778), .Y(n45586) );
  XOR2XL U43387 ( .A(n32684), .B(n36829), .Y(n43545) );
  XOR2XL U43388 ( .A(n32692), .B(n36827), .Y(n43540) );
  XOR2XL U43389 ( .A(n36735), .B(n32618), .Y(n46975) );
  XOR2XL U43390 ( .A(n32753), .B(n36783), .Y(n46664) );
  XOR2XL U43391 ( .A(n41301), .B(n32692), .Y(n46658) );
  XOR2XL U43392 ( .A(n36744), .B(n32724), .Y(n46662) );
  XOR2XL U43393 ( .A(n36743), .B(n32788), .Y(n47907) );
  XOR2XL U43394 ( .A(n36767), .B(n32817), .Y(n46640) );
  XOR2XL U43395 ( .A(n36774), .B(n32801), .Y(n46641) );
  XOR2XL U43396 ( .A(n32796), .B(n36822), .Y(n43514) );
  XOR2XL U43397 ( .A(n32788), .B(n36821), .Y(n43515) );
  XOR2XL U43398 ( .A(n32828), .B(n36822), .Y(n43501) );
  XOR2XL U43399 ( .A(n32780), .B(n36830), .Y(n43522) );
  XOR2XL U43400 ( .A(n41303), .B(n32788), .Y(n45589) );
  XOR2XL U43401 ( .A(n41300), .B(n32796), .Y(n45588) );
  XOR2XL U43402 ( .A(n32745), .B(n36777), .Y(n45617) );
  XOR2XL U43403 ( .A(n41301), .B(n32652), .Y(n45553) );
  XOR2XL U43404 ( .A(n36735), .B(n32714), .Y(n46663) );
  XOR2XL U43405 ( .A(n41305), .B(n32684), .Y(n45592) );
  XOR2XL U43406 ( .A(n36740), .B(n32780), .Y(n46666) );
  XOR2XL U43407 ( .A(n32721), .B(n36783), .Y(n45606) );
  XOR2XL U43408 ( .A(n32804), .B(n36824), .Y(n43513) );
  XOR2XL U43409 ( .A(n32617), .B(n36785), .Y(n45561) );
  XOR2XL U43410 ( .A(n36747), .B(n32796), .Y(n47912) );
  XOR2XL U43411 ( .A(n32844), .B(n36831), .Y(n43502) );
  XOR2XL U43412 ( .A(n41300), .B(n32780), .Y(n45598) );
  XOR2XL U43413 ( .A(n32801), .B(n36785), .Y(n45587) );
  XOR2XL U43414 ( .A(n36765), .B(n32825), .Y(n46639) );
  XOR2XL U43415 ( .A(n32836), .B(n36822), .Y(n43507) );
  XOR2XL U43416 ( .A(n32633), .B(n36782), .Y(n45558) );
  XOR2XL U43417 ( .A(n32761), .B(n36785), .Y(n46673) );
  XOR2XL U43418 ( .A(n41302), .B(n32676), .Y(n45597) );
  XOR2XL U43419 ( .A(n36748), .B(n32668), .Y(n46652) );
  XOR2XL U43420 ( .A(n36733), .B(n32586), .Y(n46979) );
  XOR2XL U43421 ( .A(n36740), .B(n32740), .Y(n46660) );
  XOR2XL U43422 ( .A(n36770), .B(n32841), .Y(n46633) );
  XOR2XL U43423 ( .A(n32772), .B(n36822), .Y(n43527) );
  XOR2XL U43424 ( .A(n32708), .B(n36830), .Y(n43534) );
  XOR2XL U43425 ( .A(n36766), .B(n32625), .Y(n47860) );
  XOR2XL U43426 ( .A(n36736), .B(n32610), .Y(n46974) );
  XOR2XL U43427 ( .A(n32820), .B(n36830), .Y(n43500) );
  XOR2XL U43428 ( .A(n32812), .B(n36830), .Y(n43512) );
  XOR2XL U43429 ( .A(n32833), .B(n36778), .Y(n45574) );
  XOR2XL U43430 ( .A(n32769), .B(n36784), .Y(n45603) );
  XOR2XL U43431 ( .A(n32732), .B(n36824), .Y(n43528) );
  XOR2XL U43432 ( .A(n32716), .B(n36829), .Y(n43529) );
  XOR2XL U43433 ( .A(n36747), .B(n32676), .Y(n46650) );
  XOR2XL U43434 ( .A(n36772), .B(n32745), .Y(n46665) );
  XOR2XL U43435 ( .A(n36748), .B(n32684), .Y(n46659) );
  XOR2XL U43436 ( .A(n32764), .B(n36830), .Y(n43516) );
  XOR2XL U43437 ( .A(n32700), .B(n36823), .Y(n43535) );
  XOR2XL U43438 ( .A(n36743), .B(n32692), .Y(n46649) );
  XOR2XL U43439 ( .A(n32729), .B(n36776), .Y(n45604) );
  XOR2XL U43440 ( .A(n41305), .B(n32668), .Y(n45591) );
  XOR2XL U43441 ( .A(n36750), .B(n32700), .Y(n46643) );
  XOR2XL U43442 ( .A(n36773), .B(n32857), .Y(n46616) );
  XOR2XL U43443 ( .A(n36770), .B(n32633), .Y(n47865) );
  XOR2XL U43444 ( .A(n36764), .B(n32769), .Y(n46667) );
  XOR2XL U43445 ( .A(n36733), .B(n32642), .Y(n46973) );
  XNOR2XL U43446 ( .A(n32498), .B(n36845), .Y(net213216) );
  XNOR2XL U43447 ( .A(n32562), .B(n42564), .Y(net214989) );
  XNOR2XL U43448 ( .A(n36733), .B(n32650), .Y(net211619) );
  XNOR2XL U43449 ( .A(n36735), .B(n32602), .Y(net211614) );
  XNOR2XL U43450 ( .A(n32666), .B(n42558), .Y(n44618) );
  XNOR2XL U43451 ( .A(n36736), .B(n32554), .Y(net211580) );
  XNOR2XL U43452 ( .A(n32490), .B(n42563), .Y(net215124) );
  XNOR2XL U43453 ( .A(n36840), .B(n32514), .Y(net213226) );
  XNOR2XL U43454 ( .A(n36733), .B(n32410), .Y(net211188) );
  XNOR2XL U43455 ( .A(n32442), .B(n42565), .Y(n47273) );
  XNOR2XL U43456 ( .A(n36735), .B(n32466), .Y(net211439) );
  XNOR2XL U43457 ( .A(n32554), .B(n42564), .Y(net214962) );
  XNOR2XL U43458 ( .A(n36735), .B(n32474), .Y(net211444) );
  XNOR2XL U43459 ( .A(n32450), .B(n42562), .Y(n44324) );
  XNOR2XL U43460 ( .A(n36837), .B(n32522), .Y(net213211) );
  XNOR2XL U43461 ( .A(n32570), .B(n42564), .Y(net214998) );
  XNOR2XL U43462 ( .A(n36733), .B(n32522), .Y(net211469) );
  XNOR2XL U43463 ( .A(n32418), .B(n42563), .Y(n44338) );
  XNOR2XL U43464 ( .A(n32426), .B(n42563), .Y(n44343) );
  XNOR2XL U43465 ( .A(n32458), .B(n42562), .Y(n44333) );
  XNOR2XL U43466 ( .A(n32442), .B(n36847), .Y(n47870) );
  XNOR2XL U43467 ( .A(n32506), .B(n42560), .Y(net213221) );
  XNOR2XL U43468 ( .A(n32594), .B(n42564), .Y(net215052) );
  XNOR2XL U43469 ( .A(n36838), .B(n32418), .Y(net212553) );
  XNOR2XL U43470 ( .A(n36845), .B(n32426), .Y(net212558) );
  XNOR2XL U43471 ( .A(n36838), .B(n32466), .Y(net213232) );
  XNOR2XL U43472 ( .A(n36838), .B(n32570), .Y(n45545) );
  XNOR2XL U43473 ( .A(n32498), .B(n42565), .Y(net213206) );
  XNOR2XL U43474 ( .A(n32434), .B(n36841), .Y(n47278) );
  XNOR2XL U43475 ( .A(n36843), .B(n32578), .Y(n45540) );
  XNOR2XL U43476 ( .A(n32610), .B(n42564), .Y(n44388) );
  XNOR2XL U43477 ( .A(n32514), .B(n42563), .Y(net215097) );
  XNOR2XL U43478 ( .A(n32578), .B(n42564), .Y(net215016) );
  XNOR2XL U43479 ( .A(n32746), .B(n42560), .Y(net214673) );
  XNOR2XL U43480 ( .A(n36838), .B(n32482), .Y(net213196) );
  XNOR2XL U43481 ( .A(n36837), .B(n32490), .Y(net213201) );
  XNOR2XL U43482 ( .A(n32506), .B(n36844), .Y(net213191) );
  XNOR2XL U43483 ( .A(n36736), .B(n32402), .Y(net211559) );
  XNOR2XL U43484 ( .A(n36846), .B(n32714), .Y(n45610) );
  XNOR2XL U43485 ( .A(n32618), .B(n42564), .Y(n44397) );
  XNOR2XL U43486 ( .A(n36742), .B(n32460), .Y(n46988) );
  XNOR2XL U43487 ( .A(n36736), .B(n32434), .Y(n47875) );
  XNOR2XL U43488 ( .A(n32586), .B(n42564), .Y(n44403) );
  XNOR2XL U43489 ( .A(n36845), .B(n32586), .Y(n45535) );
  XNOR2XL U43490 ( .A(n36841), .B(n32458), .Y(n45713) );
  XNOR2XL U43491 ( .A(n32522), .B(n42563), .Y(n44360) );
  XOR2XL U43492 ( .A(n41301), .B(n32484), .Y(n45796) );
  XOR2XL U43493 ( .A(n41299), .B(n32412), .Y(n46307) );
  XOR2XL U43494 ( .A(n32724), .B(n36825), .Y(n44622) );
  XOR2XL U43495 ( .A(n32489), .B(n36778), .Y(n45795) );
  XOR2XL U43496 ( .A(n36750), .B(n32404), .Y(n46991) );
  XOR2XL U43497 ( .A(n32505), .B(n36783), .Y(n45797) );
  XOR2XL U43498 ( .A(n36747), .B(n32540), .Y(n46984) );
  XOR2XL U43499 ( .A(n36773), .B(n32489), .Y(n47049) );
  XOR2XL U43500 ( .A(n32553), .B(n36786), .Y(n45567) );
  XOR2XL U43501 ( .A(n41304), .B(n32532), .Y(n45565) );
  XOR2XL U43502 ( .A(n41302), .B(n32468), .Y(n45789) );
  XOR2XL U43503 ( .A(n32444), .B(n36827), .Y(n47270) );
  XOR2XL U43504 ( .A(n32508), .B(n36828), .Y(n45791) );
  XOR2XL U43505 ( .A(n32500), .B(n36821), .Y(n45794) );
  XOR2XL U43506 ( .A(n41304), .B(n32660), .Y(n45590) );
  XOR2XL U43507 ( .A(n41305), .B(n32524), .Y(n45793) );
  XOR2XL U43508 ( .A(n41300), .B(n32460), .Y(n45710) );
  XOR2XL U43509 ( .A(n36765), .B(n32505), .Y(n47047) );
  XOR2XL U43510 ( .A(n32436), .B(n41303), .Y(n47275) );
  XOR2XL U43511 ( .A(n41303), .B(n32540), .Y(n45564) );
  XOR2XL U43512 ( .A(n32436), .B(n36831), .Y(n46306) );
  XOR2XL U43513 ( .A(n36766), .B(n32593), .Y(n46978) );
  XOR2XL U43514 ( .A(n41304), .B(n32548), .Y(n45566) );
  XOR2XL U43515 ( .A(n41301), .B(n32476), .Y(n45788) );
  XOR2XL U43516 ( .A(n36746), .B(n32732), .Y(n46661) );
  XOR2XL U43517 ( .A(n32444), .B(n41303), .Y(n47867) );
  XOR2XL U43518 ( .A(n36774), .B(n32513), .Y(n47046) );
  XOR2XL U43519 ( .A(n32748), .B(n36822), .Y(n44623) );
  XOR2XL U43520 ( .A(n32668), .B(n36829), .Y(n44615) );
  XOR2XL U43521 ( .A(n36772), .B(n32601), .Y(n46977) );
  XOR2XL U43522 ( .A(n36742), .B(n32524), .Y(n47045) );
  XOR2XL U43523 ( .A(n36740), .B(n32468), .Y(n47051) );
  XOR2XL U43524 ( .A(n41302), .B(n32420), .Y(n46309) );
  XOR2XL U43525 ( .A(n41299), .B(n32452), .Y(n45715) );
  XOR2XL U43526 ( .A(n32433), .B(n36774), .Y(n47872) );
  XOR2XL U43527 ( .A(n32497), .B(n36786), .Y(n45792) );
  XOR2XL U43528 ( .A(n32585), .B(n36783), .Y(n45532) );
  XOR2XL U43529 ( .A(n32753), .B(n36766), .Y(n46674) );
  XOR2XL U43530 ( .A(n36736), .B(n32458), .Y(n46985) );
  XOR2XL U43531 ( .A(n41300), .B(n32428), .Y(n46308) );
  XOR2XL U43532 ( .A(n32425), .B(n36765), .Y(n47280) );
  XOR2XL U43533 ( .A(n41305), .B(n32404), .Y(n45716) );
  XOR2XL U43534 ( .A(n36743), .B(n32652), .Y(n46976) );
  XOR2XL U43535 ( .A(n36750), .B(n32532), .Y(n46981) );
  XOR2XL U43536 ( .A(n32737), .B(n36784), .Y(n45605) );
  XOR2XL U43537 ( .A(n36743), .B(n32476), .Y(n47050) );
  XOR2XL U43538 ( .A(n32713), .B(n36782), .Y(n45607) );
  XOR2XL U43539 ( .A(n32481), .B(n36764), .Y(n47052) );
  XOR2XL U43540 ( .A(n36767), .B(n32497), .Y(n47048) );
  XOR2XL U43541 ( .A(n32548), .B(n36824), .Y(n44422) );
  XOR2XL U43542 ( .A(n32417), .B(n36772), .Y(n47269) );
  XOR2XL U43543 ( .A(n36741), .B(n32412), .Y(n47268) );
  XOR2XL U43544 ( .A(n36771), .B(n32561), .Y(n47859) );
  XOR2XL U43545 ( .A(n32761), .B(n36770), .Y(n46672) );
  XOR2XL U43546 ( .A(n36768), .B(n32569), .Y(n47858) );
  XOR2XL U43547 ( .A(n32441), .B(n36770), .Y(n47866) );
  XOR2XL U43548 ( .A(n32609), .B(n36782), .Y(n45563) );
  XOR2XL U43549 ( .A(n36749), .B(n32708), .Y(n46653) );
  XOR2XL U43550 ( .A(n32556), .B(n36821), .Y(n44421) );
  XOR2XL U43551 ( .A(n32532), .B(n36825), .Y(n44416) );
  XOR2XL U43552 ( .A(n32513), .B(n36783), .Y(n45790) );
  XOR2XL U43553 ( .A(n36733), .B(n32578), .Y(n46980) );
  XOR2XL U43554 ( .A(n32545), .B(n36773), .Y(n46982) );
  XOR2XL U43555 ( .A(n36736), .B(n32450), .Y(n46990) );
  XOR2XL U43556 ( .A(n36767), .B(n32553), .Y(n46983) );
  NOR2X1 U43557 ( .A(n50143), .B(state[1]), .Y(n9689) );
  XNOR2XL U43558 ( .A(n32402), .B(n42562), .Y(n44318) );
  XOR2XL U43559 ( .A(n32404), .B(n36822), .Y(n44315) );
  NOR2X1 U43560 ( .A(n50148), .B(n32398), .Y(n19376) );
  AOI31XL U43561 ( .A0(n9683), .A1(n49556), .A2(state[0]), .B0(n41736), .Y(
        n9682) );
  CLKINVX1 U43562 ( .A(data[17]), .Y(n49538) );
  CLKINVX1 U43563 ( .A(data[18]), .Y(n49537) );
  CLKINVX1 U43564 ( .A(data[19]), .Y(n49536) );
  CLKINVX1 U43565 ( .A(data[20]), .Y(n49535) );
  CLKINVX1 U43566 ( .A(data[21]), .Y(n49534) );
  CLKINVX1 U43567 ( .A(data[22]), .Y(n49533) );
  CLKINVX1 U43568 ( .A(data[23]), .Y(n49532) );
  CLKINVX1 U43569 ( .A(data[1]), .Y(n49554) );
  CLKINVX1 U43570 ( .A(data[2]), .Y(n49553) );
  CLKINVX1 U43571 ( .A(data[3]), .Y(n49552) );
  CLKINVX1 U43572 ( .A(data[4]), .Y(n49551) );
  CLKINVX1 U43573 ( .A(data[5]), .Y(n49550) );
  CLKINVX1 U43574 ( .A(data[6]), .Y(n49549) );
  CLKINVX1 U43575 ( .A(data[7]), .Y(n49548) );
  CLKINVX1 U43576 ( .A(data[0]), .Y(n49555) );
  CLKINVX1 U43577 ( .A(data[16]), .Y(n49539) );
  INVXL U43578 ( .A(n34105), .Y(n49326) );
  CLKINVX1 U43579 ( .A(reset), .Y(n49523) );
  INVX16 U43580 ( .A(n41791), .Y(out_valid) );
  OR2X4 U43581 ( .A(n50149), .B(n50143), .Y(n41791) );
  INVX3 U43582 ( .A(n40175), .Y(net217944) );
  INVX3 U43583 ( .A(n40315), .Y(net217036) );
  INVX3 U43584 ( .A(net217238), .Y(net216978) );
  CLKBUFX3 U43585 ( .A(net218244), .Y(net218174) );
  CLKBUFX3 U43586 ( .A(net218244), .Y(net218176) );
  CLKBUFX3 U43587 ( .A(net218242), .Y(net218178) );
  CLKBUFX3 U43588 ( .A(net218242), .Y(net218180) );
  CLKBUFX3 U43589 ( .A(net218240), .Y(net218182) );
  CLKBUFX3 U43590 ( .A(net218240), .Y(net218184) );
  CLKBUFX3 U43591 ( .A(net218238), .Y(net218186) );
  CLKBUFX3 U43592 ( .A(net218250), .Y(net218164) );
  CLKBUFX3 U43593 ( .A(net218250), .Y(net218162) );
  CLKBUFX3 U43594 ( .A(net218248), .Y(net218166) );
  CLKBUFX3 U43595 ( .A(net218248), .Y(net218168) );
  CLKBUFX3 U43596 ( .A(net218246), .Y(net218170) );
  CLKBUFX3 U43597 ( .A(net218246), .Y(net218172) );
  CLKBUFX3 U43598 ( .A(net218230), .Y(net218204) );
  CLKBUFX3 U43599 ( .A(net218228), .Y(net218206) );
  CLKBUFX3 U43600 ( .A(net218228), .Y(net218208) );
  CLKBUFX3 U43601 ( .A(net218226), .Y(net218210) );
  CLKBUFX3 U43602 ( .A(net218226), .Y(net218212) );
  CLKBUFX3 U43603 ( .A(net218238), .Y(net218188) );
  CLKBUFX3 U43604 ( .A(net218236), .Y(net218190) );
  CLKBUFX3 U43605 ( .A(net218236), .Y(net218192) );
  CLKBUFX3 U43606 ( .A(net218234), .Y(net218194) );
  CLKBUFX3 U43607 ( .A(net218234), .Y(net218196) );
  CLKBUFX3 U43608 ( .A(net218232), .Y(net218198) );
  CLKBUFX3 U43609 ( .A(net218232), .Y(net218200) );
  CLKBUFX3 U43610 ( .A(net218230), .Y(net218202) );
  CLKINVX1 U43611 ( .A(n43033), .Y(n42735) );
  CLKBUFX3 U43612 ( .A(net217236), .Y(net217144) );
  CLKBUFX3 U43613 ( .A(net217234), .Y(net217146) );
  CLKBUFX3 U43614 ( .A(net217234), .Y(net217148) );
  CLKBUFX3 U43615 ( .A(net217232), .Y(net217150) );
  CLKBUFX3 U43616 ( .A(net217232), .Y(net217152) );
  CLKBUFX3 U43617 ( .A(net217230), .Y(net217154) );
  CLKBUFX3 U43618 ( .A(net217230), .Y(net217156) );
  CLKBUFX3 U43619 ( .A(net217228), .Y(net217158) );
  CLKBUFX3 U43620 ( .A(net217228), .Y(net217160) );
  CLKBUFX3 U43621 ( .A(net217226), .Y(net217162) );
  CLKBUFX3 U43622 ( .A(net217244), .Y(net217128) );
  CLKBUFX3 U43623 ( .A(net217244), .Y(net217126) );
  CLKBUFX3 U43624 ( .A(net217246), .Y(net217124) );
  CLKBUFX3 U43625 ( .A(net217246), .Y(net217122) );
  CLKBUFX3 U43626 ( .A(net217242), .Y(net217132) );
  CLKBUFX3 U43627 ( .A(net217240), .Y(net217134) );
  CLKBUFX3 U43628 ( .A(net217240), .Y(net217136) );
  CLKBUFX3 U43629 ( .A(net217238), .Y(net217138) );
  CLKBUFX3 U43630 ( .A(net217238), .Y(net217140) );
  CLKBUFX3 U43631 ( .A(net217236), .Y(net217142) );
  CLKBUFX3 U43632 ( .A(net217222), .Y(net217172) );
  CLKBUFX3 U43633 ( .A(net217220), .Y(net217174) );
  CLKBUFX3 U43634 ( .A(net217220), .Y(net217176) );
  CLKBUFX3 U43635 ( .A(net217222), .Y(net217170) );
  CLKBUFX3 U43636 ( .A(net217224), .Y(net217168) );
  CLKBUFX3 U43637 ( .A(net217224), .Y(net217166) );
  CLKBUFX3 U43638 ( .A(net217226), .Y(net217164) );
  CLKBUFX3 U43639 ( .A(net218224), .Y(net218214) );
  CLKBUFX3 U43640 ( .A(net218224), .Y(net218216) );
  CLKBUFX3 U43641 ( .A(net218262), .Y(net218258) );
  CLKBUFX3 U43642 ( .A(net218264), .Y(net218256) );
  CLKBUFX3 U43643 ( .A(net218264), .Y(net218254) );
  CLKBUFX3 U43644 ( .A(net218262), .Y(net218260) );
  CLKBUFX3 U43645 ( .A(net218270), .Y(net218244) );
  CLKBUFX3 U43646 ( .A(net218270), .Y(net218242) );
  CLKBUFX3 U43647 ( .A(net218272), .Y(net218240) );
  CLKBUFX3 U43648 ( .A(net218266), .Y(net218250) );
  CLKBUFX3 U43649 ( .A(net218266), .Y(net218252) );
  CLKBUFX3 U43650 ( .A(net218268), .Y(net218248) );
  CLKBUFX3 U43651 ( .A(net218268), .Y(net218246) );
  CLKBUFX3 U43652 ( .A(net218278), .Y(net218228) );
  CLKBUFX3 U43653 ( .A(net218278), .Y(net218226) );
  CLKBUFX3 U43654 ( .A(net218272), .Y(net218238) );
  CLKBUFX3 U43655 ( .A(net218274), .Y(net218236) );
  CLKBUFX3 U43656 ( .A(net218274), .Y(net218234) );
  CLKBUFX3 U43657 ( .A(net218276), .Y(net218232) );
  CLKBUFX3 U43658 ( .A(net217212), .Y(net217190) );
  CLKBUFX3 U43659 ( .A(net217214), .Y(net217188) );
  CLKBUFX3 U43660 ( .A(net217216), .Y(net217184) );
  CLKBUFX3 U43661 ( .A(net217216), .Y(net217182) );
  CLKBUFX3 U43662 ( .A(net217178), .Y(net217180) );
  CLKBUFX3 U43663 ( .A(net217214), .Y(net217186) );
  CLKBUFX3 U43664 ( .A(net217206), .Y(net217202) );
  CLKBUFX3 U43665 ( .A(net217210), .Y(net217196) );
  CLKBUFX3 U43666 ( .A(net218910), .Y(net218694) );
  CLKBUFX3 U43667 ( .A(net218910), .Y(net218696) );
  CLKBUFX3 U43668 ( .A(net218910), .Y(net218698) );
  CLKBUFX3 U43669 ( .A(net218908), .Y(net218700) );
  CLKBUFX3 U43670 ( .A(net218908), .Y(net218702) );
  CLKBUFX3 U43671 ( .A(net218908), .Y(net218704) );
  CLKBUFX3 U43672 ( .A(net218914), .Y(net218676) );
  CLKBUFX3 U43673 ( .A(net218914), .Y(net218678) );
  CLKBUFX3 U43674 ( .A(net218914), .Y(net218680) );
  CLKBUFX3 U43675 ( .A(net218912), .Y(net218684) );
  CLKBUFX3 U43676 ( .A(net218912), .Y(net218688) );
  CLKBUFX3 U43677 ( .A(net218902), .Y(net218724) );
  CLKBUFX3 U43678 ( .A(net218902), .Y(net218728) );
  CLKBUFX3 U43679 ( .A(net218902), .Y(net218730) );
  CLKBUFX3 U43680 ( .A(net218900), .Y(net218732) );
  CLKBUFX3 U43681 ( .A(net218900), .Y(net218736) );
  CLKBUFX3 U43682 ( .A(net218906), .Y(net218708) );
  CLKBUFX3 U43683 ( .A(net218906), .Y(net218710) );
  CLKBUFX3 U43684 ( .A(net218906), .Y(net218712) );
  CLKBUFX3 U43685 ( .A(net218904), .Y(net218716) );
  CLKBUFX3 U43686 ( .A(net218904), .Y(net218720) );
  CLKBUFX3 U43687 ( .A(net218904), .Y(net218722) );
  CLKBUFX3 U43688 ( .A(net218926), .Y(net218628) );
  CLKBUFX3 U43689 ( .A(net218926), .Y(net218632) );
  CLKBUFX3 U43690 ( .A(net218926), .Y(net218634) );
  CLKBUFX3 U43691 ( .A(net218924), .Y(net218636) );
  CLKBUFX3 U43692 ( .A(net218924), .Y(net218640) );
  CLKBUFX3 U43693 ( .A(net218930), .Y(net218612) );
  CLKBUFX3 U43694 ( .A(net218930), .Y(net218614) );
  CLKBUFX3 U43695 ( .A(net218930), .Y(net218616) );
  CLKBUFX3 U43696 ( .A(net218930), .Y(net218618) );
  CLKBUFX3 U43697 ( .A(net218928), .Y(net218620) );
  CLKBUFX3 U43698 ( .A(net218928), .Y(net218622) );
  CLKBUFX3 U43699 ( .A(net218928), .Y(net218624) );
  CLKBUFX3 U43700 ( .A(net218928), .Y(net218626) );
  CLKBUFX3 U43701 ( .A(net218918), .Y(net218660) );
  CLKBUFX3 U43702 ( .A(net218918), .Y(net218664) );
  CLKBUFX3 U43703 ( .A(net218918), .Y(net218666) );
  CLKBUFX3 U43704 ( .A(net218916), .Y(net218668) );
  CLKBUFX3 U43705 ( .A(net218916), .Y(net218670) );
  CLKBUFX3 U43706 ( .A(net218916), .Y(net218672) );
  CLKBUFX3 U43707 ( .A(net218916), .Y(net218674) );
  CLKBUFX3 U43708 ( .A(net218924), .Y(net218642) );
  CLKBUFX3 U43709 ( .A(net218922), .Y(net218644) );
  CLKBUFX3 U43710 ( .A(net218922), .Y(net218646) );
  CLKBUFX3 U43711 ( .A(net218922), .Y(net218648) );
  CLKBUFX3 U43712 ( .A(net218922), .Y(net218650) );
  CLKBUFX3 U43713 ( .A(net218920), .Y(net218652) );
  CLKBUFX3 U43714 ( .A(net218920), .Y(net218654) );
  CLKBUFX3 U43715 ( .A(net218920), .Y(net218656) );
  CLKBUFX3 U43716 ( .A(net218920), .Y(net218658) );
  CLKBUFX3 U43717 ( .A(net218878), .Y(net218820) );
  CLKBUFX3 U43718 ( .A(net218878), .Y(net218822) );
  CLKBUFX3 U43719 ( .A(net218878), .Y(net218824) );
  CLKBUFX3 U43720 ( .A(net218876), .Y(net218828) );
  CLKBUFX3 U43721 ( .A(net218876), .Y(net218830) );
  CLKBUFX3 U43722 ( .A(net218876), .Y(net218832) );
  CLKBUFX3 U43723 ( .A(net218882), .Y(net218804) );
  CLKBUFX3 U43724 ( .A(net218882), .Y(net218806) );
  CLKBUFX3 U43725 ( .A(net218882), .Y(net218808) );
  CLKBUFX3 U43726 ( .A(net218882), .Y(net218810) );
  CLKBUFX3 U43727 ( .A(net218880), .Y(net218812) );
  CLKBUFX3 U43728 ( .A(net218880), .Y(net218814) );
  CLKBUFX3 U43729 ( .A(net218880), .Y(net218816) );
  CLKBUFX3 U43730 ( .A(net218880), .Y(net218818) );
  CLKBUFX3 U43731 ( .A(net218870), .Y(net218852) );
  CLKBUFX3 U43732 ( .A(net218870), .Y(net218854) );
  CLKBUFX3 U43733 ( .A(net218870), .Y(net218856) );
  CLKBUFX3 U43734 ( .A(net218876), .Y(net218834) );
  CLKBUFX3 U43735 ( .A(net218874), .Y(net218836) );
  CLKBUFX3 U43736 ( .A(net218874), .Y(net218838) );
  CLKBUFX3 U43737 ( .A(net218874), .Y(net218840) );
  CLKBUFX3 U43738 ( .A(net218874), .Y(net218842) );
  CLKBUFX3 U43739 ( .A(net218872), .Y(net218844) );
  CLKBUFX3 U43740 ( .A(net218872), .Y(net218846) );
  CLKBUFX3 U43741 ( .A(net218872), .Y(net218848) );
  CLKBUFX3 U43742 ( .A(net218872), .Y(net218850) );
  CLKBUFX3 U43743 ( .A(net218894), .Y(net218756) );
  CLKBUFX3 U43744 ( .A(net218894), .Y(net218758) );
  CLKBUFX3 U43745 ( .A(net218894), .Y(net218760) );
  CLKBUFX3 U43746 ( .A(net218894), .Y(net218762) );
  CLKBUFX3 U43747 ( .A(net218892), .Y(net218764) );
  CLKBUFX3 U43748 ( .A(net218892), .Y(net218766) );
  CLKBUFX3 U43749 ( .A(net218892), .Y(net218768) );
  CLKBUFX3 U43750 ( .A(net218900), .Y(net218738) );
  CLKBUFX3 U43751 ( .A(net218898), .Y(net218740) );
  CLKBUFX3 U43752 ( .A(net218898), .Y(net218742) );
  CLKBUFX3 U43753 ( .A(net218898), .Y(net218744) );
  CLKBUFX3 U43754 ( .A(net218898), .Y(net218746) );
  CLKBUFX3 U43755 ( .A(net218896), .Y(net218748) );
  CLKBUFX3 U43756 ( .A(net218896), .Y(net218750) );
  CLKBUFX3 U43757 ( .A(net218896), .Y(net218752) );
  CLKBUFX3 U43758 ( .A(net218896), .Y(net218754) );
  CLKBUFX3 U43759 ( .A(net218888), .Y(net218786) );
  CLKBUFX3 U43760 ( .A(net218886), .Y(net218788) );
  CLKBUFX3 U43761 ( .A(net218886), .Y(net218790) );
  CLKBUFX3 U43762 ( .A(net218886), .Y(net218792) );
  CLKBUFX3 U43763 ( .A(net218886), .Y(net218794) );
  CLKBUFX3 U43764 ( .A(net218884), .Y(net218796) );
  CLKBUFX3 U43765 ( .A(net218884), .Y(net218798) );
  CLKBUFX3 U43766 ( .A(net218884), .Y(net218800) );
  CLKBUFX3 U43767 ( .A(net218884), .Y(net218802) );
  CLKBUFX3 U43768 ( .A(net218892), .Y(net218770) );
  CLKBUFX3 U43769 ( .A(net218890), .Y(net218772) );
  CLKBUFX3 U43770 ( .A(net218890), .Y(net218774) );
  CLKBUFX3 U43771 ( .A(net218890), .Y(net218776) );
  CLKBUFX3 U43772 ( .A(net218890), .Y(net218778) );
  CLKBUFX3 U43773 ( .A(net218888), .Y(net218780) );
  CLKBUFX3 U43774 ( .A(net218888), .Y(net218782) );
  CLKBUFX3 U43775 ( .A(net218868), .Y(net218860) );
  CLKBUFX3 U43776 ( .A(net218868), .Y(net218862) );
  CLKBUFX3 U43777 ( .A(net218868), .Y(net218864) );
  CLKBUFX3 U43778 ( .A(n43031), .Y(n43009) );
  CLKBUFX3 U43779 ( .A(n43025), .Y(n43021) );
  CLKBUFX3 U43780 ( .A(n43025), .Y(n43022) );
  CLKBUFX3 U43781 ( .A(n43027), .Y(n43018) );
  CLKBUFX3 U43782 ( .A(n43026), .Y(n43019) );
  CLKBUFX3 U43783 ( .A(n43026), .Y(n43020) );
  CLKBUFX3 U43784 ( .A(n43029), .Y(n43014) );
  CLKBUFX3 U43785 ( .A(n43027), .Y(n43017) );
  CLKBUFX3 U43786 ( .A(n43028), .Y(n43015) );
  CLKBUFX3 U43787 ( .A(n43028), .Y(n43016) );
  CLKBUFX3 U43788 ( .A(n43031), .Y(n43010) );
  CLKBUFX3 U43789 ( .A(n43029), .Y(n43013) );
  CLKBUFX3 U43790 ( .A(n43030), .Y(n43011) );
  CLKBUFX3 U43791 ( .A(n43030), .Y(n43012) );
  CLKBUFX3 U43792 ( .A(net218868), .Y(net218866) );
  CLKBUFX3 U43793 ( .A(net218284), .Y(net218270) );
  CLKBUFX3 U43794 ( .A(net218286), .Y(net218278) );
  CLKBUFX3 U43795 ( .A(net218284), .Y(net218272) );
  CLKBUFX3 U43796 ( .A(net218286), .Y(net218274) );
  CLKBUFX3 U43797 ( .A(net218286), .Y(net218276) );
  CLKBUFX3 U43798 ( .A(net217262), .Y(net217234) );
  CLKBUFX3 U43799 ( .A(net217264), .Y(net217232) );
  CLKBUFX3 U43800 ( .A(net217264), .Y(net217230) );
  CLKBUFX3 U43801 ( .A(net217266), .Y(net217228) );
  CLKBUFX3 U43802 ( .A(net217258), .Y(net217244) );
  CLKBUFX3 U43803 ( .A(net217260), .Y(net217240) );
  CLKBUFX3 U43804 ( .A(net218274), .Y(net218224) );
  CLKBUFX3 U43805 ( .A(net217260), .Y(net217238) );
  CLKBUFX3 U43806 ( .A(net217262), .Y(net217236) );
  CLKBUFX3 U43807 ( .A(net218274), .Y(net218222) );
  CLKBUFX3 U43808 ( .A(net217268), .Y(net217222) );
  CLKBUFX3 U43809 ( .A(net217268), .Y(net217224) );
  CLKBUFX3 U43810 ( .A(n43032), .Y(n42992) );
  CLKBUFX3 U43811 ( .A(n43032), .Y(n42999) );
  CLKBUFX3 U43812 ( .A(n43032), .Y(n42998) );
  CLKBUFX3 U43813 ( .A(n43032), .Y(n42997) );
  CLKBUFX3 U43814 ( .A(n43009), .Y(n42995) );
  CLKBUFX3 U43815 ( .A(n43032), .Y(n42994) );
  CLKBUFX3 U43816 ( .A(n43032), .Y(n42993) );
  CLKBUFX3 U43817 ( .A(n43009), .Y(n42996) );
  CLKBUFX3 U43818 ( .A(n43032), .Y(n43008) );
  CLKBUFX3 U43819 ( .A(n43032), .Y(n43007) );
  CLKBUFX3 U43820 ( .A(n43032), .Y(n43006) );
  CLKBUFX3 U43821 ( .A(n43032), .Y(n43004) );
  CLKBUFX3 U43822 ( .A(n43032), .Y(n43003) );
  CLKBUFX3 U43823 ( .A(n43032), .Y(n43005) );
  CLKBUFX3 U43824 ( .A(n43032), .Y(n43002) );
  CLKBUFX3 U43825 ( .A(n43032), .Y(n43001) );
  CLKBUFX3 U43826 ( .A(n43032), .Y(n43000) );
  CLKBUFX3 U43827 ( .A(net217272), .Y(net217216) );
  CLKBUFX3 U43828 ( .A(net217272), .Y(net217214) );
  CLKBUFX3 U43829 ( .A(net217274), .Y(net217210) );
  CLKBUFX3 U43830 ( .A(net217274), .Y(net217212) );
  CLKBUFX3 U43831 ( .A(net218934), .Y(net218932) );
  CLKBUFX3 U43832 ( .A(net218940), .Y(net218910) );
  CLKBUFX3 U43833 ( .A(net218940), .Y(net218914) );
  CLKBUFX3 U43834 ( .A(net218940), .Y(net218912) );
  CLKBUFX3 U43835 ( .A(net218944), .Y(net218902) );
  CLKBUFX3 U43836 ( .A(net218942), .Y(net218908) );
  CLKBUFX3 U43837 ( .A(net218942), .Y(net218906) );
  CLKBUFX3 U43838 ( .A(net218942), .Y(net218904) );
  CLKBUFX3 U43839 ( .A(net218936), .Y(net218926) );
  CLKBUFX3 U43840 ( .A(net218938), .Y(net218918) );
  CLKBUFX3 U43841 ( .A(net218938), .Y(net218916) );
  CLKBUFX3 U43842 ( .A(net218936), .Y(net218924) );
  CLKBUFX3 U43843 ( .A(net218936), .Y(net218922) );
  CLKBUFX3 U43844 ( .A(net218938), .Y(net218920) );
  CLKBUFX3 U43845 ( .A(net218952), .Y(net218878) );
  CLKBUFX3 U43846 ( .A(net218950), .Y(net218882) );
  CLKBUFX3 U43847 ( .A(net218950), .Y(net218880) );
  CLKBUFX3 U43848 ( .A(net218954), .Y(net218870) );
  CLKBUFX3 U43849 ( .A(net218952), .Y(net218876) );
  CLKBUFX3 U43850 ( .A(net218952), .Y(net218874) );
  CLKBUFX3 U43851 ( .A(net218954), .Y(net218872) );
  CLKBUFX3 U43852 ( .A(net218946), .Y(net218894) );
  CLKBUFX3 U43853 ( .A(net218944), .Y(net218900) );
  CLKBUFX3 U43854 ( .A(net218944), .Y(net218898) );
  CLKBUFX3 U43855 ( .A(net218946), .Y(net218896) );
  CLKBUFX3 U43856 ( .A(net218950), .Y(net218884) );
  CLKBUFX3 U43857 ( .A(net218946), .Y(net218892) );
  CLKBUFX3 U43858 ( .A(net218954), .Y(net218868) );
  CLKBUFX3 U43859 ( .A(net217278), .Y(net217254) );
  CLKBUFX3 U43860 ( .A(net217280), .Y(net217264) );
  CLKBUFX3 U43861 ( .A(net217278), .Y(net217256) );
  CLKBUFX3 U43862 ( .A(net217278), .Y(net217258) );
  CLKBUFX3 U43863 ( .A(net217280), .Y(net217260) );
  CLKBUFX3 U43864 ( .A(net217280), .Y(net217262) );
  CLKBUFX3 U43865 ( .A(net217282), .Y(net217270) );
  CLKBUFX3 U43866 ( .A(net217282), .Y(net217268) );
  CLKBUFX3 U43867 ( .A(net217282), .Y(net217266) );
  CLKBUFX3 U43868 ( .A(net218292), .Y(net218282) );
  CLKBUFX3 U43869 ( .A(net218292), .Y(net218284) );
  CLKBUFX3 U43870 ( .A(n43036), .Y(n43025) );
  CLKBUFX3 U43871 ( .A(n43036), .Y(n43024) );
  CLKBUFX3 U43872 ( .A(n43035), .Y(n43026) );
  CLKBUFX3 U43873 ( .A(n43035), .Y(n43027) );
  CLKBUFX3 U43874 ( .A(n43035), .Y(n43028) );
  CLKBUFX3 U43875 ( .A(net218562), .Y(net218368) );
  CLKBUFX3 U43876 ( .A(net218562), .Y(net218370) );
  CLKBUFX3 U43877 ( .A(net218560), .Y(net218376) );
  CLKBUFX3 U43878 ( .A(net218560), .Y(net218378) );
  CLKBUFX3 U43879 ( .A(net218566), .Y(net218352) );
  CLKBUFX3 U43880 ( .A(net218566), .Y(net218354) );
  CLKBUFX3 U43881 ( .A(net218564), .Y(net218360) );
  CLKBUFX3 U43882 ( .A(net218556), .Y(net218394) );
  CLKBUFX3 U43883 ( .A(net218554), .Y(net218400) );
  CLKBUFX3 U43884 ( .A(net218554), .Y(net218402) );
  CLKBUFX3 U43885 ( .A(net218558), .Y(net218384) );
  CLKBUFX3 U43886 ( .A(net218558), .Y(net218386) );
  CLKBUFX3 U43887 ( .A(net218556), .Y(net218392) );
  CLKBUFX3 U43888 ( .A(net218576), .Y(net218312) );
  CLKBUFX3 U43889 ( .A(net218576), .Y(net218314) );
  CLKBUFX3 U43890 ( .A(net218574), .Y(net218320) );
  CLKBUFX3 U43891 ( .A(net218578), .Y(net218304) );
  CLKBUFX3 U43892 ( .A(net218570), .Y(net218338) );
  CLKBUFX3 U43893 ( .A(net218568), .Y(net218344) );
  CLKBUFX3 U43894 ( .A(net218568), .Y(net218346) );
  CLKBUFX3 U43895 ( .A(net218574), .Y(net218322) );
  CLKBUFX3 U43896 ( .A(net218572), .Y(net218328) );
  CLKBUFX3 U43897 ( .A(net218572), .Y(net218330) );
  CLKBUFX3 U43898 ( .A(net218570), .Y(net218336) );
  CLKBUFX3 U43899 ( .A(net218534), .Y(net218480) );
  CLKBUFX3 U43900 ( .A(net218534), .Y(net218482) );
  CLKBUFX3 U43901 ( .A(net218532), .Y(net218488) );
  CLKBUFX3 U43902 ( .A(net218532), .Y(net218490) );
  CLKBUFX3 U43903 ( .A(net218536), .Y(net218472) );
  CLKBUFX3 U43904 ( .A(net218536), .Y(net218474) );
  CLKBUFX3 U43905 ( .A(net218530), .Y(net218496) );
  CLKBUFX3 U43906 ( .A(net218528), .Y(net218504) );
  CLKBUFX3 U43907 ( .A(net218528), .Y(net218506) );
  CLKBUFX3 U43908 ( .A(net218548), .Y(net218424) );
  CLKBUFX3 U43909 ( .A(net218548), .Y(net218426) );
  CLKBUFX3 U43910 ( .A(net218546), .Y(net218432) );
  CLKBUFX3 U43911 ( .A(net218546), .Y(net218434) );
  CLKBUFX3 U43912 ( .A(net218552), .Y(net218408) );
  CLKBUFX3 U43913 ( .A(net218552), .Y(net218410) );
  CLKBUFX3 U43914 ( .A(net218550), .Y(net218416) );
  CLKBUFX3 U43915 ( .A(net218550), .Y(net218418) );
  CLKBUFX3 U43916 ( .A(net218540), .Y(net218456) );
  CLKBUFX3 U43917 ( .A(net218540), .Y(net218458) );
  CLKBUFX3 U43918 ( .A(net218538), .Y(net218464) );
  CLKBUFX3 U43919 ( .A(net218544), .Y(net218440) );
  CLKBUFX3 U43920 ( .A(net218544), .Y(net218442) );
  CLKBUFX3 U43921 ( .A(net218542), .Y(net218450) );
  CLKBUFX3 U43922 ( .A(net218294), .Y(net218296) );
  CLKBUFX3 U43923 ( .A(net218294), .Y(net218298) );
  CLKBUFX3 U43924 ( .A(net218562), .Y(net218366) );
  CLKBUFX3 U43925 ( .A(net218560), .Y(net218372) );
  CLKBUFX3 U43926 ( .A(net218560), .Y(net218374) );
  CLKBUFX3 U43927 ( .A(net218564), .Y(net218356) );
  CLKBUFX3 U43928 ( .A(net218564), .Y(net218358) );
  CLKBUFX3 U43929 ( .A(net218562), .Y(net218364) );
  CLKBUFX3 U43930 ( .A(net218554), .Y(net218396) );
  CLKBUFX3 U43931 ( .A(net218554), .Y(net218398) );
  CLKBUFX3 U43932 ( .A(net218552), .Y(net218404) );
  CLKBUFX3 U43933 ( .A(net218552), .Y(net218406) );
  CLKBUFX3 U43934 ( .A(net218558), .Y(net218380) );
  CLKBUFX3 U43935 ( .A(net218556), .Y(net218388) );
  CLKBUFX3 U43936 ( .A(net218576), .Y(net218310) );
  CLKBUFX3 U43937 ( .A(net218574), .Y(net218316) );
  CLKBUFX3 U43938 ( .A(net218578), .Y(net218300) );
  CLKBUFX3 U43939 ( .A(net218578), .Y(net218302) );
  CLKBUFX3 U43940 ( .A(net218576), .Y(net218308) );
  CLKBUFX3 U43941 ( .A(net218568), .Y(net218340) );
  CLKBUFX3 U43942 ( .A(net218568), .Y(net218342) );
  CLKBUFX3 U43943 ( .A(net218566), .Y(net218348) );
  CLKBUFX3 U43944 ( .A(net218566), .Y(net218350) );
  CLKBUFX3 U43945 ( .A(net218572), .Y(net218324) );
  CLKBUFX3 U43946 ( .A(net218572), .Y(net218326) );
  CLKBUFX3 U43947 ( .A(net218570), .Y(net218332) );
  CLKBUFX3 U43948 ( .A(net218570), .Y(net218334) );
  CLKBUFX3 U43949 ( .A(net218532), .Y(net218484) );
  CLKBUFX3 U43950 ( .A(net218532), .Y(net218486) );
  CLKBUFX3 U43951 ( .A(net218536), .Y(net218468) );
  CLKBUFX3 U43952 ( .A(net218534), .Y(net218476) );
  CLKBUFX3 U43953 ( .A(net218534), .Y(net218478) );
  CLKBUFX3 U43954 ( .A(net218530), .Y(net218494) );
  CLKBUFX3 U43955 ( .A(net218528), .Y(net218500) );
  CLKBUFX3 U43956 ( .A(net218528), .Y(net218502) );
  CLKBUFX3 U43957 ( .A(net218546), .Y(net218428) );
  CLKBUFX3 U43958 ( .A(net218546), .Y(net218430) );
  CLKBUFX3 U43959 ( .A(net218550), .Y(net218412) );
  CLKBUFX3 U43960 ( .A(net218550), .Y(net218414) );
  CLKBUFX3 U43961 ( .A(net218548), .Y(net218420) );
  CLKBUFX3 U43962 ( .A(net218548), .Y(net218422) );
  CLKBUFX3 U43963 ( .A(net218540), .Y(net218452) );
  CLKBUFX3 U43964 ( .A(net218540), .Y(net218454) );
  CLKBUFX3 U43965 ( .A(net218538), .Y(net218462) );
  CLKBUFX3 U43966 ( .A(net218544), .Y(net218438) );
  CLKBUFX3 U43967 ( .A(net218542), .Y(net218446) );
  CLKBUFX3 U43968 ( .A(net217284), .Y(net217272) );
  CLKBUFX3 U43969 ( .A(net217284), .Y(net217274) );
  CLKBUFX3 U43970 ( .A(net217284), .Y(net217276) );
  CLKBUFX3 U43971 ( .A(n43024), .Y(n43032) );
  CLKBUFX3 U43972 ( .A(net218582), .Y(net218580) );
  CLKBUFX3 U43973 ( .A(net218962), .Y(net218952) );
  CLKBUFX3 U43974 ( .A(net218962), .Y(net218954) );
  CLKBUFX3 U43975 ( .A(net218958), .Y(net218940) );
  CLKBUFX3 U43976 ( .A(net218958), .Y(net218942) );
  CLKBUFX3 U43977 ( .A(net218956), .Y(net218934) );
  CLKBUFX3 U43978 ( .A(net218956), .Y(net218936) );
  CLKBUFX3 U43979 ( .A(net218956), .Y(net218938) );
  CLKBUFX3 U43980 ( .A(net218958), .Y(net218944) );
  CLKBUFX3 U43981 ( .A(net218960), .Y(net218950) );
  CLKBUFX3 U43982 ( .A(net218960), .Y(net218946) );
  CLKBUFX3 U43983 ( .A(net218960), .Y(net218948) );
  CLKBUFX3 U43984 ( .A(net217288), .Y(net217280) );
  CLKBUFX3 U43985 ( .A(n43037), .Y(n43035) );
  CLKBUFX3 U43986 ( .A(n43037), .Y(n43034) );
  CLKBUFX3 U43987 ( .A(n43037), .Y(n43036) );
  CLKBUFX3 U43988 ( .A(net218526), .Y(net218512) );
  CLKBUFX3 U43989 ( .A(net218524), .Y(net218518) );
  CLKBUFX3 U43990 ( .A(net218524), .Y(net218520) );
  CLKBUFX3 U43991 ( .A(net218588), .Y(net218560) );
  CLKBUFX3 U43992 ( .A(net218586), .Y(net218564) );
  CLKBUFX3 U43993 ( .A(net218588), .Y(net218562) );
  CLKBUFX3 U43994 ( .A(net218590), .Y(net218554) );
  CLKBUFX3 U43995 ( .A(net218588), .Y(net218558) );
  CLKBUFX3 U43996 ( .A(net218590), .Y(net218556) );
  CLKBUFX3 U43997 ( .A(net218582), .Y(net218578) );
  CLKBUFX3 U43998 ( .A(net218582), .Y(net218576) );
  CLKBUFX3 U43999 ( .A(net218586), .Y(net218568) );
  CLKBUFX3 U44000 ( .A(net218586), .Y(net218566) );
  CLKBUFX3 U44001 ( .A(net218584), .Y(net218574) );
  CLKBUFX3 U44002 ( .A(net218584), .Y(net218572) );
  CLKBUFX3 U44003 ( .A(net218584), .Y(net218570) );
  CLKBUFX3 U44004 ( .A(net218598), .Y(net218532) );
  CLKBUFX3 U44005 ( .A(net218596), .Y(net218536) );
  CLKBUFX3 U44006 ( .A(net218596), .Y(net218534) );
  CLKBUFX3 U44007 ( .A(net218598), .Y(net218530) );
  CLKBUFX3 U44008 ( .A(net218598), .Y(net218528) );
  CLKBUFX3 U44009 ( .A(net218592), .Y(net218546) );
  CLKBUFX3 U44010 ( .A(net218590), .Y(net218552) );
  CLKBUFX3 U44011 ( .A(net218592), .Y(net218550) );
  CLKBUFX3 U44012 ( .A(net218592), .Y(net218548) );
  CLKBUFX3 U44013 ( .A(net218594), .Y(net218540) );
  CLKBUFX3 U44014 ( .A(net218596), .Y(net218538) );
  CLKBUFX3 U44015 ( .A(net218594), .Y(net218544) );
  CLKBUFX3 U44016 ( .A(net218594), .Y(net218542) );
  CLKBUFX3 U44017 ( .A(net218526), .Y(net218508) );
  CLKBUFX3 U44018 ( .A(net218526), .Y(net218510) );
  CLKBUFX3 U44019 ( .A(net218524), .Y(net218516) );
  CLKBUFX3 U44020 ( .A(n43037), .Y(n43033) );
  INVX3 U44021 ( .A(net221974), .Y(net221788) );
  CLKINVX1 U44022 ( .A(n9790), .Y(n49493) );
  NAND2BX1 U44023 ( .AN(net210705), .B(net171380), .Y(n9874) );
  CLKBUFX3 U44024 ( .A(n9782), .Y(net217288) );
  CLKBUFX3 U44025 ( .A(n9782), .Y(net217286) );
  NAND4X1 U44026 ( .A(n9931), .B(n24671), .C(n9825), .D(n49494), .Y(n9790) );
  NOR2X1 U44027 ( .A(n9829), .B(n9820), .Y(n24671) );
  NOR2X1 U44028 ( .A(net264532), .B(net171380), .Y(n9754) );
  CLKINVX1 U44029 ( .A(n9935), .Y(n49519) );
  CLKINVX1 U44030 ( .A(n47842), .Y(n47845) );
  CLKBUFX3 U44031 ( .A(net218588), .Y(net218526) );
  CLKBUFX3 U44032 ( .A(net221976), .Y(net221906) );
  CLKINVX1 U44033 ( .A(n9791), .Y(n50118) );
  CLKBUFX3 U44034 ( .A(net218590), .Y(net218524) );
  CLKBUFX3 U44035 ( .A(net218604), .Y(net218588) );
  CLKBUFX3 U44036 ( .A(net218606), .Y(net218598) );
  CLKBUFX3 U44037 ( .A(net218604), .Y(net218590) );
  CLKBUFX3 U44038 ( .A(net218604), .Y(net218592) );
  CLKBUFX3 U44039 ( .A(net218606), .Y(net218596) );
  CLKBUFX3 U44040 ( .A(net218606), .Y(net218594) );
  CLKINVX1 U44041 ( .A(n9852), .Y(n43037) );
  CLKINVX1 U44042 ( .A(n9943), .Y(n50120) );
  CLKINVX1 U44043 ( .A(n9931), .Y(n50126) );
  CLKINVX1 U44044 ( .A(n9825), .Y(n50125) );
  CLKBUFX3 U44045 ( .A(net221972), .Y(net221920) );
  CLKBUFX3 U44046 ( .A(net221972), .Y(net221922) );
  CLKBUFX3 U44047 ( .A(net221970), .Y(net221924) );
  CLKBUFX3 U44048 ( .A(net221970), .Y(net221926) );
  CLKBUFX3 U44049 ( .A(net221970), .Y(net221928) );
  CLKBUFX3 U44050 ( .A(net221968), .Y(net221930) );
  CLKBUFX3 U44051 ( .A(net221976), .Y(net221910) );
  CLKBUFX3 U44052 ( .A(net221976), .Y(net221908) );
  CLKBUFX3 U44053 ( .A(net221974), .Y(net221912) );
  CLKBUFX3 U44054 ( .A(net221974), .Y(net221914) );
  CLKBUFX3 U44055 ( .A(net221974), .Y(net221916) );
  CLKBUFX3 U44056 ( .A(net221972), .Y(net221918) );
  CLKBUFX3 U44057 ( .A(net221964), .Y(net221946) );
  CLKBUFX3 U44058 ( .A(net221962), .Y(net221948) );
  CLKBUFX3 U44059 ( .A(net221962), .Y(net221950) );
  CLKBUFX3 U44060 ( .A(net221962), .Y(net221952) );
  CLKBUFX3 U44061 ( .A(net221960), .Y(net221954) );
  CLKBUFX3 U44062 ( .A(net221960), .Y(net221956) );
  CLKBUFX3 U44063 ( .A(net221968), .Y(net221932) );
  CLKBUFX3 U44064 ( .A(net221968), .Y(net221934) );
  CLKBUFX3 U44065 ( .A(net221966), .Y(net221936) );
  CLKBUFX3 U44066 ( .A(net221966), .Y(net221938) );
  CLKBUFX3 U44067 ( .A(net221966), .Y(net221940) );
  CLKBUFX3 U44068 ( .A(net221964), .Y(net221942) );
  CLKBUFX3 U44069 ( .A(net221964), .Y(net221944) );
  CLKBUFX3 U44070 ( .A(n42647), .Y(n42651) );
  CLKBUFX3 U44071 ( .A(n42498), .Y(n42493) );
  OAI21XL U44072 ( .A0(n48382), .A1(n48381), .B0(n48380), .Y(n48385) );
  NOR4X1 U44073 ( .A(n48379), .B(n48378), .C(n48377), .D(n48376), .Y(n48380)
         );
  OAI21XL U44074 ( .A0(net209504), .A1(n48375), .B0(n48374), .Y(n48381) );
  AOI21X1 U44075 ( .A0(n48366), .A1(n48365), .B0(n48364), .Y(n48382) );
  CLKBUFX3 U44076 ( .A(n42480), .Y(n42492) );
  CLKINVX1 U44077 ( .A(net207642), .Y(net171301) );
  CLKBUFX3 U44078 ( .A(n42490), .Y(n42486) );
  CLKINVX1 U44079 ( .A(n10094), .Y(net151263) );
  CLKBUFX3 U44080 ( .A(n42667), .Y(n42657) );
  CLKINVX1 U44081 ( .A(net209402), .Y(net172112) );
  AOI211X1 U44082 ( .A0(n9942), .A1(n10071), .B0(n10072), .C0(n10073), .Y(
        n10069) );
  OAI21XL U44083 ( .A0(n10074), .A1(n10075), .B0(n10076), .Y(n10071) );
  NOR4BX1 U44084 ( .AN(n10077), .B(n10078), .C(n40404), .D(n10080), .Y(n10074)
         );
  AOI211X1 U44085 ( .A0(n9931), .A1(n10081), .B0(n10082), .C0(n10083), .Y(
        n10078) );
  NOR4X1 U44086 ( .A(n10099), .B(net171198), .C(n10101), .D(n10102), .Y(n10095) );
  AOI211X1 U44087 ( .A0(n10103), .A1(n10104), .B0(n10105), .C0(n40403), .Y(
        n10099) );
  OAI21XL U44088 ( .A0(n10107), .A1(n10108), .B0(n10109), .Y(n10104) );
  AOI211X1 U44089 ( .A0(n10110), .A1(n10111), .B0(n10112), .C0(n10113), .Y(
        n10107) );
  OAI31XL U44090 ( .A0(n9815), .A1(n9816), .A2(n9817), .B0(n50119), .Y(n9813)
         );
  CLKINVX1 U44091 ( .A(n9819), .Y(n50119) );
  OAI31XL U44092 ( .A0(n9820), .A1(n9821), .A2(n50125), .B0(n50123), .Y(n9815)
         );
  NAND2X1 U44093 ( .A(net266235), .B(n43043), .Y(n9744) );
  OAI21XL U44094 ( .A0(n42697), .A1(n40176), .B0(n13063), .Y(n48715) );
  CLKBUFX3 U44095 ( .A(n42696), .Y(n42694) );
  CLKBUFX3 U44096 ( .A(n42661), .Y(n42654) );
  CLKBUFX3 U44097 ( .A(n36711), .Y(n42606) );
  CLKINVX1 U44098 ( .A(n48873), .Y(n48553) );
  CLKBUFX3 U44099 ( .A(n10058), .Y(net218602) );
  CLKBUFX3 U44100 ( .A(n10197), .Y(net218966) );
  CLKBUFX3 U44101 ( .A(n10197), .Y(net218964) );
  NAND3BX1 U44102 ( .AN(n10112), .B(net168850), .C(n10110), .Y(n9794) );
  NOR3BX1 U44103 ( .AN(n10293), .B(n10295), .C(net171280), .Y(n9943) );
  NOR2BX1 U44104 ( .AN(n10076), .B(n10075), .Y(n9825) );
  NAND4X1 U44105 ( .A(net151263), .B(net151265), .C(n10091), .D(n24675), .Y(
        n9829) );
  NOR4X1 U44106 ( .A(net151264), .B(net151266), .C(n10093), .D(n10085), .Y(
        n24675) );
  NAND3BX1 U44107 ( .AN(n10105), .B(n10103), .C(net151404), .Y(n9791) );
  NAND3BX1 U44108 ( .AN(n10082), .B(n10077), .C(n24672), .Y(n9820) );
  NOR3X1 U44109 ( .A(n10080), .B(n10083), .C(n40404), .Y(n24672) );
  OAI31XL U44110 ( .A0(n50120), .A1(n9924), .A2(n9819), .B0(n50117), .Y(n9923)
         );
  CLKINVX1 U44111 ( .A(n9812), .Y(n50117) );
  AOI211X1 U44112 ( .A0(n50124), .A1(n9927), .B0(n9816), .C0(n9824), .Y(n9924)
         );
  CLKINVX1 U44113 ( .A(n9817), .Y(n50124) );
  NOR4X1 U44114 ( .A(n10311), .B(net171169), .C(n_cell_301249_net269488), .D(
        net171168), .Y(n10129) );
  CLKINVX1 U44115 ( .A(net260384), .Y(net171349) );
  NOR2X1 U44116 ( .A(n10334), .B(n10338), .Y(n9931) );
  NOR2BX1 U44117 ( .AN(n10109), .B(n10108), .Y(n9935) );
  NAND2X1 U44118 ( .A(n24683), .B(n24684), .Y(n9781) );
  NOR4X1 U44119 ( .A(n9824), .B(n9816), .C(n9819), .D(n9812), .Y(n24684) );
  AND4X1 U44120 ( .A(net168846), .B(net168848), .C(n10129), .D(n9943), .Y(
        n24683) );
  NOR4X1 U44121 ( .A(n9826), .B(n50126), .C(n9828), .D(n9829), .Y(n9821) );
  NOR3X1 U44122 ( .A(n9792), .B(n9830), .C(n9791), .Y(n9826) );
  AOI211X1 U44123 ( .A0(n49495), .A1(n9832), .B0(n9794), .C0(n49519), .Y(n9830) );
  CLKINVX1 U44124 ( .A(n47847), .Y(n49495) );
  CLKINVX1 U44125 ( .A(n9828), .Y(n49494) );
  OR2X1 U44126 ( .A(n41737), .B(n9938), .Y(n47847) );
  OR2X1 U44127 ( .A(n9939), .B(n47839), .Y(n41737) );
  OAI21XL U44128 ( .A0(n9928), .A1(n9820), .B0(n9825), .Y(n9927) );
  AOI211X1 U44129 ( .A0(n50127), .A1(n9930), .B0(n9828), .C0(n50126), .Y(n9928) );
  CLKINVX1 U44130 ( .A(n9829), .Y(n50127) );
  AO21X1 U44131 ( .A0(n50118), .A1(n9933), .B0(n9792), .Y(n9930) );
  CLKBUFX3 U44132 ( .A(n50114), .Y(n42454) );
  CLKBUFX3 U44133 ( .A(n50082), .Y(n42450) );
  CLKBUFX3 U44134 ( .A(n50082), .Y(n42451) );
  CLKBUFX3 U44135 ( .A(n42483), .Y(n42488) );
  CLKBUFX3 U44136 ( .A(n50114), .Y(n42453) );
  CLKBUFX3 U44137 ( .A(n50114), .Y(n42452) );
  CLKBUFX3 U44138 ( .A(n42465), .Y(n42464) );
  CLKBUFX3 U44139 ( .A(n42465), .Y(n42463) );
  NAND2BX1 U44140 ( .AN(n47824), .B(n41744), .Y(n47842) );
  CLKBUFX3 U44141 ( .A(n10058), .Y(net218604) );
  CLKBUFX3 U44142 ( .A(n10058), .Y(net218606) );
  CLKBUFX3 U44143 ( .A(net221982), .Y(net221980) );
  CLKBUFX3 U44144 ( .A(net221982), .Y(net221976) );
  NAND3X1 U44145 ( .A(net168848), .B(net168846), .C(n9942), .Y(n9817) );
  CLKINVX1 U44146 ( .A(n9816), .Y(n50121) );
  CLKINVX1 U44147 ( .A(n9824), .Y(n50123) );
  CLKBUFX3 U44148 ( .A(net221982), .Y(net221978) );
  CLKBUFX3 U44149 ( .A(net221984), .Y(net221970) );
  CLKBUFX3 U44150 ( .A(net221984), .Y(net221974) );
  CLKBUFX3 U44151 ( .A(net221984), .Y(net221972) );
  CLKBUFX3 U44152 ( .A(net221986), .Y(net221968) );
  CLKBUFX3 U44153 ( .A(net221986), .Y(net221966) );
  CLKBUFX3 U44154 ( .A(net221986), .Y(net221964) );
  CLKBUFX3 U44155 ( .A(net221988), .Y(net221962) );
  CLKBUFX3 U44156 ( .A(net221988), .Y(net221960) );
  CLKBUFX3 U44157 ( .A(n42413), .Y(n42412) );
  CLKBUFX3 U44158 ( .A(n42414), .Y(n42411) );
  CLKBUFX3 U44159 ( .A(n42414), .Y(n42410) );
  CLKBUFX3 U44160 ( .A(n42414), .Y(n42409) );
  CLKBUFX3 U44161 ( .A(n42415), .Y(n42408) );
  CLKBUFX3 U44162 ( .A(n42415), .Y(n42407) );
  CLKBUFX3 U44163 ( .A(n42415), .Y(n42406) );
  CLKBUFX3 U44164 ( .A(n42415), .Y(n42405) );
  CLKBUFX3 U44165 ( .A(n42416), .Y(n42404) );
  CLKBUFX3 U44166 ( .A(n42416), .Y(n42403) );
  CLKBUFX3 U44167 ( .A(n42416), .Y(n42402) );
  CLKBUFX3 U44168 ( .A(n42417), .Y(n42401) );
  CLKBUFX3 U44169 ( .A(n42418), .Y(n42400) );
  CLKBUFX3 U44170 ( .A(n42419), .Y(n42399) );
  CLKBUFX3 U44171 ( .A(n42419), .Y(n42398) );
  CLKBUFX3 U44172 ( .A(n42420), .Y(n42397) );
  CLKBUFX3 U44173 ( .A(n42420), .Y(n42396) );
  CLKBUFX3 U44174 ( .A(n42420), .Y(n42395) );
  CLKBUFX3 U44175 ( .A(n42420), .Y(n42394) );
  CLKBUFX3 U44176 ( .A(n42421), .Y(n42393) );
  CLKBUFX3 U44177 ( .A(n42421), .Y(n42392) );
  CLKBUFX3 U44178 ( .A(n42421), .Y(n42391) );
  CLKBUFX3 U44179 ( .A(n42446), .Y(n42390) );
  CLKBUFX3 U44180 ( .A(n49523), .Y(n42389) );
  CLKBUFX3 U44181 ( .A(n42446), .Y(n42388) );
  CLKBUFX3 U44182 ( .A(n42417), .Y(n42387) );
  CLKBUFX3 U44183 ( .A(n42422), .Y(n42386) );
  CLKBUFX3 U44184 ( .A(n42422), .Y(n42385) );
  CLKBUFX3 U44185 ( .A(n42422), .Y(n42384) );
  CLKBUFX3 U44186 ( .A(n42422), .Y(n42383) );
  CLKBUFX3 U44187 ( .A(n42423), .Y(n42382) );
  CLKBUFX3 U44188 ( .A(n42423), .Y(n42381) );
  CLKBUFX3 U44189 ( .A(n42423), .Y(n42380) );
  CLKBUFX3 U44190 ( .A(n42423), .Y(n42379) );
  CLKBUFX3 U44191 ( .A(n42424), .Y(n42378) );
  CLKBUFX3 U44192 ( .A(n42424), .Y(n42377) );
  CLKBUFX3 U44193 ( .A(n42424), .Y(n42376) );
  CLKBUFX3 U44194 ( .A(n42424), .Y(n42375) );
  CLKBUFX3 U44195 ( .A(n42444), .Y(n42374) );
  CLKBUFX3 U44196 ( .A(n42418), .Y(n42373) );
  CLKBUFX3 U44197 ( .A(n42425), .Y(n42372) );
  CLKBUFX3 U44198 ( .A(n42425), .Y(n42371) );
  CLKBUFX3 U44199 ( .A(n42425), .Y(n42370) );
  CLKBUFX3 U44200 ( .A(n42425), .Y(n42369) );
  CLKBUFX3 U44201 ( .A(n42426), .Y(n42368) );
  CLKBUFX3 U44202 ( .A(n42426), .Y(n42367) );
  CLKBUFX3 U44203 ( .A(n42426), .Y(n42366) );
  CLKBUFX3 U44204 ( .A(n42426), .Y(n42365) );
  CLKBUFX3 U44205 ( .A(n42436), .Y(n42364) );
  CLKBUFX3 U44206 ( .A(n42443), .Y(n42363) );
  CLKBUFX3 U44207 ( .A(n42442), .Y(n42362) );
  CLKBUFX3 U44208 ( .A(n42438), .Y(n42361) );
  CLKBUFX3 U44209 ( .A(n42427), .Y(n42360) );
  CLKBUFX3 U44210 ( .A(n42427), .Y(n42359) );
  CLKBUFX3 U44211 ( .A(n42427), .Y(n42358) );
  CLKBUFX3 U44212 ( .A(n42427), .Y(n42357) );
  CLKBUFX3 U44213 ( .A(n42428), .Y(n42356) );
  CLKBUFX3 U44214 ( .A(n42428), .Y(n42355) );
  CLKBUFX3 U44215 ( .A(n42428), .Y(n42354) );
  CLKBUFX3 U44216 ( .A(n42428), .Y(n42353) );
  CLKBUFX3 U44217 ( .A(n42429), .Y(n42352) );
  CLKBUFX3 U44218 ( .A(n42429), .Y(n42351) );
  CLKBUFX3 U44219 ( .A(n42429), .Y(n42350) );
  CLKBUFX3 U44220 ( .A(n42413), .Y(n42349) );
  CLKBUFX3 U44221 ( .A(n42430), .Y(n42348) );
  CLKBUFX3 U44222 ( .A(n42430), .Y(n42347) );
  CLKBUFX3 U44223 ( .A(n42430), .Y(n42346) );
  CLKBUFX3 U44224 ( .A(n42431), .Y(n42345) );
  CLKBUFX3 U44225 ( .A(n42431), .Y(n42344) );
  CLKBUFX3 U44226 ( .A(n42431), .Y(n42343) );
  CLKBUFX3 U44227 ( .A(n42431), .Y(n42342) );
  CLKBUFX3 U44228 ( .A(n42432), .Y(n42341) );
  CLKBUFX3 U44229 ( .A(n42432), .Y(n42340) );
  CLKBUFX3 U44230 ( .A(n42432), .Y(n42339) );
  CLKBUFX3 U44231 ( .A(n42439), .Y(n42338) );
  CLKBUFX3 U44232 ( .A(n42438), .Y(n42337) );
  CLKBUFX3 U44233 ( .A(n42433), .Y(n42336) );
  CLKBUFX3 U44234 ( .A(n42433), .Y(n42335) );
  CLKBUFX3 U44235 ( .A(n42433), .Y(n42334) );
  CLKBUFX3 U44236 ( .A(n42433), .Y(n42333) );
  CLKBUFX3 U44237 ( .A(n42434), .Y(n42332) );
  CLKBUFX3 U44238 ( .A(n42434), .Y(n42331) );
  CLKBUFX3 U44239 ( .A(n42434), .Y(n42330) );
  CLKBUFX3 U44240 ( .A(n42434), .Y(n42329) );
  CLKBUFX3 U44241 ( .A(n42435), .Y(n42328) );
  CLKBUFX3 U44242 ( .A(n42435), .Y(n42327) );
  CLKBUFX3 U44243 ( .A(n42435), .Y(n42326) );
  CLKBUFX3 U44244 ( .A(n42435), .Y(n42325) );
  CLKBUFX3 U44245 ( .A(n42436), .Y(n42324) );
  CLKBUFX3 U44246 ( .A(n42439), .Y(n42323) );
  CLKBUFX3 U44247 ( .A(n42436), .Y(n42322) );
  NAND2X1 U44248 ( .A(n11723), .B(net207642), .Y(n11720) );
  NAND2X1 U44249 ( .A(n11699), .B(n11700), .Y(n11696) );
  CLKINVX1 U44250 ( .A(n11705), .Y(net151330) );
  NAND2X1 U44251 ( .A(n11661), .B(n11662), .Y(n11660) );
  NAND2X1 U44252 ( .A(n11651), .B(n11652), .Y(n11648) );
  CLKINVX1 U44253 ( .A(n11658), .Y(net151271) );
  AND2X2 U44254 ( .A(n11849), .B(n11850), .Y(n11745) );
  CLKINVX1 U44255 ( .A(n11646), .Y(net151249) );
  NAND2X1 U44256 ( .A(n11687), .B(n11688), .Y(n11684) );
  CLKINVX1 U44257 ( .A(n12582), .Y(net171231) );
  CLKINVX1 U44258 ( .A(n48337), .Y(n48295) );
  CLKBUFX3 U44259 ( .A(n41629), .Y(n42572) );
  CLKINVX1 U44260 ( .A(n10394), .Y(net151340) );
  CLKBUFX3 U44261 ( .A(n42528), .Y(n42525) );
  INVX3 U44262 ( .A(n42509), .Y(n42507) );
  INVX3 U44263 ( .A(n42585), .Y(n42582) );
  INVX3 U44264 ( .A(n42621), .Y(n42619) );
  INVX3 U44265 ( .A(n42545), .Y(n42543) );
  INVX3 U44266 ( .A(n42555), .Y(n42553) );
  INVX3 U44267 ( .A(n42685), .Y(n42683) );
  INVX3 U44268 ( .A(n42677), .Y(n42674) );
  INVX3 U44269 ( .A(n42713), .Y(n42710) );
  INVX3 U44270 ( .A(n36920), .Y(n42504) );
  INVX3 U44271 ( .A(n42555), .Y(n42554) );
  INVX3 U44272 ( .A(n42585), .Y(n42584) );
  INVX3 U44273 ( .A(n42556), .Y(n42547) );
  INVX3 U44274 ( .A(n42726), .Y(n42725) );
  INVX3 U44275 ( .A(n42621), .Y(n42620) );
  INVX3 U44276 ( .A(n42509), .Y(n42508) );
  CLKBUFX3 U44277 ( .A(n42512), .Y(n42531) );
  CLKBUFX3 U44278 ( .A(n42477), .Y(n42497) );
  CLKBUFX3 U44279 ( .A(n42455), .Y(n42474) );
  CLKINVX1 U44280 ( .A(n10384), .Y(net171237) );
  CLKINVX1 U44281 ( .A(n12583), .Y(net171189) );
  CLKINVX1 U44282 ( .A(n12530), .Y(n49507) );
  CLKINVX1 U44283 ( .A(n12479), .Y(n48394) );
  CLKINVX1 U44284 ( .A(n12476), .Y(n48397) );
  CLKINVX1 U44285 ( .A(n11651), .Y(net209469) );
  CLKINVX1 U44286 ( .A(n11669), .Y(net209482) );
  NAND2X1 U44287 ( .A(n11685), .B(n48383), .Y(n48384) );
  CLKINVX1 U44288 ( .A(n12486), .Y(net209486) );
  NOR4X1 U44289 ( .A(n48358), .B(n48357), .C(n48356), .D(n48355), .Y(n48359)
         );
  NAND2X1 U44290 ( .A(n12539), .B(n12542), .Y(n11761) );
  CLKINVX1 U44291 ( .A(n10385), .Y(net171238) );
  CLKBUFX3 U44292 ( .A(n42573), .Y(n42571) );
  INVX3 U44293 ( .A(n42509), .Y(n42506) );
  INVX3 U44294 ( .A(n42545), .Y(n42541) );
  INVX3 U44295 ( .A(n42585), .Y(n42581) );
  INVX3 U44296 ( .A(n42545), .Y(n42540) );
  INVX3 U44297 ( .A(n42545), .Y(n42535) );
  INVX3 U44298 ( .A(n42687), .Y(n42682) );
  CLKBUFX3 U44299 ( .A(n42456), .Y(n42476) );
  CLKINVX1 U44300 ( .A(n12585), .Y(net171309) );
  CLKINVX1 U44301 ( .A(n10422), .Y(net209517) );
  CLKINVX1 U44302 ( .A(n11722), .Y(net209504) );
  CLKINVX1 U44303 ( .A(n48383), .Y(n49506) );
  CLKINVX1 U44304 ( .A(n48370), .Y(n49504) );
  CLKINVX1 U44305 ( .A(n12587), .Y(net171211) );
  CLKINVX1 U44306 ( .A(n12586), .Y(n49505) );
  CLKINVX1 U44307 ( .A(n44598), .Y(n49502) );
  CLKINVX1 U44308 ( .A(n12542), .Y(n48354) );
  CLKINVX1 U44309 ( .A(n11687), .Y(net209663) );
  CLKINVX1 U44310 ( .A(n11693), .Y(net209664) );
  CLKINVX1 U44311 ( .A(n10382), .Y(net209543) );
  OAI21XL U44312 ( .A0(net171237), .A1(n48350), .B0(n10385), .Y(n48351) );
  CLKINVX1 U44313 ( .A(n11700), .Y(net209669) );
  CLKINVX1 U44314 ( .A(n10424), .Y(net209516) );
  NAND2X1 U44315 ( .A(n11744), .B(n11741), .Y(n48286) );
  CLKINVX1 U44316 ( .A(n10393), .Y(net209549) );
  CLKINVX1 U44317 ( .A(n12535), .Y(net209661) );
  CLKINVX1 U44318 ( .A(n11712), .Y(net209676) );
  CLKINVX1 U44319 ( .A(n11717), .Y(net209675) );
  CLKINVX1 U44320 ( .A(n10369), .Y(net209520) );
  CLKINVX1 U44321 ( .A(n10387), .Y(net209557) );
  NAND4X1 U44322 ( .A(n48344), .B(n48343), .C(n48342), .D(n12549), .Y(n48345)
         );
  NOR2X1 U44323 ( .A(net151348), .B(n48354), .Y(n48344) );
  NOR2X1 U44324 ( .A(net171237), .B(net209557), .Y(n48343) );
  NOR2X1 U44325 ( .A(net209547), .B(net151340), .Y(n48342) );
  NOR2X1 U44326 ( .A(net171309), .B(net209507), .Y(n48374) );
  CLKINVX1 U44327 ( .A(n11721), .Y(net209507) );
  NAND4X1 U44328 ( .A(n48363), .B(n48362), .C(n48361), .D(n48360), .Y(n48364)
         );
  NOR3X1 U44329 ( .A(net209509), .B(net209504), .C(net171301), .Y(n48363) );
  NOR2X1 U44330 ( .A(n49504), .B(net209513), .Y(n48362) );
  AOI21X1 U44331 ( .A0(n11741), .A1(net209528), .B0(net209529), .Y(n48360) );
  NAND3X1 U44332 ( .A(n11699), .B(n11697), .C(n11706), .Y(n48377) );
  CLKINVX1 U44333 ( .A(n10383), .Y(net209546) );
  CLKINVX1 U44334 ( .A(n10423), .Y(net151356) );
  CLKINVX1 U44335 ( .A(n11742), .Y(net209528) );
  CLKINVX1 U44336 ( .A(n11849), .Y(n48283) );
  NOR2BX1 U44337 ( .AN(n12539), .B(net209537), .Y(n48352) );
  CLKINVX1 U44338 ( .A(n12506), .Y(n49500) );
  INVX3 U44339 ( .A(n42555), .Y(n42551) );
  INVX3 U44340 ( .A(n42545), .Y(n42539) );
  INVX3 U44341 ( .A(n42622), .Y(n42617) );
  INVX3 U44342 ( .A(n36920), .Y(n42503) );
  INVX3 U44343 ( .A(n42715), .Y(n42708) );
  CLKINVX1 U44344 ( .A(n11718), .Y(net151401) );
  CLKINVX1 U44345 ( .A(net214730), .Y(net171129) );
  CLKINVX1 U44346 ( .A(net214729), .Y(net171119) );
  CLKINVX1 U44347 ( .A(n11661), .Y(net171114) );
  CLKINVX1 U44348 ( .A(n11662), .Y(net171319) );
  CLKINVX1 U44349 ( .A(n10340), .Y(net171328) );
  CLKINVX1 U44350 ( .A(n12490), .Y(net151258) );
  CLKINVX1 U44351 ( .A(n12493), .Y(net151261) );
  CLKINVX1 U44352 ( .A(n12501), .Y(net171196) );
  INVX3 U44353 ( .A(n42727), .Y(n42720) );
  CLKINVX1 U44354 ( .A(n11706), .Y(net151333) );
  INVX3 U44355 ( .A(n42585), .Y(n42578) );
  INVX3 U44356 ( .A(n42593), .Y(n42588) );
  INVX3 U44357 ( .A(n42593), .Y(n42589) );
  CLKINVX1 U44358 ( .A(n11694), .Y(net151327) );
  CLKINVX1 U44359 ( .A(n12589), .Y(net171099) );
  CLKINVX1 U44360 ( .A(n12588), .Y(net171101) );
  CLKINVX1 U44361 ( .A(net209476), .Y(net171113) );
  CLKINVX1 U44362 ( .A(n12461), .Y(net171104) );
  CLKINVX1 U44363 ( .A(n12466), .Y(net171143) );
  NAND2X1 U44364 ( .A(n12476), .B(n12479), .Y(n10086) );
  CLKINVX1 U44365 ( .A(n12474), .Y(net151253) );
  NAND2X1 U44366 ( .A(n11668), .B(n11669), .Y(n11667) );
  CLKINVX1 U44367 ( .A(n11657), .Y(net151270) );
  OAI31XL U44368 ( .A0(n9780), .A1(n9781), .A2(n40313), .B0(n9783), .Y(n9779)
         );
  OAI21XL U44369 ( .A0(n9789), .A1(n9790), .B0(net260527), .Y(n9780) );
  NOR4X1 U44370 ( .A(n9791), .B(n9792), .C(n49519), .D(n9794), .Y(n9789) );
  AOI211X1 U44371 ( .A0(n9757), .A1(n9795), .B0(n50086), .C0(n9797), .Y(n9778)
         );
  NAND4X1 U44372 ( .A(n9798), .B(n9799), .C(n41758), .D(n50084), .Y(n9795) );
  NOR3BXL U44373 ( .AN(n50118), .B(n9781), .C(n49519), .Y(net213661) );
  NOR2X1 U44374 ( .A(n9790), .B(n47847), .Y(net213659) );
  NOR4BX1 U44375 ( .AN(net260527), .B(n9792), .C(n9794), .D(n9832), .Y(
        net213660) );
  OAI31XL U44376 ( .A0(n50083), .A1(n50104), .A2(n9763), .B0(n9764), .Y(n9760)
         );
  NAND4X1 U44377 ( .A(net216970), .B(n49497), .C(n49493), .D(net260527), .Y(
        n9764) );
  CLKINVX1 U44378 ( .A(n9770), .Y(n50083) );
  CLKINVX1 U44379 ( .A(n9781), .Y(n49497) );
  AOI21X1 U44380 ( .A0(n41742), .A1(n47840), .B0(n47815), .Y(n47817) );
  OAI21XL U44381 ( .A0(n50133), .A1(n43041), .B0(n43043), .Y(n9721) );
  NOR4BX1 U44382 ( .AN(n10064), .B(n10065), .C(n10066), .D(n10067), .Y(n10061)
         );
  AOI21X1 U44383 ( .A0(n9943), .A1(n10068), .B0(n9819), .Y(n10065) );
  OAI21XL U44384 ( .A0(n10069), .A1(n9824), .B0(n50121), .Y(n10068) );
  OAI31XL U44385 ( .A0(n10084), .A1(n10085), .A2(n10086), .B0(n49494), .Y(
        n10081) );
  NOR4BX1 U44386 ( .AN(n10091), .B(n10092), .C(n10093), .D(n10094), .Y(n10088)
         );
  NOR4X1 U44387 ( .A(n10095), .B(net171207), .C(n10097), .D(n10098), .Y(n10092) );
  NAND2X1 U44388 ( .A(net217930), .B(n42726), .Y(n49335) );
  NAND2X1 U44389 ( .A(n40192), .B(n42713), .Y(n49490) );
  NOR2X1 U44390 ( .A(net210516), .B(net210520), .Y(n41744) );
  NAND2X1 U44391 ( .A(n40272), .B(n41280), .Y(n48873) );
  NAND3X1 U44392 ( .A(n11685), .B(n11686), .C(n11679), .Y(n10097) );
  CLKINVX1 U44393 ( .A(net210481), .Y(net210435) );
  OAI21XL U44394 ( .A0(n10114), .A1(n9939), .B0(n50122), .Y(n10111) );
  CLKINVX1 U44395 ( .A(n9938), .Y(n50122) );
  NOR2X1 U44396 ( .A(n47821), .B(n47820), .Y(n10114) );
  NAND2X1 U44397 ( .A(n41743), .B(n10128), .Y(n47820) );
  NAND3X1 U44398 ( .A(n41750), .B(n45529), .C(n41742), .Y(n9832) );
  INVXL U44399 ( .A(n47840), .Y(n45529) );
  CLKINVX1 U44400 ( .A(net210494), .Y(net210443) );
  CLKINVX1 U44401 ( .A(n47843), .Y(n47846) );
  NAND3BX1 U44402 ( .AN(n9804), .B(n47844), .C(n47846), .Y(n47709) );
  CLKINVX1 U44403 ( .A(n12457), .Y(net151243) );
  CLKINVX1 U44404 ( .A(n12459), .Y(net151246) );
  NOR2X1 U44405 ( .A(n47819), .B(n47818), .Y(n47821) );
  NAND2X1 U44406 ( .A(net210424), .B(n37125), .Y(n47818) );
  NOR2X1 U44407 ( .A(n47817), .B(n47816), .Y(n47819) );
  NAND2X1 U44408 ( .A(n40276), .B(net219472), .Y(n49180) );
  NOR2X1 U44409 ( .A(net210416), .B(net210417), .Y(n47828) );
  CLKBUFX3 U44410 ( .A(n9719), .Y(n43043) );
  INVX3 U44411 ( .A(n41789), .Y(n43038) );
  INVX3 U44412 ( .A(n41790), .Y(n43041) );
  INVX3 U44413 ( .A(n41251), .Y(n42639) );
  INVX3 U44414 ( .A(n42622), .Y(n42616) );
  INVX3 U44415 ( .A(n42594), .Y(n42587) );
  NOR2BX1 U44416 ( .AN(n41760), .B(n47834), .Y(n41745) );
  OAI31XL U44417 ( .A0(n9804), .A1(n49517), .A2(n9806), .B0(n9772), .Y(n9802)
         );
  NOR3X1 U44418 ( .A(n10102), .B(n10101), .C(n10098), .Y(n24722) );
  NOR2X1 U44419 ( .A(net151299), .B(net171318), .Y(n24712) );
  NOR2X1 U44420 ( .A(net151304), .B(n10301), .Y(n24711) );
  NAND4BX1 U44421 ( .AN(n10066), .B(net168849), .C(n10064), .D(n24685), .Y(
        n9812) );
  NOR2X1 U44422 ( .A(n10067), .B(n10063), .Y(n24685) );
  OAI211X1 U44423 ( .A0(n9865), .A1(n41745), .B0(n9799), .C0(n41758), .Y(n9864) );
  OR2X1 U44424 ( .A(n41746), .B(n41747), .Y(n9819) );
  OR4X1 U44425 ( .A(net171297), .B(net171270), .C(net171294), .D(net151380),
        .Y(n41746) );
  NAND4X1 U44426 ( .A(net259677), .B(n10434), .C(n10436), .D(n10292), .Y(
        n41747) );
  AND2X2 U44427 ( .A(n10336), .B(n37470), .Y(n24678) );
  CLKINVX1 U44428 ( .A(n9747), .Y(net171523) );
  NOR2X1 U44429 ( .A(n45523), .B(n45522), .Y(n45526) );
  NOR4X1 U44430 ( .A(n9763), .B(n9846), .C(n9787), .D(n9788), .Y(n45525) );
  NOR2BX1 U44431 ( .AN(n9845), .B(n50104), .Y(n45524) );
  NAND4X1 U44432 ( .A(n10387), .B(n10385), .C(net151347), .D(n24717), .Y(n9938) );
  NAND4X1 U44433 ( .A(n11543), .B(n11544), .C(n11549), .D(n11550), .Y(n10062)
         );
  NOR2X1 U44434 ( .A(net151275), .B(n10331), .Y(n24680) );
  NAND4BX1 U44435 ( .AN(net210426), .B(n10128), .C(n37125), .D(n41743), .Y(
        n47839) );
  NAND4X1 U44436 ( .A(n11594), .B(n11595), .C(n40418), .D(n40422), .Y(n10073)
         );
  NAND4X1 U44437 ( .A(n12433), .B(net260376), .C(n40415), .D(n40411), .Y(
        n10072) );
  NAND3X1 U44438 ( .A(n10134), .B(net151812), .C(net151819), .Y(n9945) );
  OAI21XL U44439 ( .A0(n9934), .A1(n9794), .B0(n9935), .Y(n9933) );
  AOI211X1 U44440 ( .A0(n49496), .A1(n9937), .B0(n9938), .C0(n9939), .Y(n9934)
         );
  CLKINVX1 U44441 ( .A(n47839), .Y(n49496) );
  OAI31XL U44442 ( .A0(net210390), .A1(n47840), .A2(net210392), .B0(n41750),
        .Y(n9937) );
  CLKINVX1 U44443 ( .A(n9798), .Y(n50090) );
  CLKINVX1 U44444 ( .A(n9908), .Y(n49517) );
  CLKINVX1 U44445 ( .A(n9862), .Y(n50084) );
  NOR2X1 U44446 ( .A(net151349), .B(n10419), .Y(n24718) );
  NAND2X1 U44447 ( .A(n9851), .B(n9958), .Y(n45523) );
  CLKINVX1 U44448 ( .A(n9841), .Y(n49521) );
  CLKINVX1 U44449 ( .A(n9844), .Y(n50111) );
  CLKINVX1 U44450 ( .A(n9847), .Y(n45522) );
  CLKINVX1 U44451 ( .A(n9707), .Y(n50087) );
  INVX3 U44452 ( .A(n41789), .Y(n43040) );
  CLKBUFX3 U44453 ( .A(n9719), .Y(n43044) );
  INVX3 U44454 ( .A(n41789), .Y(n43039) );
  INVX3 U44455 ( .A(n41218), .Y(n42673) );
  NOR2X1 U44456 ( .A(n41748), .B(n41749), .Y(n10076) );
  OR4X1 U44457 ( .A(net171151), .B(net171158), .C(net151283), .D(net151279),
        .Y(n41748) );
  NAND4X1 U44458 ( .A(net259653), .B(net259649), .C(n39470), .D(n39444), .Y(
        n41749) );
  NOR2X1 U44459 ( .A(n47816), .B(n47815), .Y(n41750) );
  CLKINVX1 U44460 ( .A(n9806), .Y(n50094) );
  INVX3 U44461 ( .A(n41790), .Y(n43042) );
  OA21X2 U44462 ( .A0(n19522), .A1(n19487), .B0(n50142), .Y(n19492) );
  NAND2BX2 U44463 ( .AN(n19487), .B(n19411), .Y(n19456) );
  OA21X2 U44464 ( .A0(n19411), .A1(n19487), .B0(n50142), .Y(n19457) );
  INVX3 U44465 ( .A(n19450), .Y(n50128) );
  OAI31XL U44466 ( .A0(n50136), .A1(n19411), .A2(n19412), .B0(n50142), .Y(
        n19450) );
  CLKINVX1 U44467 ( .A(n19449), .Y(n50136) );
  NOR4X1 U44468 ( .A(n49520), .B(n45522), .C(n9787), .D(n9788), .Y(n9784) );
  CLKINVX1 U44469 ( .A(n9958), .Y(n49520) );
  CLKINVX1 U44470 ( .A(n50104), .Y(n49499) );
  AND2X2 U44471 ( .A(n10129), .B(net260527), .Y(n9942) );
  CLKINVX1 U44472 ( .A(n9797), .Y(n50105) );
  CLKINVX1 U44473 ( .A(n9871), .Y(n50092) );
  OAI21X2 U44474 ( .A0(n19281), .A1(n19238), .B0(n50142), .Y(n19247) );
  NAND2X2 U44475 ( .A(n19449), .B(n19411), .Y(n19419) );
  NAND2X2 U44476 ( .A(n19449), .B(n19412), .Y(n19417) );
  NOR2X2 U44477 ( .A(n50129), .B(n50146), .Y(n19411) );
  CLKINVX2 U44478 ( .A(n37520), .Y(n50131) );
  AND2X2 U44479 ( .A(n32368), .B(n50138), .Y(n19187) );
  CLKINVX3 U44480 ( .A(n37530), .Y(n50130) );
  NOR2X1 U44481 ( .A(n19412), .B(n19281), .Y(n19336) );
  INVX3 U44482 ( .A(n42734), .Y(n42732) );
  CLKINVX1 U44483 ( .A(net221992), .Y(net221988) );
  CLKBUFX3 U44484 ( .A(n42449), .Y(n42413) );
  CLKBUFX3 U44485 ( .A(n42449), .Y(n42414) );
  CLKBUFX3 U44486 ( .A(n42449), .Y(n42415) );
  CLKBUFX3 U44487 ( .A(n42448), .Y(n42416) );
  CLKBUFX3 U44488 ( .A(n42448), .Y(n42417) );
  CLKBUFX3 U44489 ( .A(n42448), .Y(n42418) );
  CLKBUFX3 U44490 ( .A(n42447), .Y(n42419) );
  CLKBUFX3 U44491 ( .A(n42447), .Y(n42420) );
  CLKBUFX3 U44492 ( .A(n42447), .Y(n42421) );
  CLKBUFX3 U44493 ( .A(n42445), .Y(n42422) );
  CLKBUFX3 U44494 ( .A(n42445), .Y(n42423) );
  CLKBUFX3 U44495 ( .A(n42445), .Y(n42424) );
  CLKBUFX3 U44496 ( .A(n42444), .Y(n42425) );
  CLKBUFX3 U44497 ( .A(n42443), .Y(n42426) );
  CLKBUFX3 U44498 ( .A(n42442), .Y(n42427) );
  CLKBUFX3 U44499 ( .A(n42441), .Y(n42428) );
  CLKBUFX3 U44500 ( .A(n42441), .Y(n42429) );
  CLKBUFX3 U44501 ( .A(n42440), .Y(n42430) );
  CLKBUFX3 U44502 ( .A(n42440), .Y(n42431) );
  CLKBUFX3 U44503 ( .A(n42439), .Y(n42432) );
  CLKBUFX3 U44504 ( .A(n42438), .Y(n42433) );
  CLKBUFX3 U44505 ( .A(n42437), .Y(n42434) );
  CLKBUFX3 U44506 ( .A(n42437), .Y(n42435) );
  NOR4X1 U44507 ( .A(n27602), .B(n27603), .C(n27604), .D(n27605), .Y(net215466) );
  NOR4X1 U44508 ( .A(n27606), .B(n27607), .C(n27608), .D(n27609), .Y(net215467) );
  NOR4X1 U44509 ( .A(n27297), .B(n27298), .C(n27299), .D(n27300), .Y(net215348) );
  NOR4X1 U44510 ( .A(n27301), .B(n27302), .C(n27303), .D(n27304), .Y(net215349) );
  NOR4X1 U44511 ( .A(n27237), .B(n27238), .C(n27239), .D(n27240), .Y(net215402) );
  NOR4X1 U44512 ( .A(n27241), .B(n27242), .C(n27243), .D(n27244), .Y(net215403) );
  NOR4X1 U44513 ( .A(n27245), .B(n27246), .C(n27247), .D(n27248), .Y(net215404) );
  NOR4X1 U44514 ( .A(n27542), .B(n27543), .C(n27544), .D(n27545), .Y(net215430) );
  NOR4X1 U44515 ( .A(n27512), .B(n27513), .C(n27514), .D(n27515), .Y(net215421) );
  NOR4X1 U44516 ( .A(n27207), .B(n27208), .C(n27209), .D(n27210), .Y(net215375) );
  NOR4X1 U44517 ( .A(n27211), .B(n27212), .C(n27213), .D(n27214), .Y(net215376) );
  NOR4X1 U44518 ( .A(n27215), .B(n27216), .C(n27217), .D(n27218), .Y(net215377) );
  NOR4X1 U44519 ( .A(n27388), .B(n27389), .C(n27390), .D(n27391), .Y(net215438) );
  NOR4X1 U44520 ( .A(n27392), .B(n27393), .C(n27394), .D(n27395), .Y(net215439) );
  NOR4X1 U44521 ( .A(n27418), .B(n27419), .C(n27420), .D(n27421), .Y(n44181)
         );
  NOR4X1 U44522 ( .A(n27422), .B(n27423), .C(n27424), .D(n27425), .Y(n44180)
         );
  NOR4X1 U44523 ( .A(n27426), .B(n27427), .C(n27428), .D(n27429), .Y(n44179)
         );
  NOR4X1 U44524 ( .A(n28019), .B(n28020), .C(n28021), .D(n28022), .Y(net215818) );
  NOR4X1 U44525 ( .A(n28023), .B(n28024), .C(n28025), .D(n28026), .Y(net215819) );
  NOR4X1 U44526 ( .A(n28031), .B(n28032), .C(n28033), .D(n28034), .Y(net215821) );
  NOR4X1 U44527 ( .A(n27357), .B(n27358), .C(n27359), .D(n27360), .Y(net215366) );
  NOR4X1 U44528 ( .A(n27361), .B(n27362), .C(n27363), .D(n27364), .Y(net215367) );
  NOR4X1 U44529 ( .A(n27147), .B(n27148), .C(n27149), .D(n27150), .Y(net215386) );
  NOR4X1 U44530 ( .A(n27151), .B(n27152), .C(n27153), .D(n27154), .Y(net215387) );
  NOR4X1 U44531 ( .A(n27267), .B(n27268), .C(n27269), .D(n27270), .Y(n44201)
         );
  NOR4X1 U44532 ( .A(n27271), .B(n27272), .C(n27273), .D(n27274), .Y(n44200)
         );
  NOR4X1 U44533 ( .A(n27275), .B(n27276), .C(n27277), .D(n27278), .Y(n44199)
         );
  NOR4X1 U44534 ( .A(n27693), .B(n27694), .C(n27695), .D(n27696), .Y(n43836)
         );
  NOR4X1 U44535 ( .A(n27697), .B(n27698), .C(n27699), .D(n27700), .Y(n43835)
         );
  NOR4X1 U44536 ( .A(n27989), .B(n27990), .C(n27991), .D(n27992), .Y(n43828)
         );
  NOR4X1 U44537 ( .A(n27993), .B(n27994), .C(n27995), .D(n27996), .Y(n43827)
         );
  NOR4X1 U44538 ( .A(n27997), .B(n27998), .C(n27999), .D(n28000), .Y(n43826)
         );
  NOR4X1 U44539 ( .A(n27568), .B(n27569), .C(n27570), .D(n27571), .Y(n44172)
         );
  NOR4X1 U44540 ( .A(n27572), .B(n27573), .C(n27574), .D(n27575), .Y(n44171)
         );
  NOR4X1 U44541 ( .A(n27482), .B(n27483), .C(n27484), .D(n27485), .Y(n44577)
         );
  NOR4X1 U44542 ( .A(n27486), .B(n27487), .C(n27488), .D(n27489), .Y(n44576)
         );
  NOR4X1 U44543 ( .A(n29222), .B(n29223), .C(n29224), .D(n29225), .Y(n43581)
         );
  NOR4X1 U44544 ( .A(n29234), .B(n29235), .C(n29236), .D(n29237), .Y(n43578)
         );
  NOR4X1 U44545 ( .A(n28079), .B(n28080), .C(n28081), .D(n28082), .Y(n43817)
         );
  NOR4X1 U44546 ( .A(n27335), .B(n27336), .C(n27337), .D(n27338), .Y(n44225)
         );
  NOR4X1 U44547 ( .A(n27452), .B(n27453), .C(n27454), .D(n27455), .Y(n44574)
         );
  NOR4X1 U44548 ( .A(n27456), .B(n27457), .C(n27458), .D(n27459), .Y(n44573)
         );
  CLKINVX1 U44549 ( .A(n45530), .Y(n48291) );
  NAND4X1 U44550 ( .A(n46568), .B(n46567), .C(n46566), .D(n46565), .Y(n46575)
         );
  NOR2X1 U44551 ( .A(n45048), .B(n45047), .Y(n45053) );
  NOR2X1 U44552 ( .A(n45050), .B(n45049), .Y(n45051) );
  CLKINVX1 U44553 ( .A(net210492), .Y(net210690) );
  NOR2BX1 U44554 ( .AN(net209572), .B(net209570), .Y(n47747) );
  NOR2X1 U44555 ( .A(net209591), .B(net209582), .Y(n47739) );
  NOR2BX1 U44556 ( .AN(net209595), .B(n39479), .Y(n47744) );
  NAND2X1 U44557 ( .A(n48326), .B(n48325), .Y(net210646) );
  NAND2X1 U44558 ( .A(n48289), .B(n48334), .Y(net210639) );
  AND2X2 U44559 ( .A(n48145), .B(n48146), .Y(net234998) );
  CLKINVX1 U44560 ( .A(net210669), .Y(net209633) );
  CLKBUFX3 U44561 ( .A(n42574), .Y(n42570) );
  CLKINVX1 U44562 ( .A(n41630), .Y(n42574) );
  NOR2X1 U44563 ( .A(net210667), .B(net210668), .Y(n47735) );
  CLKBUFX3 U44564 ( .A(n42650), .Y(n42646) );
  NOR4X1 U44565 ( .A(n29342), .B(n29343), .C(n29344), .D(n29345), .Y(net216043) );
  NOR4X1 U44566 ( .A(n29346), .B(n29347), .C(n29348), .D(n29349), .Y(net216044) );
  NOR4X1 U44567 ( .A(n29354), .B(n29355), .C(n29356), .D(n29357), .Y(net216046) );
  NOR4X1 U44568 ( .A(n26815), .B(n26816), .C(n26817), .D(n26818), .Y(net215209) );
  NOR4X1 U44569 ( .A(n29105), .B(n29106), .C(n29107), .D(n29108), .Y(n43647)
         );
  NOR4X1 U44570 ( .A(n29113), .B(n29114), .C(n29115), .D(n29116), .Y(n43645)
         );
  NOR4X1 U44571 ( .A(n29372), .B(n29373), .C(n29374), .D(n29375), .Y(n43572)
         );
  NOR4X1 U44572 ( .A(n26845), .B(n26846), .C(n26847), .D(n26848), .Y(n44312)
         );
  NOR4X1 U44573 ( .A(n26849), .B(n26850), .C(n26851), .D(n26852), .Y(n44311)
         );
  NOR4X1 U44574 ( .A(n27086), .B(n27087), .C(n27088), .D(n27089), .Y(net215312) );
  NOR4X1 U44575 ( .A(n27090), .B(n27091), .C(n27092), .D(n27093), .Y(net215313) );
  NOR4X1 U44576 ( .A(n29282), .B(n29283), .C(n29284), .D(n29285), .Y(net216025) );
  NOR4X1 U44577 ( .A(n29414), .B(n29415), .C(n29416), .D(n29417), .Y(net216138) );
  NAND4X2 U44578 ( .A(n44271), .B(n44270), .C(n44269), .D(n44268), .Y(n11733)
         );
  NOR4X1 U44579 ( .A(n26996), .B(n26997), .C(n26998), .D(n26999), .Y(n44271)
         );
  NOR4X1 U44580 ( .A(n27000), .B(n27001), .C(n27002), .D(n27003), .Y(n44270)
         );
  NOR4X1 U44581 ( .A(n27004), .B(n27005), .C(n27006), .D(n27007), .Y(n44269)
         );
  NOR4X1 U44582 ( .A(n26966), .B(n26967), .C(n26968), .D(n26969), .Y(net215305) );
  NOR4X1 U44583 ( .A(n26970), .B(n26971), .C(n26972), .D(n26973), .Y(net215306) );
  NOR4X1 U44584 ( .A(n26766), .B(n26764), .C(n26763), .D(n26765), .Y(n44600)
         );
  NOR4X1 U44585 ( .A(n29011), .B(n29012), .C(n29013), .D(n29014), .Y(n43670)
         );
  NOR4X1 U44586 ( .A(n29015), .B(n29016), .C(n29017), .D(n29018), .Y(n43669)
         );
  NOR4X1 U44587 ( .A(n26906), .B(n26907), .C(n26908), .D(n26909), .Y(net215276) );
  NOR4X1 U44588 ( .A(n26910), .B(n26911), .C(n26912), .D(n26913), .Y(net215277) );
  NOR4X1 U44589 ( .A(n26729), .B(n26730), .C(n26731), .D(n26732), .Y(n44605)
         );
  NOR4X1 U44590 ( .A(n26733), .B(n26734), .C(n26735), .D(n26736), .Y(n44604)
         );
  NOR4X1 U44591 ( .A(n26936), .B(n26937), .C(n26938), .D(n26939), .Y(net215294) );
  NOR4X1 U44592 ( .A(n26940), .B(n26941), .C(n26942), .D(n26943), .Y(net215295) );
  NOR4X1 U44593 ( .A(n29075), .B(n29076), .C(n29077), .D(n29078), .Y(n43655)
         );
  NOR4X1 U44594 ( .A(n29083), .B(n29084), .C(n29085), .D(n29086), .Y(n43653)
         );
  NOR4X1 U44595 ( .A(n26785), .B(n26786), .C(n26787), .D(n26788), .Y(n44281)
         );
  NOR4X1 U44596 ( .A(n29462), .B(n29463), .C(n29464), .D(n29465), .Y(n43549)
         );
  NOR4X1 U44597 ( .A(n29466), .B(n29467), .C(n29468), .D(n29469), .Y(n43548)
         );
  NOR4X1 U44598 ( .A(n26699), .B(n26700), .C(n26701), .D(n26702), .Y(n44609)
         );
  NOR4X1 U44599 ( .A(n26703), .B(n26704), .C(n26705), .D(n26706), .Y(n44608)
         );
  NOR4X1 U44600 ( .A(n29196), .B(n29197), .C(n29198), .D(n29199), .Y(n43589)
         );
  NOR4X1 U44601 ( .A(n29204), .B(n29205), .C(n29206), .D(n29207), .Y(n43587)
         );
  NOR4X1 U44602 ( .A(n29045), .B(n29046), .C(n29047), .D(n29048), .Y(n43663)
         );
  NOR4X1 U44603 ( .A(n29053), .B(n29054), .C(n29055), .D(n29056), .Y(n43661)
         );
  NOR4X1 U44604 ( .A(n27026), .B(n27027), .C(n27028), .D(n27029), .Y(n44246)
         );
  NOR4X1 U44605 ( .A(n27030), .B(n27031), .C(n27032), .D(n27033), .Y(n44245)
         );
  NOR4X1 U44606 ( .A(n27116), .B(n27117), .C(n27118), .D(n27119), .Y(n44255)
         );
  NOR4X1 U44607 ( .A(n27120), .B(n27121), .C(n27122), .D(n27123), .Y(n44254)
         );
  NOR4X1 U44608 ( .A(n27124), .B(n27125), .C(n27126), .D(n27127), .Y(n44253)
         );
  NOR4X1 U44609 ( .A(n29312), .B(n29313), .C(n29314), .D(n29315), .Y(n43638)
         );
  NOR4X1 U44610 ( .A(n29316), .B(n29317), .C(n29318), .D(n29319), .Y(n43637)
         );
  NOR4X1 U44611 ( .A(n29324), .B(n29325), .C(n29326), .D(n29327), .Y(n43635)
         );
  NOR4X1 U44612 ( .A(n29252), .B(n29253), .C(n29254), .D(n29255), .Y(n43628)
         );
  NOR4X1 U44613 ( .A(n29256), .B(n29257), .C(n29258), .D(n29259), .Y(n43627)
         );
  NAND4X1 U44614 ( .A(n44597), .B(n44596), .C(n44595), .D(n44594), .Y(n12538)
         );
  NOR4X1 U44615 ( .A(n29139), .B(n29136), .C(n29137), .D(n29138), .Y(n44596)
         );
  NOR4X1 U44616 ( .A(n29147), .B(n29145), .C(n29144), .D(n29146), .Y(n44594)
         );
  NAND4X1 U44617 ( .A(n44593), .B(n44592), .C(n44591), .D(n44590), .Y(n11763)
         );
  NOR4X1 U44618 ( .A(n29169), .B(n29166), .C(n29167), .D(n29168), .Y(n44592)
         );
  NOR4X1 U44619 ( .A(n29165), .B(n29163), .C(n29162), .D(n29164), .Y(n44593)
         );
  NOR4X1 U44620 ( .A(n29174), .B(n29175), .C(n29177), .D(n29176), .Y(n44590)
         );
  NOR4X1 U44621 ( .A(n29143), .B(n29140), .C(n29141), .D(n29142), .Y(n44595)
         );
  NAND3X1 U44622 ( .A(n44297), .B(n44296), .C(n44295), .Y(n44298) );
  NOR2X1 U44623 ( .A(n26746), .B(n26769), .Y(n44297) );
  NOR3X1 U44624 ( .A(n26770), .B(n26762), .C(n26758), .Y(n44295) );
  NOR2X1 U44625 ( .A(n48315), .B(n48314), .Y(n48316) );
  NOR3X1 U44626 ( .A(n48340), .B(n48339), .C(n48338), .Y(n48341) );
  NAND2BX1 U44627 ( .AN(n48237), .B(n48236), .Y(n48238) );
  OR3X2 U44628 ( .A(n41753), .B(n29165), .C(n29162), .Y(n43602) );
  OR2X1 U44629 ( .A(n29177), .B(n29169), .Y(n41753) );
  OR3X2 U44630 ( .A(n41754), .B(n29135), .C(n29138), .Y(n43619) );
  OR3X2 U44631 ( .A(n26763), .B(n26747), .C(n26761), .Y(n44288) );
  OR2X1 U44632 ( .A(n41755), .B(n29142), .Y(n43618) );
  OR2X1 U44633 ( .A(n41756), .B(n29168), .Y(n43605) );
  CLKINVX1 U44634 ( .A(n29134), .Y(n43612) );
  CLKINVX1 U44635 ( .A(n29166), .Y(n43599) );
  CLKINVX1 U44636 ( .A(n29144), .Y(n43613) );
  CLKBUFX3 U44637 ( .A(n42692), .Y(n42690) );
  NOR4X1 U44638 ( .A(n28294), .B(n28295), .C(n28296), .D(n28297), .Y(n43753)
         );
  NAND4X2 U44639 ( .A(n44502), .B(n44501), .C(n44500), .D(n44499), .Y(n11711)
         );
  NOR4X1 U44640 ( .A(n24952), .B(n24953), .C(n24954), .D(n24955), .Y(n44502)
         );
  NOR4X1 U44641 ( .A(n24956), .B(n24957), .C(n24958), .D(n24959), .Y(n44501)
         );
  NOR4X1 U44642 ( .A(n24960), .B(n24961), .C(n24962), .D(n24963), .Y(n44500)
         );
  NOR4X1 U44643 ( .A(n28200), .B(n28201), .C(n28202), .D(n28203), .Y(n43781)
         );
  NOR4X1 U44644 ( .A(n28204), .B(n28205), .C(n28206), .D(n28207), .Y(n43780)
         );
  NOR4X1 U44645 ( .A(n28530), .B(n28531), .C(n28532), .D(n28533), .Y(n43690)
         );
  NOR4X1 U44646 ( .A(n28534), .B(n28535), .C(n28536), .D(n28537), .Y(n43689)
         );
  NOR4X1 U44647 ( .A(n28350), .B(n28351), .C(n28352), .D(n28353), .Y(n43744)
         );
  NOR4X1 U44648 ( .A(n28354), .B(n28355), .C(n28356), .D(n28357), .Y(n43743)
         );
  NOR4X1 U44649 ( .A(n28362), .B(n28363), .C(n28364), .D(n28365), .Y(n43741)
         );
  NOR4X1 U44650 ( .A(n28110), .B(n28111), .C(n28112), .D(n28113), .Y(n43808)
         );
  NOR4X1 U44651 ( .A(n24742), .B(n24743), .C(n24744), .D(n24745), .Y(n44564)
         );
  NOR4X1 U44652 ( .A(n24746), .B(n24747), .C(n24748), .D(n24749), .Y(n44563)
         );
  NOR4X1 U44653 ( .A(n24750), .B(n24751), .C(n24752), .D(n24753), .Y(n44562)
         );
  NOR4X1 U44654 ( .A(n28500), .B(n28501), .C(n28502), .D(n28503), .Y(n43699)
         );
  NOR4X1 U44655 ( .A(n28504), .B(n28505), .C(n28506), .D(n28507), .Y(n43698)
         );
  NOR4X1 U44656 ( .A(n31179), .B(n31180), .C(n31181), .D(n31182), .Y(n43329)
         );
  NOR4X1 U44657 ( .A(n31183), .B(n31184), .C(n31185), .D(n31186), .Y(n43328)
         );
  NOR4X1 U44658 ( .A(n31191), .B(n31192), .C(n31193), .D(n31194), .Y(n43326)
         );
  NOR4X1 U44659 ( .A(n28320), .B(n28321), .C(n28322), .D(n28323), .Y(n43749)
         );
  NOR4X1 U44660 ( .A(n28324), .B(n28325), .C(n28326), .D(n28327), .Y(n43748)
         );
  NOR4X1 U44661 ( .A(n28332), .B(n28333), .C(n28334), .D(n28335), .Y(n43746)
         );
  NOR4X1 U44662 ( .A(n24892), .B(n24893), .C(n24894), .D(n24895), .Y(n44520)
         );
  NOR4X1 U44663 ( .A(n24896), .B(n24897), .C(n24898), .D(n24899), .Y(n44519)
         );
  NOR4X1 U44664 ( .A(n24900), .B(n24901), .C(n24902), .D(n24903), .Y(n44518)
         );
  NOR4X1 U44665 ( .A(n28410), .B(n28411), .C(n28412), .D(n28413), .Y(n43726)
         );
  NOR4X1 U44666 ( .A(n28414), .B(n28415), .C(n28416), .D(n28417), .Y(n43725)
         );
  NOR4X1 U44667 ( .A(n28422), .B(n28423), .C(n28424), .D(n28425), .Y(n43723)
         );
  NOR4X1 U44668 ( .A(n28170), .B(n28171), .C(n28172), .D(n28173), .Y(n43790)
         );
  NOR4X1 U44669 ( .A(n28174), .B(n28175), .C(n28176), .D(n28177), .Y(n43789)
         );
  NOR4X1 U44670 ( .A(n28560), .B(n28561), .C(n28562), .D(n28563), .Y(n43679)
         );
  NOR4X1 U44671 ( .A(n28564), .B(n28565), .C(n28566), .D(n28567), .Y(n43678)
         );
  NOR4X1 U44672 ( .A(n28572), .B(n28573), .C(n28574), .D(n28575), .Y(n43680)
         );
  NOR4X1 U44673 ( .A(n28440), .B(n28441), .C(n28442), .D(n28443), .Y(n43717)
         );
  NOR4X1 U44674 ( .A(n28444), .B(n28445), .C(n28446), .D(n28447), .Y(n43716)
         );
  NOR4X1 U44675 ( .A(n28470), .B(n28471), .C(n28472), .D(n28473), .Y(n43708)
         );
  NOR4X1 U44676 ( .A(n28474), .B(n28475), .C(n28476), .D(n28477), .Y(n43707)
         );
  NOR4X1 U44677 ( .A(n28482), .B(n28483), .C(n28484), .D(n28485), .Y(n43705)
         );
  NOR4X1 U44678 ( .A(n24930), .B(n24931), .C(n24932), .D(n24933), .Y(n44509)
         );
  NOR4X1 U44679 ( .A(n24840), .B(n24841), .C(n24842), .D(n24843), .Y(n44537)
         );
  NOR4X1 U44680 ( .A(n24844), .B(n24845), .C(n24846), .D(n24847), .Y(n44536)
         );
  NOR4X1 U44681 ( .A(n24832), .B(n24833), .C(n24834), .D(n24835), .Y(n44535)
         );
  NOR4X1 U44682 ( .A(n24780), .B(n24781), .C(n24782), .D(n24783), .Y(n44553)
         );
  NOR4X1 U44683 ( .A(n28230), .B(n28231), .C(n28232), .D(n28233), .Y(n43772)
         );
  NOR4X1 U44684 ( .A(n28234), .B(n28235), .C(n28236), .D(n28237), .Y(n43771)
         );
  NOR4X1 U44685 ( .A(n28242), .B(n28243), .C(n28244), .D(n28245), .Y(n43769)
         );
  NOR4X1 U44686 ( .A(n31269), .B(n31270), .C(n31271), .D(n31272), .Y(n43302)
         );
  NOR4X1 U44687 ( .A(n31273), .B(n31274), .C(n31275), .D(n31276), .Y(n43301)
         );
  NOR4X1 U44688 ( .A(n31281), .B(n31282), .C(n31283), .D(n31284), .Y(n43299)
         );
  NOR4X1 U44689 ( .A(n25192), .B(n25193), .C(n25194), .D(n25195), .Y(n44426)
         );
  NOR4X1 U44690 ( .A(n25200), .B(n25201), .C(n25202), .D(n25203), .Y(n44424)
         );
  NOR4X1 U44691 ( .A(n25012), .B(n25013), .C(n25014), .D(n25015), .Y(n44488)
         );
  NOR4X1 U44692 ( .A(n25016), .B(n25017), .C(n25018), .D(n25019), .Y(n44487)
         );
  NOR4X1 U44693 ( .A(n25020), .B(n25021), .C(n25022), .D(n25023), .Y(n44486)
         );
  NOR4X1 U44694 ( .A(n31629), .B(n31630), .C(n31631), .D(n31632), .Y(n43195)
         );
  NOR4X1 U44695 ( .A(n31633), .B(n31634), .C(n31635), .D(n31636), .Y(n43194)
         );
  NOR4X1 U44696 ( .A(n31641), .B(n31642), .C(n31643), .D(n31644), .Y(n43192)
         );
  NOR4X1 U44697 ( .A(n28260), .B(n28261), .C(n28262), .D(n28263), .Y(n43763)
         );
  NOR4X1 U44698 ( .A(n28264), .B(n28265), .C(n28266), .D(n28267), .Y(n43762)
         );
  NOR4X1 U44699 ( .A(n24866), .B(n24867), .C(n24868), .D(n24869), .Y(n44528)
         );
  NOR4X1 U44700 ( .A(n24870), .B(n24871), .C(n24872), .D(n24873), .Y(n44527)
         );
  NOR4X1 U44701 ( .A(n31393), .B(n31394), .C(n31395), .D(n31396), .Y(n43266)
         );
  NOR4X1 U44702 ( .A(n31401), .B(n31402), .C(n31403), .D(n31404), .Y(n43264)
         );
  NOR4X1 U44703 ( .A(n25166), .B(n25167), .C(n25168), .D(n25169), .Y(n44434)
         );
  NOR4X1 U44704 ( .A(n25170), .B(n25171), .C(n25172), .D(n25173), .Y(n44433)
         );
  NOR4X1 U44705 ( .A(n27056), .B(n27057), .C(n27058), .D(n27059), .Y(n44237)
         );
  NOR4X1 U44706 ( .A(n27060), .B(n27061), .C(n27062), .D(n27063), .Y(n44236)
         );
  NOR4X1 U44707 ( .A(n27064), .B(n27065), .C(n27066), .D(n27067), .Y(n44235)
         );
  NOR4X1 U44708 ( .A(n25042), .B(n25043), .C(n25044), .D(n25045), .Y(n44479)
         );
  NOR4X1 U44709 ( .A(n25046), .B(n25047), .C(n25048), .D(n25049), .Y(n44478)
         );
  NOR4X1 U44710 ( .A(n25050), .B(n25051), .C(n25052), .D(n25053), .Y(n44477)
         );
  NOR4X1 U44711 ( .A(n31569), .B(n31570), .C(n31571), .D(n31572), .Y(n43213)
         );
  NOR4X1 U44712 ( .A(n31573), .B(n31574), .C(n31575), .D(n31576), .Y(n43212)
         );
  NOR4X1 U44713 ( .A(n31581), .B(n31582), .C(n31583), .D(n31584), .Y(n43210)
         );
  NOR4X1 U44714 ( .A(n28380), .B(n28381), .C(n28382), .D(n28383), .Y(n43735)
         );
  NOR4X1 U44715 ( .A(n28384), .B(n28385), .C(n28386), .D(n28387), .Y(n43734)
         );
  CLKINVX1 U44716 ( .A(n12063), .Y(net171252) );
  NOR2X1 U44717 ( .A(n25114), .B(n25115), .Y(n44456) );
  NOR2X1 U44718 ( .A(n25110), .B(n25111), .Y(n44458) );
  NOR4X1 U44719 ( .A(n25072), .B(n25073), .C(n25074), .D(n25075), .Y(n44470)
         );
  NOR4X1 U44720 ( .A(n25076), .B(n25077), .C(n25078), .D(n25079), .Y(n44469)
         );
  NOR4X1 U44721 ( .A(n25080), .B(n25081), .C(n25082), .D(n25083), .Y(n44468)
         );
  NOR4X1 U44722 ( .A(n31599), .B(n31600), .C(n31601), .D(n31602), .Y(n43204)
         );
  NOR4X1 U44723 ( .A(n31603), .B(n31604), .C(n31605), .D(n31606), .Y(n43203)
         );
  NOR4X1 U44724 ( .A(n31611), .B(n31612), .C(n31613), .D(n31614), .Y(n43201)
         );
  NOR4X1 U44725 ( .A(n31359), .B(n31360), .C(n31361), .D(n31362), .Y(n43275)
         );
  NOR4X1 U44726 ( .A(n31363), .B(n31364), .C(n31365), .D(n31366), .Y(n43274)
         );
  NOR4X1 U44727 ( .A(n31371), .B(n31372), .C(n31373), .D(n31374), .Y(n43272)
         );
  CLKINVX1 U44728 ( .A(n48319), .Y(n48327) );
  NOR4X1 U44729 ( .A(n24982), .B(n24983), .C(n24984), .D(n24985), .Y(n44493)
         );
  NOR4X1 U44730 ( .A(n24986), .B(n24987), .C(n24988), .D(n24989), .Y(n44492)
         );
  NOR4X1 U44731 ( .A(n24990), .B(n24991), .C(n24992), .D(n24993), .Y(n44491)
         );
  NAND4X1 U44732 ( .A(n44455), .B(n44454), .C(n44453), .D(n44452), .Y(n44570)
         );
  NOR2X1 U44733 ( .A(n25102), .B(n25103), .Y(n44454) );
  NOR2X1 U44734 ( .A(n25106), .B(n25107), .Y(n44452) );
  NOR2X1 U44735 ( .A(n25104), .B(n25105), .Y(n44455) );
  NOR2X1 U44736 ( .A(n25132), .B(n25133), .Y(n44446) );
  NOR2X1 U44737 ( .A(n25136), .B(n25137), .Y(n44444) );
  NOR2X1 U44738 ( .A(n25134), .B(n25135), .Y(n44447) );
  NOR2X1 U44739 ( .A(n25144), .B(n25145), .Y(n44440) );
  NOR2X1 U44740 ( .A(n25140), .B(n25141), .Y(n44442) );
  NOR2X1 U44741 ( .A(n25142), .B(n25143), .Y(n44443) );
  OAI21XL U44742 ( .A0(n48295), .A1(n48294), .B0(n48293), .Y(n48296) );
  CLKINVX1 U44743 ( .A(n48145), .Y(n48148) );
  CLKINVX1 U44744 ( .A(n48325), .Y(n48331) );
  NOR2X1 U44745 ( .A(n48328), .B(n48327), .Y(n48329) );
  CLKINVX1 U44746 ( .A(net210526), .Y(net210205) );
  NOR2X1 U44747 ( .A(net209591), .B(net209592), .Y(n48321) );
  OA21XL U44748 ( .A0(n48327), .A1(n48320), .B0(net209595), .Y(n41757) );
  NOR2X1 U44749 ( .A(net209280), .B(net209302), .Y(n48456) );
  CLKINVX1 U44750 ( .A(n48326), .Y(n48328) );
  NOR2X1 U44751 ( .A(net151662), .B(net171458), .Y(n11067) );
  NOR4X1 U44752 ( .A(n31239), .B(n31240), .C(n31241), .D(n31242), .Y(n43311)
         );
  NOR4X1 U44753 ( .A(n31243), .B(n31244), .C(n31245), .D(n31246), .Y(n43310)
         );
  NOR4X1 U44754 ( .A(n31251), .B(n31252), .C(n31253), .D(n31254), .Y(n43308)
         );
  NOR4X1 U44755 ( .A(n31672), .B(n31673), .C(n31674), .D(n31675), .Y(net216759) );
  NOR4X1 U44756 ( .A(n31732), .B(n31733), .C(n31734), .D(n31735), .Y(net216750) );
  NOR4X1 U44757 ( .A(n31088), .B(n31089), .C(n31090), .D(n31091), .Y(n43351)
         );
  NOR4X1 U44758 ( .A(n31092), .B(n31093), .C(n31094), .D(n31095), .Y(n43350)
         );
  NOR4X1 U44759 ( .A(n31100), .B(n31101), .C(n31102), .D(n31103), .Y(n43348)
         );
  NOR4X1 U44760 ( .A(n31122), .B(n31123), .C(n31124), .D(n31125), .Y(n43342)
         );
  NOR4X1 U44761 ( .A(n31130), .B(n31131), .C(n31132), .D(n31133), .Y(n43340)
         );
  NOR4X1 U44762 ( .A(n31509), .B(n31510), .C(n31511), .D(n31512), .Y(n43231)
         );
  NOR4X1 U44763 ( .A(n31513), .B(n31514), .C(n31515), .D(n31516), .Y(n43230)
         );
  NOR4X1 U44764 ( .A(n31521), .B(n31522), .C(n31523), .D(n31524), .Y(n43228)
         );
  NOR4X1 U44765 ( .A(n30968), .B(n30969), .C(n30970), .D(n30971), .Y(n43384)
         );
  NOR4X1 U44766 ( .A(n30972), .B(n30973), .C(n30974), .D(n30975), .Y(n43383)
         );
  NOR4X1 U44767 ( .A(n30980), .B(n30981), .C(n30982), .D(n30983), .Y(n43385)
         );
  NOR4X1 U44768 ( .A(n31419), .B(n31420), .C(n31421), .D(n31422), .Y(n43258)
         );
  NOR4X1 U44769 ( .A(n31423), .B(n31424), .C(n31425), .D(n31426), .Y(n43257)
         );
  NOR4X1 U44770 ( .A(n31431), .B(n31432), .C(n31433), .D(n31434), .Y(n43255)
         );
  NOR4X1 U44771 ( .A(n31028), .B(n31029), .C(n31030), .D(n31031), .Y(n43368)
         );
  NOR4X1 U44772 ( .A(n31032), .B(n31033), .C(n31034), .D(n31035), .Y(n43367)
         );
  NOR4X1 U44773 ( .A(n31040), .B(n31041), .C(n31042), .D(n31043), .Y(n43365)
         );
  NOR4X1 U44774 ( .A(n31062), .B(n31063), .C(n31064), .D(n31065), .Y(n43359)
         );
  NOR4X1 U44775 ( .A(n31070), .B(n31071), .C(n31072), .D(n31073), .Y(n43357)
         );
  NOR4X1 U44776 ( .A(n30998), .B(n30999), .C(n31000), .D(n31001), .Y(n43377)
         );
  NOR4X1 U44777 ( .A(n31002), .B(n31003), .C(n31004), .D(n31005), .Y(n43376)
         );
  NOR4X1 U44778 ( .A(n31010), .B(n31011), .C(n31012), .D(n31013), .Y(n43374)
         );
  NOR4X1 U44779 ( .A(n31479), .B(n31480), .C(n31481), .D(n31482), .Y(n43240)
         );
  NOR4X1 U44780 ( .A(n31483), .B(n31484), .C(n31485), .D(n31486), .Y(n43239)
         );
  NOR4X1 U44781 ( .A(n31491), .B(n31492), .C(n31493), .D(n31494), .Y(n43237)
         );
  NOR4X1 U44782 ( .A(n31822), .B(n31823), .C(n31824), .D(n31825), .Y(net214663) );
  NOR4X1 U44783 ( .A(n31148), .B(n31149), .C(n31150), .D(n31151), .Y(net216594) );
  NOR4X1 U44784 ( .A(n31152), .B(n31153), .C(n31154), .D(n31155), .Y(net216595) );
  NOR4X1 U44785 ( .A(n31160), .B(n31161), .C(n31162), .D(n31163), .Y(net216597) );
  NOR4X1 U44786 ( .A(n31870), .B(n31871), .C(n31872), .D(n31873), .Y(n44639)
         );
  NOR4X1 U44787 ( .A(n31874), .B(n31875), .C(n31876), .D(n31877), .Y(n44638)
         );
  NOR4X1 U44788 ( .A(n31882), .B(n31883), .C(n31884), .D(n31885), .Y(n44636)
         );
  NOR4X1 U44789 ( .A(n31329), .B(n31330), .C(n31331), .D(n31332), .Y(n43284)
         );
  NOR4X1 U44790 ( .A(n31333), .B(n31334), .C(n31335), .D(n31336), .Y(n43283)
         );
  NOR4X1 U44791 ( .A(n31341), .B(n31342), .C(n31343), .D(n31344), .Y(n43281)
         );
  NOR4X1 U44792 ( .A(n31750), .B(n31751), .C(n31752), .D(n31753), .Y(n43167)
         );
  NOR4X1 U44793 ( .A(n31754), .B(n31755), .C(n31756), .D(n31757), .Y(n43166)
         );
  NOR4X1 U44794 ( .A(n31762), .B(n31763), .C(n31764), .D(n31765), .Y(n43164)
         );
  NOR4X1 U44795 ( .A(n31449), .B(n31450), .C(n31451), .D(n31452), .Y(n43249)
         );
  NOR4X1 U44796 ( .A(n31453), .B(n31454), .C(n31455), .D(n31456), .Y(n43248)
         );
  NOR4X1 U44797 ( .A(n31461), .B(n31462), .C(n31463), .D(n31464), .Y(n43246)
         );
  NOR4X1 U44798 ( .A(n31690), .B(n31691), .C(n31692), .D(n31693), .Y(n43176)
         );
  NOR4X1 U44799 ( .A(n31694), .B(n31695), .C(n31696), .D(n31697), .Y(n43175)
         );
  NOR4X1 U44800 ( .A(n31702), .B(n31703), .C(n31704), .D(n31705), .Y(n43173)
         );
  NOR4X1 U44801 ( .A(n31780), .B(n31781), .C(n31782), .D(n31783), .Y(n43158)
         );
  NOR4X1 U44802 ( .A(n31784), .B(n31785), .C(n31786), .D(n31787), .Y(n43157)
         );
  NOR4X1 U44803 ( .A(n31792), .B(n31793), .C(n31794), .D(n31795), .Y(n43155)
         );
  NOR4X1 U44804 ( .A(n31209), .B(n31210), .C(n31211), .D(n31212), .Y(n43320)
         );
  NOR4X1 U44805 ( .A(n31213), .B(n31214), .C(n31215), .D(n31216), .Y(n43319)
         );
  NOR4X1 U44806 ( .A(n31221), .B(n31222), .C(n31223), .D(n31224), .Y(n43317)
         );
  NOR4X1 U44807 ( .A(n31840), .B(n31841), .C(n31842), .D(n31843), .Y(n44585)
         );
  NOR4X1 U44808 ( .A(n31844), .B(n31845), .C(n31846), .D(n31847), .Y(n44584)
         );
  NOR4X1 U44809 ( .A(n31852), .B(n31853), .C(n31854), .D(n31855), .Y(n44582)
         );
  NAND2BX1 U44810 ( .AN(n47766), .B(n41762), .Y(net211102) );
  CLKINVX1 U44811 ( .A(net210698), .Y(net214265) );
  CLKINVX1 U44812 ( .A(net210688), .Y(net213824) );
  CLKINVX1 U44813 ( .A(n11046), .Y(net151477) );
  NOR4X1 U44814 ( .A(n30890), .B(n30891), .C(n30892), .D(n30893), .Y(net216471) );
  NOR4X1 U44815 ( .A(n32111), .B(n32112), .C(n32113), .D(n32114), .Y(n43103)
         );
  NOR4X1 U44816 ( .A(n32119), .B(n32120), .C(n32121), .D(n32122), .Y(n43101)
         );
  NOR4X1 U44817 ( .A(n32115), .B(n32116), .C(n32117), .D(n32118), .Y(n43102)
         );
  NOR4X1 U44818 ( .A(n32149), .B(n32150), .C(n32151), .D(n32152), .Y(n43093)
         );
  NOR4X1 U44819 ( .A(n32145), .B(n32146), .C(n32147), .D(n32148), .Y(n43094)
         );
  NOR4X1 U44820 ( .A(n31931), .B(n31932), .C(n31933), .D(n31934), .Y(n43149)
         );
  NOR4X1 U44821 ( .A(n31939), .B(n31940), .C(n31941), .D(n31942), .Y(n43147)
         );
  NOR4X1 U44822 ( .A(n31935), .B(n31936), .C(n31937), .D(n31938), .Y(n43148)
         );
  NOR4X1 U44823 ( .A(n30740), .B(n30741), .C(n30742), .D(n30743), .Y(net216507) );
  NOR4X1 U44824 ( .A(n30770), .B(n30771), .C(n30772), .D(n30773), .Y(net216516) );
  NOR4X1 U44825 ( .A(n31991), .B(n31992), .C(n31993), .D(n31994), .Y(n43135)
         );
  NOR4X1 U44826 ( .A(n31999), .B(n32000), .C(n32001), .D(n32002), .Y(n43133)
         );
  NOR4X1 U44827 ( .A(n31995), .B(n31996), .C(n31997), .D(n31998), .Y(n43134)
         );
  NOR4X1 U44828 ( .A(n30710), .B(n30711), .C(n30712), .D(n30713), .Y(net216498) );
  NOR4X1 U44829 ( .A(n32081), .B(n32082), .C(n32083), .D(n32084), .Y(n43112)
         );
  NOR4X1 U44830 ( .A(n32089), .B(n32090), .C(n32091), .D(n32092), .Y(n43110)
         );
  NOR4X1 U44831 ( .A(n32085), .B(n32086), .C(n32087), .D(n32088), .Y(n43111)
         );
  NOR4X1 U44832 ( .A(n32051), .B(n32052), .C(n32053), .D(n32054), .Y(n43121)
         );
  NOR4X1 U44833 ( .A(n32059), .B(n32060), .C(n32061), .D(n32062), .Y(n43119)
         );
  NOR4X1 U44834 ( .A(n32055), .B(n32056), .C(n32057), .D(n32058), .Y(n43120)
         );
  NOR4X1 U44835 ( .A(n30860), .B(n30861), .C(n30862), .D(n30863), .Y(net216462) );
  NOR4X1 U44836 ( .A(n32291), .B(n32292), .C(n32293), .D(n32294), .Y(n43048)
         );
  NOR4X1 U44837 ( .A(n32299), .B(n32300), .C(n32301), .D(n32302), .Y(n43046)
         );
  NOR4X1 U44838 ( .A(n32295), .B(n32296), .C(n32297), .D(n32298), .Y(n43047)
         );
  NAND4X1 U44839 ( .A(n43140), .B(n43139), .C(n43138), .D(n43137), .Y(n12452)
         );
  NOR4X1 U44840 ( .A(n31961), .B(n31962), .C(n31963), .D(n31964), .Y(n43140)
         );
  NOR4X1 U44841 ( .A(n31969), .B(n31970), .C(n31971), .D(n31972), .Y(n43138)
         );
  NOR4X1 U44842 ( .A(n31965), .B(n31966), .C(n31967), .D(n31968), .Y(n43139)
         );
  NOR4X1 U44843 ( .A(n32201), .B(n32202), .C(n32203), .D(n32204), .Y(n43067)
         );
  NOR4X1 U44844 ( .A(n32209), .B(n32210), .C(n32211), .D(n32212), .Y(n43065)
         );
  NOR4X1 U44845 ( .A(n32205), .B(n32206), .C(n32207), .D(n32208), .Y(n43066)
         );
  NAND4X1 U44846 ( .A(n43076), .B(n43075), .C(n43074), .D(n43073), .Y(n12455)
         );
  NOR4X1 U44847 ( .A(n32351), .B(n32352), .C(n32353), .D(n32354), .Y(n43076)
         );
  NOR4X1 U44848 ( .A(n32359), .B(n32360), .C(n32361), .D(n32362), .Y(n43074)
         );
  NOR4X1 U44849 ( .A(n32355), .B(n32356), .C(n32357), .D(n32358), .Y(n43075)
         );
  NOR4X1 U44850 ( .A(n32171), .B(n32172), .C(n32173), .D(n32174), .Y(n43086)
         );
  NOR4X1 U44851 ( .A(n32179), .B(n32180), .C(n32181), .D(n32182), .Y(n43084)
         );
  NOR4X1 U44852 ( .A(n32175), .B(n32176), .C(n32177), .D(n32178), .Y(n43085)
         );
  NOR4X1 U44853 ( .A(n32231), .B(n32232), .C(n32233), .D(n32234), .Y(n43058)
         );
  NOR4X1 U44854 ( .A(n32239), .B(n32240), .C(n32241), .D(n32242), .Y(n43056)
         );
  NOR4X1 U44855 ( .A(n32235), .B(n32236), .C(n32237), .D(n32238), .Y(n43057)
         );
  NOR4X1 U44856 ( .A(n32021), .B(n32022), .C(n32023), .D(n32024), .Y(n43130)
         );
  NOR4X1 U44857 ( .A(n32029), .B(n32030), .C(n32031), .D(n32032), .Y(n43128)
         );
  NOR4X1 U44858 ( .A(n32025), .B(n32026), .C(n32027), .D(n32028), .Y(n43129)
         );
  NOR4X1 U44859 ( .A(n30938), .B(n30939), .C(n30940), .D(n30941), .Y(n43395)
         );
  NOR4X1 U44860 ( .A(n30942), .B(n30943), .C(n30944), .D(n30945), .Y(n43394)
         );
  NOR4X1 U44861 ( .A(n30950), .B(n30951), .C(n30952), .D(n30953), .Y(n43392)
         );
  NOR4X1 U44862 ( .A(n30788), .B(n30789), .C(n30790), .D(n30791), .Y(n43404)
         );
  NOR4X1 U44863 ( .A(n30792), .B(n30793), .C(n30794), .D(n30795), .Y(n43403)
         );
  NOR4X1 U44864 ( .A(n30800), .B(n30801), .C(n30802), .D(n30803), .Y(n43401)
         );
  NOR4X1 U44865 ( .A(n32321), .B(n32322), .C(n32323), .D(n32324), .Y(n43081)
         );
  NOR4X1 U44866 ( .A(n32325), .B(n32326), .C(n32327), .D(n32328), .Y(n43080)
         );
  NOR4X1 U44867 ( .A(n32333), .B(n32334), .C(n32335), .D(n32336), .Y(n43078)
         );
  NAND4X1 U44868 ( .A(n43053), .B(n43052), .C(n43051), .D(n43050), .Y(
        net214724) );
  NOR4X1 U44869 ( .A(n32261), .B(n32262), .C(n32263), .D(n32264), .Y(n43053)
         );
  NOR4X1 U44870 ( .A(n32265), .B(n32266), .C(n32267), .D(n32268), .Y(n43052)
         );
  NOR4X1 U44871 ( .A(n32269), .B(n32270), .C(n32271), .D(n32272), .Y(n43051)
         );
  NOR4X1 U44872 ( .A(n31901), .B(n31902), .C(n31903), .D(n31904), .Y(n44589)
         );
  NOR4X1 U44873 ( .A(n31909), .B(n31910), .C(n31911), .D(n31912), .Y(n44587)
         );
  NOR4X1 U44874 ( .A(n31905), .B(n31906), .C(n31907), .D(n31908), .Y(n44588)
         );
  NOR2X1 U44875 ( .A(net151494), .B(net151491), .Y(n11019) );
  NAND4BX2 U44876 ( .AN(n46609), .B(n46608), .C(n46607), .D(n46606), .Y(n9747)
         );
  NOR2X1 U44877 ( .A(n10198), .B(n9865), .Y(n46608) );
  NOR2X1 U44878 ( .A(n9797), .B(n9871), .Y(n46607) );
  NAND3X1 U44879 ( .A(n9799), .B(n41745), .C(n41758), .Y(n46609) );
  NOR3BX1 U44880 ( .AN(n9898), .B(n9901), .C(n9900), .Y(n9771) );
  NOR4X1 U44881 ( .A(n30275), .B(n30276), .C(n30277), .D(n30278), .Y(n43485)
         );
  NOR4X1 U44882 ( .A(n30279), .B(n30280), .C(n30281), .D(n30282), .Y(n43484)
         );
  NOR4X1 U44883 ( .A(n30287), .B(n30288), .C(n30289), .D(n30290), .Y(n43482)
         );
  NOR4X1 U44884 ( .A(n26303), .B(n26304), .C(n26305), .D(n26306), .Y(net215119) );
  NOR4X1 U44885 ( .A(n26307), .B(n26308), .C(n26309), .D(n26310), .Y(net215120) );
  NOR4X1 U44886 ( .A(n26311), .B(n26312), .C(n26313), .D(n26314), .Y(net215121) );
  NOR4X1 U44887 ( .A(n25921), .B(n25922), .C(n25923), .D(n25924), .Y(net215004) );
  NOR4X1 U44888 ( .A(n25853), .B(n25854), .C(n25855), .D(n25856), .Y(net215020) );
  NOR4X1 U44889 ( .A(n25857), .B(n25858), .C(n25859), .D(n25860), .Y(net215021) );
  NOR4X1 U44890 ( .A(n25861), .B(n25862), .C(n25863), .D(n25864), .Y(net215022) );
  NOR3BX1 U44891 ( .AN(n9875), .B(n9876), .C(n9877), .Y(n9773) );
  NOR4X1 U44892 ( .A(n29523), .B(n29524), .C(n29525), .D(n29526), .Y(net216180) );
  NOR4X1 U44893 ( .A(n29535), .B(n29536), .C(n29537), .D(n29538), .Y(net216183) );
  AOI211X1 U44894 ( .A0(n10140), .A1(n10141), .B0(n10142), .C0(n10143), .Y(
        n10138) );
  OAI21XL U44895 ( .A0(n10144), .A1(n9954), .B0(n50106), .Y(n10141) );
  AOI211X1 U44896 ( .A0(n9844), .A1(n10149), .B0(n10150), .C0(net171111), .Y(
        n10147) );
  NOR4X1 U44897 ( .A(n9884), .B(n9880), .C(n9885), .D(n21123), .Y(n9772) );
  OR3X2 U44898 ( .A(n9882), .B(n9881), .C(n9886), .Y(n21123) );
  NOR4X1 U44899 ( .A(n30559), .B(n30560), .C(n30561), .D(n30562), .Y(net216444) );
  NOR4X1 U44900 ( .A(n10024), .B(net171548), .C(n10028), .D(n19852), .Y(n9908)
         );
  NAND2X1 U44901 ( .A(net151666), .B(net151653), .Y(n19852) );
  NOR4X1 U44902 ( .A(n29824), .B(n29825), .C(n29826), .D(n29827), .Y(net216243) );
  NOR4X1 U44903 ( .A(n29836), .B(n29837), .C(n29838), .D(n29839), .Y(net216246) );
  NOR4X1 U44904 ( .A(n26401), .B(n26402), .C(n26403), .D(n26404), .Y(net215146) );
  NOR4X1 U44905 ( .A(n26393), .B(n26394), .C(n26395), .D(n26396), .Y(net215148) );
  NOR4X1 U44906 ( .A(n26397), .B(n26398), .C(n26399), .D(n26400), .Y(net215149) );
  NOR4X1 U44907 ( .A(n30649), .B(n30650), .C(n30651), .D(n30652), .Y(net216397) );
  NOR4X1 U44908 ( .A(n26011), .B(n26012), .C(n26013), .D(n26014), .Y(net215049) );
  NOR4X1 U44909 ( .A(n29673), .B(n29674), .C(n29675), .D(n29676), .Y(net214758) );
  NOR4X1 U44910 ( .A(n29677), .B(n29678), .C(n29679), .D(n29680), .Y(net214759) );
  NAND4BX1 U44911 ( .AN(n47712), .B(n9771), .C(n47711), .D(n47710), .Y(n9739)
         );
  NOR3X1 U44912 ( .A(n47842), .B(n9877), .C(n47822), .Y(n47711) );
  NAND2X1 U44913 ( .A(n9772), .B(n9908), .Y(n47712) );
  NOR3X1 U44914 ( .A(n47709), .B(n9806), .C(n9876), .Y(n47710) );
  NOR4X1 U44915 ( .A(n26514), .B(n26515), .C(n26516), .D(n26517), .Y(net215182) );
  NOR4X1 U44916 ( .A(n26518), .B(n26519), .C(n26520), .D(n26521), .Y(net215183) );
  NAND4X1 U44917 ( .A(n43417), .B(n43416), .C(n43415), .D(n43414), .Y(n10427)
         );
  NOR4X1 U44918 ( .A(n30908), .B(n30909), .C(n30910), .D(n30911), .Y(n43417)
         );
  NOR4X1 U44919 ( .A(n30912), .B(n30913), .C(n30914), .D(n30915), .Y(n43416)
         );
  NOR4X1 U44920 ( .A(n30920), .B(n30921), .C(n30922), .D(n30923), .Y(n43414)
         );
  NOR4X1 U44921 ( .A(n30016), .B(n30017), .C(n30018), .D(n30019), .Y(net216264) );
  NOR3BX1 U44922 ( .AN(n10700), .B(n10702), .C(net171551), .Y(n9909) );
  NOR2X1 U44923 ( .A(n10249), .B(n47807), .Y(n41758) );
  NOR4X1 U44924 ( .A(n30136), .B(n30137), .C(n30138), .D(n30139), .Y(net216300) );
  NAND4X1 U44925 ( .A(n43456), .B(n43455), .C(n43454), .D(n43453), .Y(n10426)
         );
  NOR4X1 U44926 ( .A(n30517), .B(n30518), .C(n30519), .D(n30520), .Y(n43456)
         );
  NOR4X1 U44927 ( .A(n30521), .B(n30522), .C(n30523), .D(n30524), .Y(n43455)
         );
  NOR4X1 U44928 ( .A(n30529), .B(n30530), .C(n30531), .D(n30532), .Y(n43453)
         );
  NAND4X1 U44929 ( .A(n43544), .B(n43543), .C(n43542), .D(n43541), .Y(n10432)
         );
  NOR4X1 U44930 ( .A(n29613), .B(n29614), .C(n29615), .D(n29616), .Y(n43544)
         );
  NOR4X1 U44931 ( .A(n29617), .B(n29618), .C(n29619), .D(n29620), .Y(n43543)
         );
  NOR4X1 U44932 ( .A(n29625), .B(n29626), .C(n29627), .D(n29628), .Y(n43541)
         );
  NOR4X1 U44933 ( .A(n30377), .B(n30378), .C(n30379), .D(n30380), .Y(net216327) );
  NOR4X1 U44934 ( .A(n26247), .B(n26248), .C(n26249), .D(n26250), .Y(net215102) );
  NAND4X1 U44935 ( .A(n43539), .B(n43538), .C(n43537), .D(n43536), .Y(n10431)
         );
  NOR4X1 U44936 ( .A(n29493), .B(n29494), .C(n29495), .D(n29496), .Y(n43539)
         );
  NOR4X1 U44937 ( .A(n29497), .B(n29498), .C(n29499), .D(n29500), .Y(n43538)
         );
  NOR4X1 U44938 ( .A(n29505), .B(n29506), .C(n29507), .D(n29508), .Y(n43536)
         );
  NOR4X1 U44939 ( .A(n30046), .B(n30047), .C(n30048), .D(n30049), .Y(net216273) );
  NOR4X1 U44940 ( .A(n29643), .B(n29644), .C(n29645), .D(n29646), .Y(net214766) );
  NOR4X1 U44941 ( .A(n29647), .B(n29648), .C(n29649), .D(n29650), .Y(net214767) );
  NOR4X1 U44942 ( .A(n26454), .B(n26455), .C(n26456), .D(n26457), .Y(net214739) );
  NOR4X1 U44943 ( .A(n26458), .B(n26459), .C(n26460), .D(n26461), .Y(net214740) );
  NOR4X1 U44944 ( .A(n26217), .B(n26218), .C(n26219), .D(n26220), .Y(net214752) );
  NOR4X1 U44945 ( .A(n30437), .B(n30438), .C(n30439), .D(n30440), .Y(net216345) );
  NOR4X1 U44946 ( .A(n30347), .B(n30348), .C(n30349), .D(n30350), .Y(net214787) );
  NOR4X1 U44947 ( .A(n30166), .B(n30167), .C(n30168), .D(n30169), .Y(net216309) );
  NAND3BX1 U44948 ( .AN(n10018), .B(n21446), .C(n10016), .Y(n9885) );
  NOR4X1 U44949 ( .A(n30106), .B(n30107), .C(n30108), .D(n30109), .Y(net216291) );
  NOR4X1 U44950 ( .A(n30830), .B(n30831), .C(n30832), .D(n30833), .Y(net216489) );
  NOR4X1 U44951 ( .A(n30469), .B(n30470), .C(n30471), .D(n30472), .Y(net216426) );
  NOR4X1 U44952 ( .A(n26037), .B(n26038), .C(n26039), .D(n26040), .Y(net215057) );
  OAI21XL U44953 ( .A0(n10178), .A1(n9963), .B0(n50095), .Y(n10175) );
  CLKINVX1 U44954 ( .A(n9964), .Y(n50095) );
  AOI211X1 U44955 ( .A0(n47814), .A1(n47813), .B0(n47812), .C0(net210434), .Y(
        n10178) );
  NOR2X1 U44956 ( .A(net210444), .B(net210445), .Y(n47814) );
  NAND4X1 U44957 ( .A(n43436), .B(n43435), .C(n43434), .D(n43433), .Y(n10428)
         );
  NOR4X1 U44958 ( .A(n30577), .B(n30578), .C(n30579), .D(n30580), .Y(n43436)
         );
  NOR4X1 U44959 ( .A(n30581), .B(n30582), .C(n30583), .D(n30584), .Y(n43435)
         );
  NOR4X1 U44960 ( .A(n30589), .B(n30590), .C(n30591), .D(n30592), .Y(n43433)
         );
  NAND4X1 U44961 ( .A(n43520), .B(n43519), .C(n43518), .D(n43517), .Y(n10303)
         );
  NOR4X1 U44962 ( .A(n29794), .B(n29795), .C(n29796), .D(n29797), .Y(n43520)
         );
  NOR4X1 U44963 ( .A(n29798), .B(n29799), .C(n29800), .D(n29801), .Y(n43519)
         );
  NOR4X1 U44964 ( .A(n29806), .B(n29807), .C(n29808), .D(n29809), .Y(n43517)
         );
  NAND4X1 U44965 ( .A(n43476), .B(n43475), .C(n43474), .D(n43473), .Y(n10429)
         );
  NOR4X1 U44966 ( .A(n30305), .B(n30306), .C(n30307), .D(n30308), .Y(n43476)
         );
  NOR4X1 U44967 ( .A(n30309), .B(n30310), .C(n30311), .D(n30312), .Y(n43475)
         );
  NOR4X1 U44968 ( .A(n30317), .B(n30318), .C(n30319), .D(n30320), .Y(n43473)
         );
  NOR4X1 U44969 ( .A(n29734), .B(n29735), .C(n29736), .D(n29737), .Y(net216216) );
  NOR4X1 U44970 ( .A(n29738), .B(n29739), .C(n29740), .D(n29741), .Y(net216217) );
  NOR4X1 U44971 ( .A(n29553), .B(n29554), .C(n29555), .D(n29556), .Y(net216189) );
  NOR3X1 U44972 ( .A(n9870), .B(n9871), .C(n9872), .Y(n9759) );
  NOR4X1 U44973 ( .A(n25981), .B(n25982), .C(n25983), .D(n25984), .Y(net215040) );
  NOR4X1 U44974 ( .A(n29764), .B(n29765), .C(n29766), .D(n29767), .Y(net216225) );
  NOR4X1 U44975 ( .A(n29768), .B(n29769), .C(n29770), .D(n29771), .Y(net216226) );
  NOR4X1 U44976 ( .A(n26337), .B(n26338), .C(n26339), .D(n26340), .Y(net215129) );
  NOR4X1 U44977 ( .A(n26157), .B(n26158), .C(n26159), .D(n26160), .Y(net215093) );
  NOR4X1 U44978 ( .A(n29974), .B(n29975), .C(n29976), .D(n29977), .Y(net216254) );
  NOR4X1 U44979 ( .A(n29986), .B(n29987), .C(n29988), .D(n29989), .Y(net216253) );
  NOR4X1 U44980 ( .A(n26187), .B(n26188), .C(n26189), .D(n26190), .Y(net214748) );
  NOR4X1 U44981 ( .A(n29703), .B(n29704), .C(n29705), .D(n29706), .Y(net214762) );
  NOR4X1 U44982 ( .A(n29707), .B(n29708), .C(n29709), .D(n29710), .Y(net214763) );
  OAI31XL U44983 ( .A0(n10018), .A1(n10019), .A2(n10020), .B0(net151479), .Y(
        n10017) );
  NOR4X1 U44984 ( .A(n10022), .B(net171548), .C(n10024), .D(n10025), .Y(n10019) );
  NOR3X1 U44985 ( .A(n10026), .B(n10027), .C(n10028), .Y(n10022) );
  AOI211X1 U44986 ( .A0(n10029), .A1(n10030), .B0(n39657), .C0(n10032), .Y(
        n10027) );
  NOR4X1 U44987 ( .A(n30395), .B(n30396), .C(n30397), .D(n30398), .Y(net216333) );
  NOR4X1 U44988 ( .A(n30399), .B(n30400), .C(n30401), .D(n30402), .Y(net216334) );
  NOR4X1 U44989 ( .A(n30407), .B(n30408), .C(n30409), .D(n30410), .Y(net216336) );
  NOR2BX1 U44990 ( .AN(n10815), .B(n10814), .Y(n9863) );
  NOR4X1 U44991 ( .A(n10671), .B(net151431), .C(net171533), .D(net171534), .Y(
        n10012) );
  NAND3BX1 U44992 ( .AN(n10032), .B(n10033), .C(n10029), .Y(n9804) );
  NAND4X1 U44993 ( .A(n37346), .B(n10204), .C(n37123), .D(n10199), .Y(n9871)
         );
  NAND4X1 U44994 ( .A(n44376), .B(n44375), .C(n44374), .D(n44373), .Y(n12415)
         );
  NOR4X1 U44995 ( .A(n26093), .B(n26094), .C(n26095), .D(n26096), .Y(n44376)
         );
  NOR4X1 U44996 ( .A(n26097), .B(n26098), .C(n26099), .D(n26100), .Y(n44375)
         );
  NOR4X1 U44997 ( .A(n26101), .B(n26102), .C(n26103), .D(n26104), .Y(n44374)
         );
  NOR4X1 U44998 ( .A(n29854), .B(n29855), .C(n29856), .D(n29857), .Y(net216207) );
  NOR4X1 U44999 ( .A(n29866), .B(n29867), .C(n29868), .D(n29869), .Y(net216210) );
  NAND2BX1 U45000 ( .AN(n10679), .B(n10677), .Y(n9886) );
  NAND4X1 U45001 ( .A(n44329), .B(n44328), .C(n44327), .D(n44326), .Y(n12591)
         );
  NOR4X1 U45002 ( .A(n26484), .B(n26485), .C(n26486), .D(n26487), .Y(n44329)
         );
  NOR4X1 U45003 ( .A(n26488), .B(n26489), .C(n26490), .D(n26491), .Y(n44328)
         );
  NOR4X1 U45004 ( .A(n26492), .B(n26493), .C(n26494), .D(n26495), .Y(n44327)
         );
  NAND4X1 U45005 ( .A(n43467), .B(n43466), .C(n43465), .D(n43464), .Y(n12445)
         );
  NOR4X1 U45006 ( .A(n30607), .B(n30608), .C(n30609), .D(n30610), .Y(n43467)
         );
  NOR4X1 U45007 ( .A(n30611), .B(n30612), .C(n30613), .D(n30614), .Y(n43466)
         );
  NOR4X1 U45008 ( .A(n30619), .B(n30620), .C(n30621), .D(n30622), .Y(n43464)
         );
  NAND4X1 U45009 ( .A(n44371), .B(n44370), .C(n44369), .D(n44368), .Y(n12417)
         );
  NOR4X1 U45010 ( .A(n26123), .B(n26124), .C(n26125), .D(n26126), .Y(n44371)
         );
  NOR4X1 U45011 ( .A(n26127), .B(n26128), .C(n26129), .D(n26130), .Y(n44370)
         );
  NOR4X1 U45012 ( .A(n26131), .B(n26132), .C(n26133), .D(n26134), .Y(n44369)
         );
  NAND4X1 U45013 ( .A(n44349), .B(n44348), .C(n44347), .D(n44346), .Y(n12403)
         );
  NOR4X1 U45014 ( .A(n26363), .B(n26364), .C(n26365), .D(n26366), .Y(n44349)
         );
  NOR4X1 U45015 ( .A(n26367), .B(n26368), .C(n26369), .D(n26370), .Y(n44348)
         );
  NOR4X1 U45016 ( .A(n26371), .B(n26372), .C(n26373), .D(n26374), .Y(n44347)
         );
  NOR4X1 U45017 ( .A(n10865), .B(n10861), .C(net171486), .D(net171489), .Y(
        n10251) );
  NOR4X1 U45018 ( .A(n29884), .B(n29885), .C(n29886), .D(n29887), .Y(net214778) );
  NOR4X1 U45019 ( .A(n29896), .B(n29897), .C(n29898), .D(n29899), .Y(net214781) );
  AOI211X1 U45020 ( .A0(n10244), .A1(n10245), .B0(n10246), .C0(n10247), .Y(
        n10241) );
  OAI21XL U45021 ( .A0(n10248), .A1(n10249), .B0(n49492), .Y(n10245) );
  CLKINVX1 U45022 ( .A(n47807), .Y(n49492) );
  AOI211X1 U45023 ( .A0(n10251), .A1(n10252), .B0(n10253), .C0(n10254), .Y(
        n10248) );
  OAI31XL U45024 ( .A0(n10130), .A1(n10131), .A2(net151789), .B0(n50093), .Y(
        n10059) );
  CLKINVX1 U45025 ( .A(n9922), .Y(n50093) );
  AOI211X1 U45026 ( .A0(n10134), .A1(n10135), .B0(n10136), .C0(n10137), .Y(
        n10131) );
  OAI21XL U45027 ( .A0(n10138), .A1(n9950), .B0(n44625), .Y(n10135) );
  NAND4X1 U45028 ( .A(n43511), .B(n43510), .C(n43509), .D(n43508), .Y(n12590)
         );
  NOR4X1 U45029 ( .A(n30064), .B(n30065), .C(n30066), .D(n30067), .Y(n43511)
         );
  NOR4X1 U45030 ( .A(n30068), .B(n30069), .C(n30070), .D(n30071), .Y(n43510)
         );
  NOR4X1 U45031 ( .A(n30076), .B(n30077), .C(n30078), .D(n30079), .Y(n43508)
         );
  NAND4X1 U45032 ( .A(n43499), .B(n43498), .C(n43497), .D(n43496), .Y(n12433)
         );
  NOR4X1 U45033 ( .A(n30184), .B(n30185), .C(n30186), .D(n30187), .Y(n43499)
         );
  NOR4X1 U45034 ( .A(n30188), .B(n30189), .C(n30190), .D(n30191), .Y(n43498)
         );
  NOR4X1 U45035 ( .A(n30196), .B(n30197), .C(n30198), .D(n30199), .Y(n43496)
         );
  NAND4BX1 U45036 ( .AN(n9915), .B(n9909), .C(n19528), .D(n50099), .Y(n9806)
         );
  NOR2X1 U45037 ( .A(n9911), .B(n9913), .Y(n19528) );
  NAND3BX1 U45038 ( .AN(n10246), .B(n10244), .C(net168852), .Y(n9862) );
  NAND4X1 U45039 ( .A(n43491), .B(n43490), .C(n43489), .D(n43488), .Y(
        net209441) );
  NOR4X1 U45040 ( .A(n30215), .B(n30216), .C(n30217), .D(n30218), .Y(n43491)
         );
  NOR4X1 U45041 ( .A(n30219), .B(n30220), .C(n30221), .D(n30222), .Y(n43490)
         );
  NOR4X1 U45042 ( .A(n30227), .B(n30228), .C(n30229), .D(n30230), .Y(n43488)
         );
  NOR4X1 U45043 ( .A(n11521), .B(n10651), .C(net171524), .D(net171525), .Y(
        n10000) );
  NOR4X1 U45044 ( .A(n30679), .B(n30680), .C(n30681), .D(n30682), .Y(net216408) );
  NOR4X1 U45045 ( .A(n30245), .B(n30246), .C(n30247), .D(n30248), .Y(net216360) );
  NOR4X1 U45046 ( .A(n30249), .B(n30250), .C(n30251), .D(n30252), .Y(net216361) );
  NOR4X1 U45047 ( .A(n30257), .B(n30258), .C(n30259), .D(n30260), .Y(net216363) );
  NOR4X1 U45048 ( .A(n30499), .B(n30500), .C(n30501), .D(n30502), .Y(net216435) );
  NOR2X1 U45049 ( .A(n47822), .B(net218294), .Y(n9875) );
  NOR4X1 U45050 ( .A(n29914), .B(n29915), .C(n29916), .D(n29917), .Y(net214774) );
  NOR4X1 U45051 ( .A(n29926), .B(n29927), .C(n29928), .D(n29929), .Y(net214777) );
  NOR4X1 U45052 ( .A(n29583), .B(n29584), .C(n29585), .D(n29586), .Y(net216198) );
  NOR4X1 U45053 ( .A(n29587), .B(n29588), .C(n29589), .D(n29590), .Y(net216199) );
  NOR4X1 U45054 ( .A(n29595), .B(n29596), .C(n29597), .D(n29598), .Y(net216201) );
  NOR3X1 U45055 ( .A(n9919), .B(n9918), .C(n47841), .Y(n47844) );
  NOR2X1 U45056 ( .A(n37241), .B(n9747), .Y(n9743) );
  NAND2BX1 U45057 ( .AN(n9968), .B(n9969), .Y(n9797) );
  NOR3X1 U45058 ( .A(net171412), .B(n10210), .C(net151586), .Y(n10208) );
  NOR4X1 U45059 ( .A(n10212), .B(net171416), .C(n39537), .D(n10215), .Y(n10210) );
  AOI211X1 U45060 ( .A0(n10216), .A1(n10217), .B0(n10218), .C0(n10219), .Y(
        n10212) );
  OAI21XL U45061 ( .A0(n10220), .A1(n9854), .B0(n50107), .Y(n10217) );
  NOR4X1 U45062 ( .A(net171218), .B(n10164), .C(n40402), .D(n10166), .Y(n10161) );
  AOI211X1 U45063 ( .A0(n10167), .A1(n10168), .B0(n10169), .C0(n10170), .Y(
        n10164) );
  OAI21XL U45064 ( .A0(n10171), .A1(n10172), .B0(n10173), .Y(n10168) );
  AOI211X1 U45065 ( .A0(n10174), .A1(n10175), .B0(n40401), .C0(n10177), .Y(
        n10171) );
  CLKINVX1 U45066 ( .A(n47836), .Y(n47810) );
  NAND4X1 U45067 ( .A(n44581), .B(n44580), .C(n44579), .D(n44578), .Y(
        net214677) );
  NOR4X1 U45068 ( .A(n29944), .B(n29945), .C(n29946), .D(n29947), .Y(n44581)
         );
  NOR4X1 U45069 ( .A(n29948), .B(n29949), .C(n29950), .D(n29951), .Y(n44580)
         );
  NOR4X1 U45070 ( .A(n29956), .B(n29957), .C(n29958), .D(n29959), .Y(n44578)
         );
  NAND4X1 U45071 ( .A(n44381), .B(n44380), .C(n44379), .D(n44378), .Y(
        net214783) );
  NOR4X1 U45072 ( .A(n26063), .B(n26064), .C(n26065), .D(n26066), .Y(n44381)
         );
  NOR4X1 U45073 ( .A(n26067), .B(n26068), .C(n26069), .D(n26070), .Y(n44380)
         );
  NOR4X1 U45074 ( .A(n26071), .B(n26072), .C(n26073), .D(n26074), .Y(n44379)
         );
  NAND4X1 U45075 ( .A(n44356), .B(n44355), .C(n44354), .D(n44353), .Y(
        net214756) );
  NOR4X1 U45076 ( .A(n26273), .B(n26274), .C(n26275), .D(n26276), .Y(n44356)
         );
  NOR4X1 U45077 ( .A(n26277), .B(n26278), .C(n26279), .D(n26280), .Y(n44355)
         );
  NOR4X1 U45078 ( .A(n26281), .B(n26282), .C(n26283), .D(n26284), .Y(n44354)
         );
  NAND3BX1 U45079 ( .AN(n9978), .B(n41788), .C(n50096), .Y(n9865) );
  NAND3X1 U45080 ( .A(n10012), .B(n10010), .C(n21285), .Y(n9882) );
  NOR3BXL U45081 ( .AN(n36926), .B(net259841), .C(net151435), .Y(n21285) );
  NAND3BX1 U45082 ( .AN(n10219), .B(n10216), .C(net151557), .Y(n9968) );
  NOR2X1 U45083 ( .A(net210550), .B(net210552), .Y(n41759) );
  NOR2X1 U45084 ( .A(n47798), .B(n47800), .Y(n41760) );
  OAI21XL U45085 ( .A0(n10034), .A1(n9911), .B0(n9909), .Y(n10030) );
  AOI211X1 U45086 ( .A0(n50099), .A1(n10036), .B0(n9915), .C0(n9913), .Y(
        n10034) );
  OAI21XL U45087 ( .A0(n10037), .A1(n9918), .B0(n50097), .Y(n10036) );
  AOI21X1 U45088 ( .A0(n47828), .A1(n47827), .B0(n47826), .Y(n10037) );
  NOR4BBX1 U45089 ( .AN(n22472), .BN(n9859), .C(n9854), .D(n9855), .Y(n9757)
         );
  NOR3BXL U45090 ( .AN(n9863), .B(n9858), .C(n9857), .Y(n22472) );
  NAND2X1 U45091 ( .A(n41759), .B(n46605), .Y(n47834) );
  CLKINVX1 U45092 ( .A(n47799), .Y(n46605) );
  NOR2X1 U45093 ( .A(n47801), .B(n47800), .Y(n47804) );
  AOI21X1 U45094 ( .A0(n41759), .A1(n47799), .B0(n47798), .Y(n47801) );
  NOR2X1 U45095 ( .A(n22098), .B(n9862), .Y(n46606) );
  NAND3BX1 U45096 ( .AN(n9870), .B(n9798), .C(n9757), .Y(n22098) );
  CLKINVX1 U45097 ( .A(n9914), .Y(n50099) );
  NAND2X1 U45098 ( .A(n40269), .B(n37544), .Y(n48701) );
  NAND2X1 U45099 ( .A(n40274), .B(n37545), .Y(n48857) );
  NAND2X1 U45100 ( .A(n40274), .B(n37546), .Y(n48860) );
  NAND2X1 U45101 ( .A(n40275), .B(n37547), .Y(n49013) );
  NAND2X1 U45102 ( .A(n40194), .B(n37548), .Y(n49016) );
  NAND2X1 U45103 ( .A(net217936), .B(n37541), .Y(n49167) );
  NAND2X1 U45104 ( .A(n40242), .B(n37542), .Y(n49322) );
  NAND2X1 U45105 ( .A(net217942), .B(n37543), .Y(n49325) );
  NAND2X1 U45106 ( .A(n40269), .B(n37549), .Y(n48722) );
  NAND2X1 U45107 ( .A(n40267), .B(n37550), .Y(n48880) );
  NAND2X1 U45108 ( .A(n40256), .B(n37551), .Y(n49032) );
  NAND2X1 U45109 ( .A(net217936), .B(n37552), .Y(n49188) );
  NAND2X1 U45110 ( .A(n40247), .B(n37553), .Y(n49343) );
  CLKINVX1 U45111 ( .A(n9979), .Y(n50096) );
  OR4X1 U45112 ( .A(n9994), .B(n9999), .C(net171528), .D(net171530), .Y(n9901)
         );
  CLKINVX1 U45113 ( .A(n10779), .Y(net151587) );
  CLKINVX1 U45114 ( .A(n9919), .Y(n50097) );
  NOR2X2 U45115 ( .A(n50144), .B(net171380), .Y(n19249) );
  NOR4X1 U45116 ( .A(n25707), .B(n25708), .C(n25709), .D(n25710), .Y(net214958) );
  NOR4X1 U45117 ( .A(n26574), .B(n26575), .C(n26576), .D(n26577), .Y(net215200) );
  NOR4X1 U45118 ( .A(n26578), .B(n26579), .C(n26580), .D(n26581), .Y(net215201) );
  NOR4X1 U45119 ( .A(n26582), .B(n26583), .C(n26584), .D(n26585), .Y(net215202) );
  NOR4X1 U45120 ( .A(n26428), .B(n26429), .C(n26430), .D(n26431), .Y(net214744) );
  NOR4X1 U45121 ( .A(n26604), .B(n26605), .C(n26606), .D(n26607), .Y(net215155) );
  NOR4X1 U45122 ( .A(n26608), .B(n26609), .C(n26610), .D(n26611), .Y(net215156) );
  NOR3BX1 U45123 ( .AN(n10167), .B(n10169), .C(n10170), .Y(n9958) );
  NOR4X1 U45124 ( .A(n26548), .B(n26549), .C(n26550), .D(n26551), .Y(net215192) );
  NOR4X1 U45125 ( .A(n25831), .B(n25832), .C(n25833), .D(n25834), .Y(net215013) );
  AO21X1 U45126 ( .A0(n9958), .A1(n9959), .B0(n9787), .Y(n9956) );
  OAI21XL U45127 ( .A0(n9960), .A1(n9788), .B0(n9847), .Y(n9959) );
  AOI211X1 U45128 ( .A0(n9961), .A1(n9962), .B0(n9963), .C0(n9964), .Y(n9960)
         );
  NAND2X1 U45129 ( .A(n47838), .B(n47837), .Y(n9962) );
  NAND4X1 U45130 ( .A(n44409), .B(n44408), .C(n44407), .D(n44406), .Y(n10435)
         );
  NOR4X1 U45131 ( .A(n25883), .B(n25884), .C(n25885), .D(n25886), .Y(n44409)
         );
  NOR4X1 U45132 ( .A(n25887), .B(n25888), .C(n25889), .D(n25890), .Y(n44408)
         );
  NOR4X1 U45133 ( .A(n25891), .B(n25892), .C(n25893), .D(n25894), .Y(n44407)
         );
  NOR4X1 U45134 ( .A(n26634), .B(n26635), .C(n26636), .D(n26637), .Y(net215164) );
  NOR4X1 U45135 ( .A(n26638), .B(n26639), .C(n26640), .D(n26641), .Y(net215165) );
  NOR4X1 U45136 ( .A(n26642), .B(n26643), .C(n26644), .D(n26645), .Y(net215166) );
  NOR4X1 U45137 ( .A(n10456), .B(n11904), .C(net171283), .D(net171288), .Y(
        n10134) );
  NOR2BX1 U45138 ( .AN(n10173), .B(n10172), .Y(n9847) );
  NOR4X1 U45139 ( .A(net171272), .B(net171274), .C(net151786), .D(net151788),
        .Y(n9946) );
  NOR4X1 U45140 ( .A(n25793), .B(n25794), .C(n25795), .D(n25796), .Y(net214984) );
  NOR4X1 U45141 ( .A(n25797), .B(n25798), .C(n25799), .D(n25800), .Y(net214985) );
  NOR4X1 U45142 ( .A(n24690), .B(n24691), .C(n24692), .D(n24693), .Y(net214735) );
  NOR4X1 U45143 ( .A(n24694), .B(n24695), .C(n24696), .D(n24697), .Y(net214736) );
  NOR4X1 U45144 ( .A(n24698), .B(n24699), .C(n24700), .D(n24701), .Y(net214737) );
  AOI211X1 U45145 ( .A0(n50101), .A1(n9906), .B0(n9886), .C0(n9884), .Y(n9902)
         );
  CLKINVX1 U45146 ( .A(n9885), .Y(n50101) );
  OAI21XL U45147 ( .A0(n9907), .A1(n9804), .B0(n9908), .Y(n9906) );
  NOR3BXL U45148 ( .AN(n9909), .B(n9910), .C(n9911), .Y(n9907) );
  NOR3BXL U45149 ( .AN(n10140), .B(n10143), .C(n10142), .Y(n9948) );
  NOR4X1 U45150 ( .A(n9922), .B(n10130), .C(net151789), .D(n9945), .Y(n9851)
         );
  NOR3X1 U45151 ( .A(n50111), .B(n9954), .C(n9837), .Y(n30441) );
  OAI31XL U45152 ( .A0(n9836), .A1(n9837), .A2(n9838), .B0(n49499), .Y(n9810)
         );
  OAI31XL U45153 ( .A0(n9839), .A1(n9840), .A2(n9841), .B0(n50109), .Y(n9836)
         );
  OAI31XL U45154 ( .A0(n9787), .A1(n9843), .A2(n49520), .B0(n9844), .Y(n9839)
         );
  AOI211X1 U45155 ( .A0(n9845), .A1(n9846), .B0(n9788), .C0(n45522), .Y(n9843)
         );
  OAI31XL U45156 ( .A0(n9853), .A1(n9854), .A2(n9855), .B0(n50105), .Y(n9809)
         );
  OAI31XL U45157 ( .A0(n9856), .A1(n9857), .A2(n9858), .B0(n9859), .Y(n9853)
         );
  OAI31XL U45158 ( .A0(n50090), .A1(n50091), .A2(n9862), .B0(n9863), .Y(n9856)
         );
  CLKINVX1 U45159 ( .A(n9864), .Y(n50091) );
  OAI211X1 U45160 ( .A0(n9944), .A1(n9945), .B0(n40387), .C0(net151779), .Y(
        n9921) );
  AOI211X1 U45161 ( .A0(n9948), .A1(n9949), .B0(n9950), .C0(n9951), .Y(n9944)
         );
  OAI211X1 U45162 ( .A0(n9952), .A1(n9838), .B0(n50109), .C0(n50106), .Y(n9949) );
  AOI211X1 U45163 ( .A0(n49521), .A1(n9956), .B0(n9840), .C0(n50111), .Y(n9952) );
  AOI211X1 U45164 ( .A0(n9898), .A1(n9899), .B0(n9900), .C0(n9901), .Y(n9896)
         );
  OAI211X1 U45165 ( .A0(n9902), .A1(n9882), .B0(n50110), .C0(n50108), .Y(n9899) );
  CLKINVX1 U45166 ( .A(n9880), .Y(n50110) );
  NOR4X1 U45167 ( .A(n10542), .B(n10609), .C(net171304), .D(net171307), .Y(
        n10167) );
  NOR2X1 U45168 ( .A(n50144), .B(n9747), .Y(n9707) );
  NOR4X1 U45169 ( .A(n9912), .B(n9913), .C(n9914), .D(n9915), .Y(n9910) );
  AOI211X1 U45170 ( .A0(n49491), .A1(n9917), .B0(n9918), .C0(n9919), .Y(n9912)
         );
  NAND2X1 U45171 ( .A(n47845), .B(n47843), .Y(n9917) );
  CLKINVX1 U45172 ( .A(n47841), .Y(n49491) );
  NOR2X1 U45173 ( .A(n9716), .B(n50144), .Y(n9748) );
  NAND4X1 U45174 ( .A(n44393), .B(n44392), .C(n44391), .D(n44390), .Y(
        net214782) );
  NOR4X1 U45175 ( .A(n25943), .B(n25944), .C(n25945), .D(n25946), .Y(n44393)
         );
  NOR4X1 U45176 ( .A(n25947), .B(n25948), .C(n25949), .D(n25950), .Y(n44392)
         );
  NOR4X1 U45177 ( .A(n25951), .B(n25952), .C(n25953), .D(n25954), .Y(n44391)
         );
  NAND4X1 U45178 ( .A(net235251), .B(net210670), .C(net210650), .D(n45527),
        .Y(n47816) );
  NAND4X1 U45179 ( .A(n44420), .B(n44419), .C(n44418), .D(n44417), .Y(
        net214757) );
  NOR4X1 U45180 ( .A(n25733), .B(n25734), .C(n25735), .D(n25736), .Y(n44420)
         );
  NOR4X1 U45181 ( .A(n25737), .B(n25738), .C(n25739), .D(n25740), .Y(n44419)
         );
  NOR4X1 U45182 ( .A(n25741), .B(n25742), .C(n25743), .D(n25744), .Y(n44418)
         );
  NAND4X1 U45183 ( .A(n44415), .B(n44414), .C(n44413), .D(n44412), .Y(
        net214755) );
  NOR4X1 U45184 ( .A(n25763), .B(n25764), .C(n25765), .D(n25766), .Y(n44415)
         );
  NOR4X1 U45185 ( .A(n25767), .B(n25768), .C(n25769), .D(n25770), .Y(n44414)
         );
  NOR4X1 U45186 ( .A(n25771), .B(n25772), .C(n25773), .D(n25774), .Y(n44413)
         );
  NAND4BX1 U45187 ( .AN(n10155), .B(n10158), .C(n10162), .D(n31164), .Y(n9841)
         );
  NOR4X1 U45188 ( .A(net171132), .B(net171134), .C(net171136), .D(net171139),
        .Y(n31164) );
  NOR2X1 U45189 ( .A(n10512), .B(n10509), .Y(n9844) );
  NOR4X1 U45190 ( .A(n9879), .B(n9880), .C(n9881), .D(n9882), .Y(n9878) );
  NOR4X1 U45191 ( .A(n9883), .B(n9884), .C(n9885), .D(n9886), .Y(n9879) );
  AOI211X1 U45192 ( .A0(n50094), .A1(n9888), .B0(n9804), .C0(n49517), .Y(n9883) );
  OAI2BB1X1 U45193 ( .A0N(n47846), .A1N(n47845), .B0(n47844), .Y(n9888) );
  NAND4X1 U45194 ( .A(net210443), .B(net213950), .C(net234007), .D(n37509),
        .Y(n47838) );
  CLKINVX1 U45195 ( .A(net210441), .Y(net213950) );
  OAI21XL U45196 ( .A0(n9974), .A1(n50098), .B0(n41758), .Y(n9973) );
  CLKINVX1 U45197 ( .A(n9799), .Y(n50098) );
  AOI211X1 U45198 ( .A0(n41788), .A1(n9977), .B0(n9978), .C0(n9979), .Y(n9974)
         );
  NAND2X1 U45199 ( .A(n41760), .B(n47834), .Y(n9977) );
  NAND3X1 U45200 ( .A(n9948), .B(n44625), .C(n44624), .Y(n50104) );
  CLKINVX1 U45201 ( .A(n9950), .Y(n44624) );
  CLKINVX1 U45202 ( .A(n9951), .Y(n44625) );
  OAI21XL U45203 ( .A0(n50141), .A1(n9716), .B0(n50137), .Y(n9732) );
  NAND3X1 U45204 ( .A(n47810), .B(n45521), .C(n45520), .Y(n9846) );
  CLKINVX1 U45205 ( .A(n47838), .Y(n45521) );
  CLKINVX1 U45206 ( .A(n47835), .Y(n45520) );
  OAI21XL U45207 ( .A0(n9967), .A1(n9968), .B0(n9969), .Y(n9966) );
  AOI211X1 U45208 ( .A0(n9859), .A1(n9970), .B0(n9855), .C0(n9854), .Y(n9967)
         );
  OAI211X1 U45209 ( .A0(n9971), .A1(n9858), .B0(n9863), .C0(n50112), .Y(n9970)
         );
  AOI21X1 U45210 ( .A0(n50084), .A1(n9973), .B0(n50090), .Y(n9971) );
  NOR2X1 U45211 ( .A(n47836), .B(n47835), .Y(n47837) );
  CLKINVX1 U45212 ( .A(n9881), .Y(n50108) );
  CLKINVX1 U45213 ( .A(n9857), .Y(n50112) );
  CLKINVX1 U45214 ( .A(n9855), .Y(n50107) );
  CLKINVX1 U45215 ( .A(n10196), .Y(n50100) );
  OAI21X1 U45216 ( .A0(n9702), .A1(n9737), .B0(n19449), .Y(n19487) );
  CLKINVX1 U45217 ( .A(n9704), .Y(n50146) );
  NOR2X1 U45218 ( .A(n50137), .B(n9702), .Y(n19523) );
  CLKINVX1 U45219 ( .A(n9877), .Y(n49518) );
  CLKINVX1 U45220 ( .A(n9837), .Y(n50106) );
  CLKINVX1 U45221 ( .A(n9954), .Y(n50109) );
  AOI21X2 U45222 ( .A0(n19283), .A1(n19336), .B0(n19180), .Y(n19290) );
  NOR2X2 U45223 ( .A(n19238), .B(n19239), .Y(n19207) );
  AOI2BB1X2 U45224 ( .A0N(n50138), .A1N(n19238), .B0(n19180), .Y(n19208) );
  OA21X2 U45225 ( .A0(n9679), .A1(n19374), .B0(n50142), .Y(n19381) );
  NAND2BX2 U45226 ( .AN(n19374), .B(n50139), .Y(n19344) );
  OA21X2 U45227 ( .A0(n50139), .A1(n19374), .B0(n50142), .Y(n19343) );
  NOR2X1 U45228 ( .A(n50137), .B(n50146), .Y(n19281) );
  NAND2X1 U45229 ( .A(n19283), .B(n19278), .Y(n19238) );
  AND4XL U45230 ( .A(n50142), .B(n19278), .C(n19335), .D(n50144), .Y(n32368)
         );
  NOR2X1 U45231 ( .A(n50129), .B(n9702), .Y(n19522) );
  CLKINVX1 U45232 ( .A(n9742), .Y(n50129) );
  CLKINVX1 U45233 ( .A(n9737), .Y(n50132) );
  CLKBUFX3 U45234 ( .A(n19382), .Y(n42729) );
  CLKINVX1 U45235 ( .A(n19334), .Y(n50139) );
  CLKBUFX3 U45236 ( .A(n19292), .Y(n42731) );
  CLKINVX1 U45237 ( .A(n19239), .Y(n50138) );
  CLKINVX1 U45238 ( .A(n9730), .Y(n50133) );
  CLKBUFX3 U45239 ( .A(n19420), .Y(n42728) );
  CLKINVX1 U45240 ( .A(n37525), .Y(n42733) );
  CLKBUFX3 U45241 ( .A(n19382), .Y(n42730) );
  CLKBUFX3 U45242 ( .A(n42321), .Y(n42449) );
  CLKBUFX3 U45243 ( .A(n42321), .Y(n42448) );
  CLKBUFX3 U45244 ( .A(n42321), .Y(n42447) );
  CLKBUFX3 U45245 ( .A(n42320), .Y(n42446) );
  CLKBUFX3 U45246 ( .A(n42320), .Y(n42445) );
  CLKBUFX3 U45247 ( .A(n42320), .Y(n42444) );
  CLKBUFX3 U45248 ( .A(n42319), .Y(n42443) );
  CLKBUFX3 U45249 ( .A(n42319), .Y(n42442) );
  CLKBUFX3 U45250 ( .A(n42319), .Y(n42441) );
  CLKBUFX3 U45251 ( .A(n42318), .Y(n42440) );
  CLKBUFX3 U45252 ( .A(n42318), .Y(n42439) );
  CLKBUFX3 U45253 ( .A(n42317), .Y(n42438) );
  CLKBUFX3 U45254 ( .A(n42317), .Y(n42437) );
  CLKBUFX3 U45255 ( .A(n42317), .Y(n42436) );
  NOR2X1 U45256 ( .A(n44031), .B(n44030), .Y(n44037) );
  NOR4X1 U45257 ( .A(n43866), .B(n43865), .C(n43864), .D(n43863), .Y(n43872)
         );
  NOR4X1 U45258 ( .A(n43862), .B(n43861), .C(n43860), .D(n43859), .Y(n43873)
         );
  NAND4X1 U45259 ( .A(n46246), .B(n46245), .C(n46244), .D(n46243), .Y(n46247)
         );
  NAND4X1 U45260 ( .A(n46242), .B(n46241), .C(n46240), .D(n46239), .Y(n46248)
         );
  NOR4X1 U45261 ( .A(n44021), .B(n44020), .C(n44019), .D(n44018), .Y(n44027)
         );
  NOR4X1 U45262 ( .A(n44043), .B(n44042), .C(n44041), .D(n44040), .Y(n44059)
         );
  NOR4X1 U45263 ( .A(n44047), .B(n44046), .C(n44045), .D(n44044), .Y(n44058)
         );
  NOR4X1 U45264 ( .A(n43920), .B(n43919), .C(n43918), .D(n43917), .Y(n43936)
         );
  NOR4X1 U45265 ( .A(n44856), .B(n44855), .C(n44854), .D(n44853), .Y(n44872)
         );
  NOR4X1 U45266 ( .A(n43951), .B(n43950), .C(n43949), .D(n43948), .Y(n43967)
         );
  NOR4X1 U45267 ( .A(n43959), .B(n43958), .C(n43957), .D(n43956), .Y(n43965)
         );
  NOR4X1 U45268 ( .A(n43955), .B(n43954), .C(n43953), .D(n43952), .Y(n43966)
         );
  CLKINVX1 U45269 ( .A(n12384), .Y(net171483) );
  NOR4X1 U45270 ( .A(n44715), .B(n44714), .C(n44713), .D(n44712), .Y(n44719)
         );
  NOR4X1 U45271 ( .A(n44711), .B(n44710), .C(n44709), .D(n44708), .Y(n44720)
         );
  NOR4X1 U45272 ( .A(n43990), .B(n43989), .C(n43988), .D(n43987), .Y(n43996)
         );
  NOR4X1 U45273 ( .A(n45473), .B(n45472), .C(n45471), .D(n45470), .Y(n45484)
         );
  XOR2X1 U45274 ( .A(n41806), .B(n36893), .Y(n45072) );
  NOR4X1 U45275 ( .A(n43889), .B(n43888), .C(n43887), .D(n43886), .Y(n43905)
         );
  CLKINVX1 U45276 ( .A(net210620), .Y(net210585) );
  CLKINVX1 U45277 ( .A(n12385), .Y(net171490) );
  NOR2X1 U45278 ( .A(net151751), .B(net151612), .Y(n11108) );
  CLKINVX1 U45279 ( .A(n10572), .Y(net151733) );
  NOR2X1 U45280 ( .A(net151848), .B(net151738), .Y(n11096) );
  CLKINVX1 U45281 ( .A(n12731), .Y(n49508) );
  NAND2X1 U45282 ( .A(n11084), .B(n11085), .Y(n11081) );
  AND2X2 U45283 ( .A(n11208), .B(n11209), .Y(n11086) );
  NAND2X1 U45284 ( .A(n11398), .B(n11399), .Y(n11395) );
  NAND2X1 U45285 ( .A(n11051), .B(n11052), .Y(n11048) );
  CLKINVX1 U45286 ( .A(n12797), .Y(net171199) );
  NAND2X1 U45287 ( .A(n12016), .B(n12017), .Y(n12013) );
  CLKINVX1 U45288 ( .A(n12692), .Y(net171200) );
  NAND2X1 U45289 ( .A(n11350), .B(n11351), .Y(n11347) );
  NOR2X1 U45290 ( .A(net171124), .B(net171122), .Y(n11998) );
  CLKINVX1 U45291 ( .A(n10518), .Y(net151456) );
  NOR2X1 U45292 ( .A(net171477), .B(net171478), .Y(n10993) );
  NAND2X1 U45293 ( .A(n10257), .B(n11149), .Y(n11146) );
  CLKINVX1 U45294 ( .A(net210584), .Y(net210557) );
  NOR4X1 U45295 ( .A(n44074), .B(n44073), .C(n44072), .D(n44071), .Y(n44090)
         );
  NOR4X1 U45296 ( .A(n44078), .B(n44077), .C(n44076), .D(n44075), .Y(n44089)
         );
  CLKINVX1 U45297 ( .A(n10570), .Y(net151723) );
  NAND3X1 U45298 ( .A(n46581), .B(n46580), .C(n46579), .Y(n46585) );
  NAND3X1 U45299 ( .A(n46578), .B(n46577), .C(n46576), .Y(n46586) );
  NOR4X1 U45300 ( .A(n44806), .B(n44805), .C(n44804), .D(n44803), .Y(n44812)
         );
  NOR2X1 U45301 ( .A(net151758), .B(net151757), .Y(n12056) );
  NOR2X1 U45302 ( .A(net151435), .B(net151431), .Y(n11308) );
  NOR4X1 U45303 ( .A(n44680), .B(n44679), .C(n44678), .D(n44677), .Y(n44691)
         );
  NAND2X1 U45304 ( .A(n10734), .B(n10733), .Y(n11436) );
  CLKINVX1 U45305 ( .A(n10751), .Y(net151847) );
  NOR2X1 U45306 ( .A(net151737), .B(net171540), .Y(n11390) );
  NOR2X1 U45307 ( .A(net171142), .B(n39335), .Y(n11980) );
  NOR2X1 U45308 ( .A(net151451), .B(net151453), .Y(n11328) );
  CLKINVX1 U45309 ( .A(n11065), .Y(net151644) );
  XNOR2X1 U45310 ( .A(n36857), .B(n42058), .Y(n46291) );
  NOR2X1 U45311 ( .A(n46284), .B(n46283), .Y(n46290) );
  NOR4X1 U45312 ( .A(n46288), .B(n46287), .C(n46286), .D(n46285), .Y(n46289)
         );
  NOR4X1 U45313 ( .A(n44736), .B(n44735), .C(n44734), .D(n44733), .Y(n44752)
         );
  NOR4X1 U45314 ( .A(n44740), .B(n44739), .C(n44738), .D(n44737), .Y(n44751)
         );
  NOR4X1 U45315 ( .A(n44744), .B(n44743), .C(n44742), .D(n44741), .Y(n44750)
         );
  XNOR2X1 U45316 ( .A(n51009), .B(n41291), .Y(n23804) );
  XNOR2X1 U45317 ( .A(n51008), .B(n41291), .Y(n23814) );
  XNOR2X1 U45318 ( .A(n51436), .B(n42698), .Y(n28033) );
  XNOR2X1 U45319 ( .A(n51434), .B(n42698), .Y(n28063) );
  XNOR2X1 U45320 ( .A(n51223), .B(n41333), .Y(n23805) );
  XNOR2X1 U45321 ( .A(n51222), .B(n41332), .Y(n23815) );
  XNOR2X1 U45322 ( .A(n50790), .B(net219466), .Y(n27458) );
  XNOR2X1 U45323 ( .A(n51430), .B(n42642), .Y(n27454) );
  XNOR2X1 U45324 ( .A(n50789), .B(n42592), .Y(n27450) );
  XNOR2X1 U45325 ( .A(n50785), .B(net219466), .Y(n27548) );
  XNOR2X1 U45326 ( .A(n51425), .B(n42642), .Y(n27544) );
  XNOR2X1 U45327 ( .A(n50784), .B(n42592), .Y(n27540) );
  XNOR2X1 U45328 ( .A(n51435), .B(n42643), .Y(n28025) );
  XNOR2X1 U45329 ( .A(n50794), .B(n42590), .Y(n28021) );
  XNOR2X1 U45330 ( .A(n51433), .B(n42643), .Y(n28055) );
  XNOR2X1 U45331 ( .A(n50795), .B(n36853), .Y(n23806) );
  XNOR2X1 U45332 ( .A(n50794), .B(n36853), .Y(n23816) );
  XNOR2X1 U45333 ( .A(n51004), .B(net219308), .Y(n27456) );
  XNOR2X1 U45334 ( .A(n50371), .B(n42675), .Y(n27452) );
  XNOR2X1 U45335 ( .A(n51003), .B(n42618), .Y(n27448) );
  XNOR2X1 U45336 ( .A(n50998), .B(n42618), .Y(n27538) );
  XNOR2X1 U45337 ( .A(n50376), .B(n36907), .Y(n28023) );
  XNOR2X1 U45338 ( .A(n51008), .B(n42619), .Y(n28019) );
  XNOR2X1 U45339 ( .A(n50375), .B(n42712), .Y(n28061) );
  XNOR2X1 U45340 ( .A(n50374), .B(n42671), .Y(n28053) );
  XNOR2X1 U45341 ( .A(n51006), .B(n42619), .Y(n28049) );
  XNOR2X1 U45342 ( .A(n50795), .B(n42508), .Y(n27681) );
  XNOR2X1 U45343 ( .A(n51218), .B(n41283), .Y(n27457) );
  XNOR2X1 U45344 ( .A(n50575), .B(n36903), .Y(n27453) );
  XNOR2X1 U45345 ( .A(n51217), .B(n42629), .Y(n27449) );
  XNOR2X1 U45346 ( .A(n50570), .B(n36903), .Y(n27543) );
  XNOR2X1 U45347 ( .A(n51212), .B(n42632), .Y(n27539) );
  XNOR2X1 U45348 ( .A(n50580), .B(n41380), .Y(n28024) );
  XNOR2X1 U45349 ( .A(n51222), .B(n42630), .Y(n28020) );
  XNOR2X1 U45350 ( .A(n50579), .B(n42725), .Y(n28062) );
  XOR2X1 U45351 ( .A(n41846), .B(n36891), .Y(n28060) );
  XOR2X1 U45352 ( .A(n42105), .B(n36885), .Y(n28064) );
  XOR2X1 U45353 ( .A(n41854), .B(n36894), .Y(n27549) );
  XOR2X1 U45354 ( .A(n41844), .B(n36894), .Y(n28030) );
  XOR2X1 U45355 ( .A(n42103), .B(n36880), .Y(n28034) );
  XOR2X1 U45356 ( .A(n42106), .B(n42655), .Y(n28056) );
  XOR2X1 U45357 ( .A(n41847), .B(n36819), .Y(n28052) );
  XOR2X1 U45358 ( .A(n41842), .B(n36894), .Y(n27700) );
  XOR2X1 U45359 ( .A(n41850), .B(n36895), .Y(n27489) );
  XOR2X1 U45360 ( .A(n42114), .B(n42663), .Y(n27545) );
  XOR2X1 U45361 ( .A(n42101), .B(n36883), .Y(n27704) );
  XOR2X1 U45362 ( .A(n42109), .B(n36887), .Y(n27493) );
  XOR2X1 U45363 ( .A(n42111), .B(n36887), .Y(n27613) );
  XOR2X1 U45364 ( .A(n41808), .B(n42519), .Y(n45055) );
  XOR2X1 U45365 ( .A(n36760), .B(n41807), .Y(n47674) );
  XOR2X1 U45366 ( .A(n41318), .B(n41808), .Y(n46587) );
  XOR2X1 U45367 ( .A(n36756), .B(n41808), .Y(n47697) );
  XOR2X1 U45368 ( .A(n36801), .B(n42098), .Y(n44002) );
  XOR2X1 U45369 ( .A(n42495), .B(n42080), .Y(n47339) );
  XOR2X1 U45370 ( .A(n42495), .B(n42084), .Y(n47427) );
  XOR2X1 U45371 ( .A(n36740), .B(n41798), .Y(n47668) );
  XOR2X1 U45372 ( .A(net219468), .B(n42058), .Y(n43863) );
  XOR2X1 U45373 ( .A(n41828), .B(n36901), .Y(n44651) );
  XOR2X1 U45374 ( .A(n41809), .B(n42597), .Y(n44881) );
  XOR2X1 U45375 ( .A(n41809), .B(n36891), .Y(n44919) );
  XOR2X1 U45376 ( .A(n41818), .B(n36898), .Y(n45501) );
  XOR2X1 U45377 ( .A(n41819), .B(n42611), .Y(n45493) );
  XOR2X1 U45378 ( .A(n41807), .B(n36900), .Y(n45091) );
  XOR2X1 U45379 ( .A(n41840), .B(n42612), .Y(n43887) );
  XOR2X1 U45380 ( .A(n42067), .B(n42659), .Y(n44885) );
  XOR2X1 U45381 ( .A(n42062), .B(n36907), .Y(n45012) );
  XOR2X1 U45382 ( .A(n42065), .B(n36801), .Y(n45000) );
  XOR2X1 U45383 ( .A(n41844), .B(n41312), .Y(n23807) );
  XOR2X1 U45384 ( .A(n42493), .B(n42065), .Y(n47679) );
  XOR2X1 U45385 ( .A(n36816), .B(n42066), .Y(n46592) );
  XOR2X1 U45386 ( .A(n42494), .B(n42066), .Y(n47702) );
  XOR2X1 U45387 ( .A(n42470), .B(n42057), .Y(n47665) );
  XOR2X1 U45388 ( .A(n42584), .B(n42060), .Y(n44003) );
  XOR2X1 U45389 ( .A(n41848), .B(n42516), .Y(n28042) );
  XOR2X1 U45390 ( .A(n42060), .B(n41319), .Y(n44017) );
  XOR2X1 U45391 ( .A(n41801), .B(n42633), .Y(n44013) );
  XOR2X1 U45392 ( .A(n41804), .B(n42614), .Y(n44012) );
  XOR2X1 U45393 ( .A(n41799), .B(n36825), .Y(n44034) );
  XOR2X1 U45394 ( .A(n36764), .B(n42059), .Y(n47671) );
  XOR2X1 U45395 ( .A(n41281), .B(n41802), .Y(n43866) );
  XOR2X1 U45396 ( .A(n36839), .B(n42063), .Y(n46288) );
  XOR2X1 U45397 ( .A(n36870), .B(n41805), .Y(n43865) );
  XOR2X1 U45398 ( .A(n36735), .B(n42062), .Y(n47670) );
  XOR2X1 U45399 ( .A(n36714), .B(n41800), .Y(n47666) );
  XOR2X1 U45400 ( .A(n36777), .B(n42060), .Y(n46276) );
  NOR2X1 U45401 ( .A(n47545), .B(n47544), .Y(n47549) );
  NOR4X1 U45402 ( .A(n20381), .B(n20382), .C(n47547), .D(n47546), .Y(n47548)
         );
  XOR2X1 U45403 ( .A(n41800), .B(n41282), .Y(n45074) );
  XOR2X1 U45404 ( .A(n42057), .B(net219434), .Y(n45071) );
  NOR4X1 U45405 ( .A(n27468), .B(n27469), .C(n27470), .D(n27473), .Y(n45688)
         );
  NOR3X1 U45406 ( .A(n45687), .B(n45686), .C(n45685), .Y(n45689) );
  XOR2X1 U45407 ( .A(n42107), .B(n36877), .Y(n28043) );
  XOR2X1 U45408 ( .A(n42057), .B(n36731), .Y(n45045) );
  XOR2X1 U45409 ( .A(n41800), .B(n36832), .Y(n45048) );
  XOR2X1 U45410 ( .A(n42544), .B(n41804), .Y(n44000) );
  XOR2X1 U45411 ( .A(n41292), .B(n41804), .Y(n46272) );
  XOR2X1 U45412 ( .A(n42554), .B(n41801), .Y(n44001) );
  XNOR2X1 U45413 ( .A(n36850), .B(n42057), .Y(n46565) );
  XNOR2X1 U45414 ( .A(n36808), .B(n42064), .Y(n46569) );
  NOR4X1 U45415 ( .A(n27730), .B(n27727), .C(n27734), .D(n27732), .Y(n43847)
         );
  NOR4X1 U45416 ( .A(n27701), .B(n27702), .C(n27703), .D(n27704), .Y(n43834)
         );
  XNOR2X1 U45417 ( .A(n50379), .B(n42711), .Y(n27701) );
  XNOR2X1 U45418 ( .A(n49511), .B(n42724), .Y(n27702) );
  XNOR2X1 U45419 ( .A(n51438), .B(n42697), .Y(n27703) );
  NOR4X1 U45420 ( .A(n28001), .B(n28002), .C(n28003), .D(n28004), .Y(n43825)
         );
  NOR4X1 U45421 ( .A(n27580), .B(n27581), .C(n27582), .D(n27583), .Y(n44169)
         );
  NOR4X1 U45422 ( .A(n27490), .B(n27491), .C(n27492), .D(n27493), .Y(n44575)
         );
  XNOR2X1 U45423 ( .A(n50371), .B(n42711), .Y(n27490) );
  XNOR2X1 U45424 ( .A(n50575), .B(n42724), .Y(n27491) );
  XNOR2X1 U45425 ( .A(n51430), .B(n42697), .Y(n27492) );
  NOR4X1 U45426 ( .A(n27610), .B(n27611), .C(n27612), .D(n27613), .Y(net215468) );
  XNOR2X1 U45427 ( .A(n50369), .B(n42711), .Y(n27610) );
  XNOR2X1 U45428 ( .A(n50573), .B(n42724), .Y(n27611) );
  XNOR2X1 U45429 ( .A(n51428), .B(n42697), .Y(n27612) );
  NOR4X1 U45430 ( .A(n27550), .B(n27551), .C(n27552), .D(n27553), .Y(net215432) );
  XNOR2X1 U45431 ( .A(n50367), .B(n42711), .Y(n27550) );
  XNOR2X1 U45432 ( .A(n50571), .B(n42724), .Y(n27551) );
  XNOR2X1 U45433 ( .A(n51426), .B(n42697), .Y(n27552) );
  NOR4X1 U45434 ( .A(n27279), .B(n27280), .C(n27281), .D(n27282), .Y(n44198)
         );
  NOR4X1 U45435 ( .A(n27249), .B(n27250), .C(n27251), .D(n27252), .Y(net215405) );
  XNOR2X1 U45436 ( .A(n50365), .B(n42710), .Y(n27249) );
  XNOR2X1 U45437 ( .A(n50569), .B(n42723), .Y(n27250) );
  XNOR2X1 U45438 ( .A(n51424), .B(n42697), .Y(n27251) );
  XNOR2X1 U45439 ( .A(n50374), .B(n42711), .Y(n27400) );
  XNOR2X1 U45440 ( .A(n50578), .B(n42724), .Y(n27401) );
  XNOR2X1 U45441 ( .A(n51433), .B(n42697), .Y(n27402) );
  NOR4X1 U45442 ( .A(n27460), .B(n27461), .C(n27462), .D(n27463), .Y(n44572)
         );
  XNOR2X1 U45443 ( .A(n50372), .B(n42711), .Y(n27460) );
  XNOR2X1 U45444 ( .A(n50576), .B(n42724), .Y(n27461) );
  XNOR2X1 U45445 ( .A(n51431), .B(n42697), .Y(n27462) );
  XNOR2X1 U45446 ( .A(n50363), .B(n42710), .Y(n27189) );
  XNOR2X1 U45447 ( .A(n50567), .B(n42723), .Y(n27190) );
  NOR4X1 U45448 ( .A(n27219), .B(n27220), .C(n27221), .D(n27222), .Y(net215378) );
  XNOR2X1 U45449 ( .A(n50362), .B(n42710), .Y(n27219) );
  XNOR2X1 U45450 ( .A(n50566), .B(n42723), .Y(n27220) );
  XNOR2X1 U45451 ( .A(n51421), .B(n42697), .Y(n27221) );
  NOR4X1 U45452 ( .A(n27430), .B(n27431), .C(n27432), .D(n27433), .Y(n44178)
         );
  XNOR2X1 U45453 ( .A(n50373), .B(n42711), .Y(n27430) );
  XNOR2X1 U45454 ( .A(n50577), .B(n42724), .Y(n27431) );
  XNOR2X1 U45455 ( .A(n51432), .B(n42697), .Y(n27432) );
  XNOR2X1 U45456 ( .A(n50361), .B(n42710), .Y(n27309) );
  XNOR2X1 U45457 ( .A(n50565), .B(n42723), .Y(n27310) );
  XNOR2X1 U45458 ( .A(n51420), .B(n42697), .Y(n27311) );
  NOR4X1 U45459 ( .A(n27369), .B(n27370), .C(n27371), .D(n27372), .Y(net215369) );
  NOR4X1 U45460 ( .A(n27339), .B(n27340), .C(n27341), .D(n27342), .Y(n44224)
         );
  XNOR2X1 U45461 ( .A(n50359), .B(n42711), .Y(n27339) );
  XNOR2X1 U45462 ( .A(n50563), .B(n42724), .Y(n27340) );
  XNOR2X1 U45463 ( .A(n51418), .B(n42697), .Y(n27341) );
  XOR2X1 U45464 ( .A(n42725), .B(n42061), .Y(n43870) );
  XNOR2X1 U45465 ( .A(n41318), .B(n41806), .Y(n46566) );
  XNOR2X1 U45466 ( .A(n41300), .B(n41798), .Y(n46570) );
  XNOR2X1 U45467 ( .A(n41810), .B(n42526), .Y(n44906) );
  NOR4X1 U45468 ( .A(n29230), .B(n29231), .C(n29232), .D(n29233), .Y(n43579)
         );
  XNOR2X1 U45469 ( .A(n50990), .B(net219314), .Y(n29230) );
  XNOR2X1 U45470 ( .A(n51204), .B(n41282), .Y(n29231) );
  XNOR2X1 U45471 ( .A(n50776), .B(net219468), .Y(n29232) );
  NOR4X1 U45472 ( .A(n28087), .B(n28088), .C(n28089), .D(n28090), .Y(n43815)
         );
  XNOR2X1 U45473 ( .A(n51008), .B(net219336), .Y(n28087) );
  XNOR2X1 U45474 ( .A(n51222), .B(n41282), .Y(n28088) );
  XNOR2X1 U45475 ( .A(n50794), .B(net219468), .Y(n28089) );
  XNOR2X1 U45476 ( .A(n51009), .B(net219310), .Y(n28027) );
  XNOR2X1 U45477 ( .A(n51223), .B(n41283), .Y(n28028) );
  XNOR2X1 U45478 ( .A(n50795), .B(net219466), .Y(n28029) );
  XNOR2X1 U45479 ( .A(n51007), .B(net219308), .Y(n28057) );
  XNOR2X1 U45480 ( .A(n51221), .B(n41281), .Y(n28058) );
  XNOR2X1 U45481 ( .A(n50793), .B(net219468), .Y(n28059) );
  XNOR2X1 U45482 ( .A(n41292), .B(n41803), .Y(n46567) );
  XNOR2X1 U45483 ( .A(n36779), .B(n42059), .Y(n46571) );
  XNOR2X1 U45484 ( .A(n42068), .B(n36873), .Y(n44903) );
  XNOR2X1 U45485 ( .A(n42067), .B(n41322), .Y(n45101) );
  XNOR2X1 U45486 ( .A(n41327), .B(n41800), .Y(n46568) );
  XNOR2X1 U45487 ( .A(n36840), .B(n42062), .Y(n46572) );
  NOR4X1 U45488 ( .A(n27159), .B(n27160), .C(n27161), .D(n27162), .Y(net215385) );
  NOR4X1 U45489 ( .A(n27731), .B(n43846), .C(n43845), .D(n43844), .Y(n43848)
         );
  NAND2X1 U45490 ( .A(n43843), .B(n43842), .Y(n43849) );
  NOR4X1 U45491 ( .A(n44767), .B(n44766), .C(n44765), .D(n44764), .Y(n44783)
         );
  NOR4X1 U45492 ( .A(n44771), .B(n44770), .C(n44769), .D(n44768), .Y(n44782)
         );
  NOR4X1 U45493 ( .A(n27438), .B(n27439), .C(n27440), .D(n27443), .Y(n45678)
         );
  CLKINVX1 U45494 ( .A(net210919), .Y(net209288) );
  CLKINVX1 U45495 ( .A(net210677), .Y(net209944) );
  NOR2X1 U45496 ( .A(n45280), .B(n45279), .Y(n45287) );
  NOR4X1 U45497 ( .A(n45239), .B(n45238), .C(n45237), .D(n45236), .Y(n45254)
         );
  NAND2X1 U45498 ( .A(n48166), .B(n48179), .Y(net210680) );
  NOR4X1 U45499 ( .A(n47648), .B(n47647), .C(n47646), .D(n47645), .Y(net210770) );
  NOR4X1 U45500 ( .A(n47652), .B(n47651), .C(n47650), .D(n47649), .Y(net210771) );
  NAND2X1 U45501 ( .A(n48188), .B(n48133), .Y(n10182) );
  NAND2X1 U45502 ( .A(n11041), .B(n10232), .Y(n11038) );
  NOR4X1 U45503 ( .A(n47671), .B(n47670), .C(n47669), .D(n47668), .Y(n47672)
         );
  XOR2X1 U45504 ( .A(n41317), .B(n41827), .Y(n46445) );
  NOR4X1 U45505 ( .A(n47677), .B(n47676), .C(n47675), .D(n47674), .Y(n47684)
         );
  XOR2X1 U45506 ( .A(n41312), .B(n41829), .Y(n46423) );
  NAND2X1 U45507 ( .A(n11030), .B(n11031), .Y(n11027) );
  XOR2X1 U45508 ( .A(n41311), .B(n41831), .Y(n46401) );
  XOR2X1 U45509 ( .A(n41834), .B(n42522), .Y(n44122) );
  XOR2X1 U45510 ( .A(n41837), .B(n42521), .Y(n43937) );
  NOR2X1 U45511 ( .A(n47532), .B(net209277), .Y(n47542) );
  NOR4X1 U45512 ( .A(n47307), .B(n47306), .C(n47305), .D(n47304), .Y(n47313)
         );
  NOR4X1 U45513 ( .A(n47311), .B(n47310), .C(n47309), .D(n47308), .Y(n47312)
         );
  XOR2X1 U45514 ( .A(n42496), .B(n42077), .Y(n47307) );
  XOR2X1 U45515 ( .A(n36755), .B(n41813), .Y(n47623) );
  XOR2X1 U45516 ( .A(n42512), .B(n41839), .Y(n43999) );
  XOR2X1 U45517 ( .A(n41841), .B(n42524), .Y(n43906) );
  XOR2X1 U45518 ( .A(n41826), .B(n42522), .Y(n44815) );
  NOR2X1 U45519 ( .A(n47543), .B(n48461), .Y(n47551) );
  XOR2X1 U45520 ( .A(n42471), .B(n42058), .Y(n47543) );
  NOR2X1 U45521 ( .A(n47521), .B(net209303), .Y(n47531) );
  XOR2X1 U45522 ( .A(n36753), .B(n41811), .Y(n47612) );
  XOR2X1 U45523 ( .A(n41311), .B(n34351), .Y(n46544) );
  XOR2X1 U45524 ( .A(n41311), .B(n41837), .Y(n46294) );
  XOR2X1 U45525 ( .A(n41316), .B(n41832), .Y(n46412) );
  XOR2X1 U45526 ( .A(n41814), .B(n42515), .Y(n45126) );
  XOR2X1 U45527 ( .A(n34351), .B(n42515), .Y(n45157) );
  XOR2X1 U45528 ( .A(n41827), .B(n42522), .Y(n44784) );
  XNOR2X1 U45529 ( .A(n41798), .B(n36824), .Y(n41765) );
  NAND2X1 U45530 ( .A(n10725), .B(n10726), .Y(n11430) );
  XOR2X1 U45531 ( .A(n41311), .B(n41826), .Y(n46463) );
  NOR2X1 U45532 ( .A(n27720), .B(n27719), .Y(n43843) );
  NOR2X1 U45533 ( .A(n27722), .B(n27721), .Y(n43842) );
  XOR2X1 U45534 ( .A(n41311), .B(n41818), .Y(n46310) );
  NAND2X1 U45535 ( .A(n41766), .B(n41767), .Y(n45677) );
  XNOR2X1 U45536 ( .A(n42110), .B(n36877), .Y(n41766) );
  XNOR2X1 U45537 ( .A(n41851), .B(n42526), .Y(n41767) );
  XNOR2X1 U45538 ( .A(n42111), .B(n41323), .Y(n41768) );
  CLKBUFX3 U45539 ( .A(n42514), .Y(n42511) );
  CLKBUFX3 U45540 ( .A(n42482), .Y(n42481) );
  CLKBUFX3 U45541 ( .A(n42458), .Y(n42457) );
  XNOR2X1 U45542 ( .A(n51414), .B(n42693), .Y(n29146) );
  XNOR2X1 U45543 ( .A(n50559), .B(n41379), .Y(n29167) );
  XNOR2X1 U45544 ( .A(n50354), .B(n36907), .Y(n29136) );
  XOR2X1 U45545 ( .A(n41865), .B(n36901), .Y(n29173) );
  XOR2X1 U45546 ( .A(n41866), .B(n36894), .Y(n29143) );
  XOR2X1 U45547 ( .A(n42126), .B(n42652), .Y(n29139) );
  XOR2X1 U45548 ( .A(n42125), .B(n36885), .Y(n29147) );
  XNOR2X1 U45549 ( .A(n51201), .B(n41283), .Y(n29141) );
  XNOR2X1 U45550 ( .A(n50988), .B(net219310), .Y(n29170) );
  XOR2X1 U45551 ( .A(n42140), .B(n42661), .Y(n26762) );
  XOR2X1 U45552 ( .A(n41880), .B(n36898), .Y(n26766) );
  XNOR2X1 U45553 ( .A(n50558), .B(n36905), .Y(n29137) );
  XOR2X1 U45554 ( .A(n41881), .B(n42607), .Y(n26758) );
  XOR2X1 U45555 ( .A(n42139), .B(n36879), .Y(n26770) );
  XNOR2X1 U45556 ( .A(n50341), .B(n42708), .Y(n26767) );
  XNOR2X1 U45557 ( .A(n50356), .B(n41642), .Y(n29174) );
  XNOR2X1 U45558 ( .A(n50340), .B(n42672), .Y(n26759) );
  XNOR2X1 U45559 ( .A(n50987), .B(n36870), .Y(n29140) );
  NAND4X1 U45560 ( .A(n43601), .B(n43600), .C(n43599), .D(n43598), .Y(n43606)
         );
  OAI21XL U45561 ( .A0(n48445), .A1(n48444), .B0(n48443), .Y(n48450) );
  XNOR2X1 U45562 ( .A(n50354), .B(n41642), .Y(n29324) );
  XNOR2X1 U45563 ( .A(n50357), .B(n42705), .Y(n29204) );
  XNOR2X1 U45564 ( .A(n50353), .B(n42704), .Y(n29354) );
  XNOR2X1 U45565 ( .A(n50556), .B(n42717), .Y(n29265) );
  XNOR2X1 U45566 ( .A(n50553), .B(n42724), .Y(n29385) );
  XNOR2X1 U45567 ( .A(n50555), .B(n42718), .Y(n29295) );
  XNOR2X1 U45568 ( .A(n50984), .B(n41297), .Y(n22396) );
  XNOR2X1 U45569 ( .A(n50999), .B(n41297), .Y(n23994) );
  XNOR2X1 U45570 ( .A(n51008), .B(n36791), .Y(n20286) );
  XNOR2X1 U45571 ( .A(n51007), .B(n36790), .Y(n20296) );
  XNOR2X1 U45572 ( .A(n50995), .B(n36795), .Y(n20152) );
  XNOR2X1 U45573 ( .A(n51004), .B(n36796), .Y(n20214) );
  XNOR2X1 U45574 ( .A(n50998), .B(n41293), .Y(n24004) );
  XNOR2X1 U45575 ( .A(n50996), .B(n36916), .Y(n23753) );
  XNOR2X1 U45576 ( .A(n50985), .B(n41297), .Y(n22436) );
  XNOR2X1 U45577 ( .A(n50992), .B(n36799), .Y(n20111) );
  XNOR2X1 U45578 ( .A(n50574), .B(n42582), .Y(n27443) );
  XNOR2X1 U45579 ( .A(n50974), .B(n42534), .Y(n29031) );
  XNOR2X1 U45580 ( .A(n50975), .B(n42534), .Y(n29091) );
  XNOR2X1 U45581 ( .A(n50997), .B(n42542), .Y(n27528) );
  XNOR2X1 U45582 ( .A(n50573), .B(n42582), .Y(n27473) );
  XNOR2X1 U45583 ( .A(n50993), .B(n42541), .Y(n27167) );
  XNOR2X1 U45584 ( .A(n51413), .B(n42693), .Y(n29326) );
  XNOR2X1 U45585 ( .A(n51416), .B(n42693), .Y(n29206) );
  XNOR2X1 U45586 ( .A(n51412), .B(n42693), .Y(n29356) );
  XNOR2X1 U45587 ( .A(n51406), .B(n42696), .Y(n29446) );
  XNOR2X1 U45588 ( .A(n51405), .B(n42695), .Y(n29085) );
  XNOR2X1 U45589 ( .A(n51198), .B(n41330), .Y(n22397) );
  XNOR2X1 U45590 ( .A(n51213), .B(n41327), .Y(n23995) );
  XNOR2X1 U45591 ( .A(n51222), .B(n36715), .Y(n20287) );
  XNOR2X1 U45592 ( .A(n51221), .B(n36714), .Y(n20297) );
  XNOR2X1 U45593 ( .A(n51209), .B(n36714), .Y(n20153) );
  XNOR2X1 U45594 ( .A(n51218), .B(n36715), .Y(n20215) );
  XNOR2X1 U45595 ( .A(n51212), .B(n41332), .Y(n24005) );
  XNOR2X1 U45596 ( .A(n51210), .B(n41327), .Y(n23754) );
  XNOR2X1 U45597 ( .A(n51199), .B(n36913), .Y(n22437) );
  XNOR2X1 U45598 ( .A(n51206), .B(n36716), .Y(n20112) );
  XNOR2X1 U45599 ( .A(n50788), .B(n42506), .Y(n27440) );
  XNOR2X1 U45600 ( .A(n50781), .B(net219442), .Y(n27187) );
  XNOR2X1 U45601 ( .A(n51421), .B(n42641), .Y(n27183) );
  XNOR2X1 U45602 ( .A(n50780), .B(n36863), .Y(n27179) );
  XNOR2X1 U45603 ( .A(n51187), .B(n42549), .Y(n29002) );
  XNOR2X1 U45604 ( .A(n51192), .B(n42552), .Y(n29453) );
  XNOR2X1 U45605 ( .A(n51211), .B(n42551), .Y(n27529) );
  XNOR2X1 U45606 ( .A(n51405), .B(n36867), .Y(n29438) );
  XNOR2X1 U45607 ( .A(n50764), .B(n42586), .Y(n29434) );
  XNOR2X1 U45608 ( .A(n51402), .B(n42644), .Y(n29047) );
  XNOR2X1 U45609 ( .A(n51403), .B(n42643), .Y(n29107) );
  XNOR2X1 U45610 ( .A(n50762), .B(n34450), .Y(n29103) );
  XNOR2X1 U45611 ( .A(n50761), .B(n42592), .Y(n29043) );
  XNOR2X1 U45612 ( .A(n51400), .B(n36867), .Y(n26791) );
  XNOR2X1 U45613 ( .A(n50759), .B(n36865), .Y(n26787) );
  XNOR2X1 U45614 ( .A(n50756), .B(net219434), .Y(n26855) );
  XNOR2X1 U45615 ( .A(n50757), .B(net219434), .Y(n26705) );
  XNOR2X1 U45616 ( .A(n51397), .B(n36867), .Y(n26701) );
  XNOR2X1 U45617 ( .A(n50756), .B(n36865), .Y(n26697) );
  XNOR2X1 U45618 ( .A(n50787), .B(n36737), .Y(n27470) );
  XNOR2X1 U45619 ( .A(n51207), .B(n42552), .Y(n27168) );
  XNOR2X1 U45620 ( .A(n50753), .B(net219442), .Y(n26675) );
  XNOR2X1 U45621 ( .A(n51393), .B(n36867), .Y(n26671) );
  XNOR2X1 U45622 ( .A(n50551), .B(n42718), .Y(n29445) );
  XNOR2X1 U45623 ( .A(n50550), .B(n42724), .Y(n29084) );
  XNOR2X1 U45624 ( .A(n50770), .B(n36850), .Y(n22398) );
  XNOR2X1 U45625 ( .A(n50785), .B(n36860), .Y(n23996) );
  XNOR2X1 U45626 ( .A(n50794), .B(n42469), .Y(n20288) );
  XNOR2X1 U45627 ( .A(n50793), .B(n42469), .Y(n20298) );
  XNOR2X1 U45628 ( .A(n50781), .B(n42468), .Y(n20154) );
  XNOR2X1 U45629 ( .A(n50790), .B(n42469), .Y(n20216) );
  XNOR2X1 U45630 ( .A(n50784), .B(n36854), .Y(n24006) );
  XNOR2X1 U45631 ( .A(n50782), .B(n36851), .Y(n23755) );
  XNOR2X1 U45632 ( .A(n50771), .B(n36860), .Y(n22438) );
  XNOR2X1 U45633 ( .A(n50778), .B(n42468), .Y(n20113) );
  XNOR2X1 U45634 ( .A(n50972), .B(net219308), .Y(n26733) );
  XNOR2X1 U45635 ( .A(n50339), .B(n42670), .Y(n26729) );
  XNOR2X1 U45636 ( .A(n50362), .B(n42674), .Y(n27181) );
  XNOR2X1 U45637 ( .A(n50994), .B(n42615), .Y(n27177) );
  XNOR2X1 U45638 ( .A(n50988), .B(n41284), .Y(n29192) );
  XNOR2X1 U45639 ( .A(n50347), .B(n41642), .Y(n29444) );
  XNOR2X1 U45640 ( .A(n50346), .B(n42671), .Y(n29436) );
  XNOR2X1 U45641 ( .A(n50978), .B(n42615), .Y(n29432) );
  XNOR2X1 U45642 ( .A(n50346), .B(n42707), .Y(n29083) );
  XNOR2X1 U45643 ( .A(n50345), .B(n42671), .Y(n29075) );
  XNOR2X1 U45644 ( .A(n50977), .B(n42614), .Y(n29071) );
  XNOR2X1 U45645 ( .A(n50975), .B(n42620), .Y(n29041) );
  XNOR2X1 U45646 ( .A(n50341), .B(n42670), .Y(n26789) );
  XNOR2X1 U45647 ( .A(n50973), .B(n42613), .Y(n26785) );
  XNOR2X1 U45648 ( .A(n50337), .B(n42670), .Y(n26849) );
  XNOR2X1 U45649 ( .A(n50969), .B(n42615), .Y(n26845) );
  XNOR2X1 U45650 ( .A(n50971), .B(n40039), .Y(n26703) );
  XNOR2X1 U45651 ( .A(n50338), .B(n42670), .Y(n26699) );
  XNOR2X1 U45652 ( .A(n50970), .B(n42615), .Y(n26695) );
  XNOR2X1 U45653 ( .A(n50984), .B(n41284), .Y(n29342) );
  XNOR2X1 U45654 ( .A(n51216), .B(n42550), .Y(n27439) );
  XNOR2X1 U45655 ( .A(n51186), .B(n41281), .Y(n26734) );
  XNOR2X1 U45656 ( .A(n50774), .B(n42502), .Y(n29214) );
  XNOR2X1 U45657 ( .A(n51209), .B(n41283), .Y(n27186) );
  XNOR2X1 U45658 ( .A(n50566), .B(n36834), .Y(n27182) );
  XNOR2X1 U45659 ( .A(n51208), .B(n42633), .Y(n27178) );
  XNOR2X1 U45660 ( .A(n50560), .B(n41319), .Y(n29197) );
  XNOR2X1 U45661 ( .A(n50769), .B(n42502), .Y(n29334) );
  XNOR2X1 U45662 ( .A(n50770), .B(n42502), .Y(n29304) );
  XNOR2X1 U45663 ( .A(n50783), .B(n36737), .Y(n27530) );
  XNOR2X1 U45664 ( .A(n50550), .B(n36728), .Y(n29437) );
  XNOR2X1 U45665 ( .A(n51192), .B(n42633), .Y(n29433) );
  XNOR2X1 U45666 ( .A(n50549), .B(n41319), .Y(n29076) );
  XNOR2X1 U45667 ( .A(n51190), .B(n42632), .Y(n29102) );
  XNOR2X1 U45668 ( .A(n50548), .B(n42725), .Y(n29054) );
  XNOR2X1 U45669 ( .A(n50547), .B(n36905), .Y(n29046) );
  XNOR2X1 U45670 ( .A(n51189), .B(n42624), .Y(n29042) );
  XNOR2X1 U45671 ( .A(n50545), .B(n36905), .Y(n26790) );
  XNOR2X1 U45672 ( .A(n51187), .B(n42633), .Y(n26786) );
  XNOR2X1 U45673 ( .A(n51184), .B(n41282), .Y(n26854) );
  XNOR2X1 U45674 ( .A(n50541), .B(n36905), .Y(n26850) );
  XNOR2X1 U45675 ( .A(n51185), .B(n41281), .Y(n26704) );
  XNOR2X1 U45676 ( .A(n50542), .B(n41319), .Y(n26700) );
  XNOR2X1 U45677 ( .A(n51184), .B(n42633), .Y(n26696) );
  XNOR2X1 U45678 ( .A(n51215), .B(n36832), .Y(n27469) );
  XNOR2X1 U45679 ( .A(n50556), .B(n36905), .Y(n29347) );
  XOR2X1 U45680 ( .A(n42123), .B(n42653), .Y(n29229) );
  XOR2X1 U45681 ( .A(n41864), .B(n42602), .Y(n29225) );
  XOR2X1 U45682 ( .A(n42140), .B(n36888), .Y(n26740) );
  XOR2X1 U45683 ( .A(n41881), .B(n36901), .Y(n26736) );
  XOR2X1 U45684 ( .A(n42141), .B(n42661), .Y(n26732) );
  XOR2X1 U45685 ( .A(n41882), .B(n42607), .Y(n26728) );
  XOR2X1 U45686 ( .A(n42126), .B(n36889), .Y(n29327) );
  XOR2X1 U45687 ( .A(n42127), .B(n42653), .Y(n29319) );
  XOR2X1 U45688 ( .A(n42147), .B(n36886), .Y(n26951) );
  XOR2X1 U45689 ( .A(n42118), .B(n42662), .Y(n27184) );
  XOR2X1 U45690 ( .A(n41859), .B(n42608), .Y(n27180) );
  XOR2X1 U45691 ( .A(n41864), .B(n36900), .Y(n29203) );
  XOR2X1 U45692 ( .A(n42123), .B(n36887), .Y(n29207) );
  XOR2X1 U45693 ( .A(n42124), .B(n42652), .Y(n29199) );
  XOR2X1 U45694 ( .A(n41865), .B(n42601), .Y(n29195) );
  XOR2X1 U45695 ( .A(n41878), .B(n42601), .Y(n29044) );
  XOR2X1 U45696 ( .A(n42138), .B(n36879), .Y(n26800) );
  XOR2X1 U45697 ( .A(n42139), .B(n42661), .Y(n26792) );
  XOR2X1 U45698 ( .A(n41880), .B(n42607), .Y(n26788) );
  XOR2X1 U45699 ( .A(n42142), .B(n36880), .Y(n26860) );
  XOR2X1 U45700 ( .A(n41883), .B(n36895), .Y(n26856) );
  XOR2X1 U45701 ( .A(n42143), .B(n42661), .Y(n26852) );
  XOR2X1 U45702 ( .A(n41884), .B(n42607), .Y(n26848) );
  XOR2X1 U45703 ( .A(n42141), .B(n36888), .Y(n26710) );
  XOR2X1 U45704 ( .A(n41882), .B(n36894), .Y(n26706) );
  XOR2X1 U45705 ( .A(n42142), .B(n42661), .Y(n26702) );
  XOR2X1 U45706 ( .A(n41883), .B(n42607), .Y(n26698) );
  XOR2X1 U45707 ( .A(n41886), .B(n36892), .Y(n26676) );
  XOR2X1 U45708 ( .A(n42146), .B(n42663), .Y(n26672) );
  XOR2X1 U45709 ( .A(n41887), .B(n42608), .Y(n26668) );
  XOR2X1 U45710 ( .A(n41868), .B(n36897), .Y(n29353) );
  XOR2X1 U45711 ( .A(n42127), .B(n36881), .Y(n29357) );
  XOR2X1 U45712 ( .A(n42128), .B(n42653), .Y(n29349) );
  XOR2X1 U45713 ( .A(n41869), .B(n42602), .Y(n29345) );
  XOR2X1 U45714 ( .A(n41866), .B(n42516), .Y(n29185) );
  XOR2X1 U45715 ( .A(n36773), .B(n42061), .Y(n47546) );
  XOR2X1 U45716 ( .A(n41869), .B(n41316), .Y(n22399) );
  XOR2X1 U45717 ( .A(n41845), .B(n36760), .Y(n20289) );
  XOR2X1 U45718 ( .A(n41840), .B(n36760), .Y(n20381) );
  XOR2X1 U45719 ( .A(n41845), .B(n41311), .Y(n23817) );
  XOR2X1 U45720 ( .A(n41858), .B(n36757), .Y(n20155) );
  XOR2X1 U45721 ( .A(n41855), .B(n41316), .Y(n24007) );
  XOR2X1 U45722 ( .A(n41857), .B(n41314), .Y(n23756) );
  XOR2X1 U45723 ( .A(n41861), .B(n36757), .Y(n20114) );
  XOR2X1 U45724 ( .A(n42099), .B(n42478), .Y(n20382) );
  XOR2X1 U45725 ( .A(n36770), .B(n42060), .Y(n47537) );
  XNOR2X1 U45726 ( .A(n51411), .B(n41303), .Y(n22401) );
  XNOR2X1 U45727 ( .A(n50566), .B(n36766), .Y(n20167) );
  XNOR2X1 U45728 ( .A(n51412), .B(n41304), .Y(n22441) );
  XNOR2X1 U45729 ( .A(n51414), .B(n41303), .Y(n22461) );
  XNOR2X1 U45730 ( .A(n51423), .B(n36748), .Y(n20147) );
  XNOR2X1 U45731 ( .A(n51438), .B(n36741), .Y(n20413) );
  XNOR2X1 U45732 ( .A(n50567), .B(n36773), .Y(n20157) );
  XNOR2X1 U45733 ( .A(n50565), .B(n36783), .Y(n23708) );
  XNOR2X1 U45734 ( .A(n50576), .B(n36768), .Y(n20219) );
  XNOR2X1 U45735 ( .A(n50564), .B(n36776), .Y(n23718) );
  XNOR2X1 U45736 ( .A(n51423), .B(n41305), .Y(n23758) );
  XNOR2X1 U45737 ( .A(n50577), .B(n36768), .Y(n20281) );
  XNOR2X1 U45738 ( .A(n50985), .B(n42535), .Y(n29122) );
  XNOR2X1 U45739 ( .A(n50565), .B(n42581), .Y(n27172) );
  XOR2X1 U45740 ( .A(n42128), .B(n36809), .Y(n22400) );
  XOR2X1 U45741 ( .A(n42104), .B(n36808), .Y(n23818) );
  XOR2X1 U45742 ( .A(n42117), .B(n42492), .Y(n20156) );
  XOR2X1 U45743 ( .A(n42116), .B(n36810), .Y(n23757) );
  XOR2X1 U45744 ( .A(n42127), .B(n36815), .Y(n22440) );
  XOR2X1 U45745 ( .A(n36792), .B(n41804), .Y(n47533) );
  XOR2X1 U45746 ( .A(n36722), .B(n41801), .Y(n47534) );
  NOR4X1 U45747 ( .A(n19606), .B(n19605), .C(n19604), .D(n19603), .Y(n47239)
         );
  NOR4X1 U45748 ( .A(n19596), .B(n19595), .C(n19594), .D(n19593), .Y(n47244)
         );
  XOR2X1 U45749 ( .A(n41866), .B(n36757), .Y(n19596) );
  XNOR2X1 U45750 ( .A(n50773), .B(n42465), .Y(n19595) );
  XNOR2X1 U45751 ( .A(n51201), .B(n36714), .Y(n19594) );
  XNOR2X1 U45752 ( .A(n50333), .B(n42710), .Y(n26948) );
  XNOR2X1 U45753 ( .A(n50537), .B(n42723), .Y(n26949) );
  XNOR2X1 U45754 ( .A(n51392), .B(n42697), .Y(n26950) );
  NOR4X1 U45755 ( .A(n26857), .B(n26858), .C(n26859), .D(n26860), .Y(n44309)
         );
  XNOR2X1 U45756 ( .A(n50338), .B(n42707), .Y(n26857) );
  NOR4X1 U45757 ( .A(n26707), .B(n26708), .C(n26709), .D(n26710), .Y(n44607)
         );
  XNOR2X1 U45758 ( .A(n50339), .B(n41641), .Y(n26707) );
  XNOR2X1 U45759 ( .A(n50543), .B(n34435), .Y(n26708) );
  XNOR2X1 U45760 ( .A(n51398), .B(n42696), .Y(n26709) );
  XNOR2X1 U45761 ( .A(n50335), .B(n42708), .Y(n26677) );
  XNOR2X1 U45762 ( .A(n50539), .B(n42717), .Y(n26678) );
  XNOR2X1 U45763 ( .A(n50337), .B(n41641), .Y(n26887) );
  XNOR2X1 U45764 ( .A(n50541), .B(n36875), .Y(n26888) );
  XNOR2X1 U45765 ( .A(n51396), .B(n42697), .Y(n26889) );
  NOR4X1 U45766 ( .A(n26918), .B(n26919), .C(n26920), .D(n26921), .Y(net215279) );
  NOR4X1 U45767 ( .A(n26737), .B(n26738), .C(n26739), .D(n26740), .Y(n44603)
         );
  XNOR2X1 U45768 ( .A(n50340), .B(n42707), .Y(n26737) );
  XNOR2X1 U45769 ( .A(n50544), .B(n42717), .Y(n26738) );
  XNOR2X1 U45770 ( .A(n51399), .B(n42696), .Y(n26739) );
  NOR4X1 U45771 ( .A(n26797), .B(n26798), .C(n26799), .D(n26800), .Y(n44278)
         );
  XNOR2X1 U45772 ( .A(n50342), .B(n41642), .Y(n26797) );
  XNOR2X1 U45773 ( .A(n50546), .B(n34435), .Y(n26798) );
  XNOR2X1 U45774 ( .A(n51401), .B(n42696), .Y(n26799) );
  NOR4X1 U45775 ( .A(n27008), .B(n27009), .C(n27010), .D(n27011), .Y(n44268)
         );
  XNOR2X1 U45776 ( .A(n50331), .B(n42710), .Y(n27008) );
  XNOR2X1 U45777 ( .A(n50535), .B(n42723), .Y(n27009) );
  XNOR2X1 U45778 ( .A(n51390), .B(n42697), .Y(n27010) );
  NOR4X1 U45779 ( .A(n27098), .B(n27099), .C(n27100), .D(n27101), .Y(net215315) );
  NOR4X1 U45780 ( .A(n27038), .B(n27039), .C(n27040), .D(n27041), .Y(n44243)
         );
  XNOR2X1 U45781 ( .A(n50328), .B(n42710), .Y(n27038) );
  XNOR2X1 U45782 ( .A(n50532), .B(n42723), .Y(n27039) );
  XNOR2X1 U45783 ( .A(n51387), .B(n42697), .Y(n27040) );
  NOR4X1 U45784 ( .A(n27128), .B(n27129), .C(n27130), .D(n27131), .Y(n44252)
         );
  XNOR2X1 U45785 ( .A(n50329), .B(n42710), .Y(n27128) );
  XNOR2X1 U45786 ( .A(n50533), .B(n42723), .Y(n27129) );
  XNOR2X1 U45787 ( .A(n51388), .B(n42697), .Y(n27130) );
  XNOR2X1 U45788 ( .A(n50986), .B(net219314), .Y(n29320) );
  NOR4X1 U45789 ( .A(n29260), .B(n29261), .C(n29262), .D(n29263), .Y(n43626)
         );
  NOR4X1 U45790 ( .A(n29470), .B(n29471), .C(n29472), .D(n29473), .Y(n43547)
         );
  NOR4X1 U45791 ( .A(n29380), .B(n29381), .C(n29382), .D(n29383), .Y(n43570)
         );
  XNOR2X1 U45792 ( .A(n51195), .B(n41282), .Y(n29381) );
  XNOR2X1 U45793 ( .A(n50767), .B(net258207), .Y(n29382) );
  NOR4X1 U45794 ( .A(n29200), .B(n29201), .C(n29202), .D(n29203), .Y(n43588)
         );
  XNOR2X1 U45795 ( .A(n50989), .B(net219336), .Y(n29200) );
  XNOR2X1 U45796 ( .A(n51203), .B(n41282), .Y(n29201) );
  XNOR2X1 U45797 ( .A(n50775), .B(net258207), .Y(n29202) );
  XNOR2X1 U45798 ( .A(n50979), .B(net219330), .Y(n29440) );
  XNOR2X1 U45799 ( .A(n51193), .B(n41283), .Y(n29441) );
  NOR4X1 U45800 ( .A(n29079), .B(n29080), .C(n29081), .D(n29082), .Y(n43654)
         );
  XNOR2X1 U45801 ( .A(n50978), .B(net219310), .Y(n29079) );
  XNOR2X1 U45802 ( .A(n51192), .B(n41282), .Y(n29080) );
  XNOR2X1 U45803 ( .A(n50764), .B(net219468), .Y(n29081) );
  XNOR2X1 U45804 ( .A(n51190), .B(n41282), .Y(n29050) );
  NOR4X1 U45805 ( .A(n29350), .B(n29351), .C(n29352), .D(n29353), .Y(net216045) );
  XNOR2X1 U45806 ( .A(n51199), .B(n41282), .Y(n29351) );
  XNOR2X1 U45807 ( .A(n50771), .B(net219468), .Y(n29352) );
  XNOR2X1 U45808 ( .A(n50983), .B(net219314), .Y(n29290) );
  XNOR2X1 U45809 ( .A(n51197), .B(n41282), .Y(n29291) );
  XNOR2X1 U45810 ( .A(n50769), .B(net258207), .Y(n29292) );
  NOR4X1 U45811 ( .A(n29410), .B(n29411), .C(n29412), .D(n29413), .Y(net216137) );
  NOR4X1 U45812 ( .A(n26978), .B(n26979), .C(n26980), .D(n26981), .Y(net215304) );
  XOR2X1 U45813 ( .A(n42141), .B(n41322), .Y(n26749) );
  NOR4X1 U45814 ( .A(n29019), .B(n29020), .C(n29021), .D(n29022), .Y(n43672)
         );
  AOI21X1 U45815 ( .A0(n48459), .A1(n48458), .B0(n48457), .Y(n48473) );
  CLKINVX1 U45816 ( .A(n12386), .Y(net171418) );
  XNOR2X1 U45817 ( .A(n50557), .B(n42577), .Y(n29127) );
  NOR3X1 U45818 ( .A(n29172), .B(n29170), .C(n29154), .Y(n43598) );
  CLKINVX1 U45819 ( .A(n10487), .Y(net209736) );
  AOI21X1 U45820 ( .A0(n48534), .A1(n10820), .B0(net209179), .Y(n48535) );
  OAI221XL U45821 ( .A0(n10233), .A1(n10231), .B0(n10232), .B1(net209182),
        .C0(n11039), .Y(n48532) );
  NOR2X1 U45822 ( .A(n29184), .B(n29187), .Y(n43594) );
  NOR2X1 U45823 ( .A(n29182), .B(n29183), .Y(n43593) );
  CLKINVX1 U45824 ( .A(n10903), .Y(net209144) );
  CLKINVX1 U45825 ( .A(n11034), .Y(net209175) );
  CLKINVX1 U45826 ( .A(n11217), .Y(net209161) );
  AOI21X1 U45827 ( .A0(n48248), .A1(n12006), .B0(net209781), .Y(n48249) );
  CLKINVX1 U45828 ( .A(n11007), .Y(net209158) );
  XNOR2X1 U45829 ( .A(n50971), .B(n42540), .Y(n26745) );
  AOI21X1 U45830 ( .A0(n48170), .A1(n48169), .B0(n48168), .Y(n48193) );
  AOI21X1 U45831 ( .A0(n48480), .A1(n48479), .B0(n48478), .Y(n48490) );
  NAND4BBXL U45832 ( .AN(n48494), .BN(n48493), .C(n48492), .D(n48491), .Y(
        n48495) );
  AOI21X1 U45833 ( .A0(n48425), .A1(n12385), .B0(net209355), .Y(n48497) );
  AOI21X1 U45834 ( .A0(n48516), .A1(n48515), .B0(n48514), .Y(n48526) );
  AOI21X1 U45835 ( .A0(n48200), .A1(n48199), .B0(n48198), .Y(n48211) );
  NAND2X1 U45836 ( .A(n48197), .B(n48196), .Y(n48198) );
  CLKINVX1 U45837 ( .A(n12723), .Y(net151758) );
  CLKINVX1 U45838 ( .A(n12940), .Y(net151744) );
  CLKINVX1 U45839 ( .A(n12333), .Y(net171482) );
  NOR4X1 U45840 ( .A(n44292), .B(n26760), .C(n26764), .D(n26768), .Y(n44301)
         );
  CLKINVX1 U45841 ( .A(n12942), .Y(net151746) );
  XOR2X1 U45842 ( .A(n42127), .B(n36873), .Y(n29126) );
  NOR2X1 U45843 ( .A(n29156), .B(n29173), .Y(n43597) );
  NAND2X1 U45844 ( .A(n43616), .B(n43615), .Y(n43617) );
  XNOR2X1 U45845 ( .A(n50771), .B(n42501), .Y(n29124) );
  XNOR2X1 U45846 ( .A(n50543), .B(n42577), .Y(n26750) );
  OR2X1 U45847 ( .A(n41774), .B(n29157), .Y(n43604) );
  OR2X1 U45848 ( .A(n29164), .B(n29171), .Y(n41774) );
  XNOR2X1 U45849 ( .A(n50558), .B(n42577), .Y(n29157) );
  XNOR2X1 U45850 ( .A(n51199), .B(n36832), .Y(n29123) );
  CLKBUFX3 U45851 ( .A(n42482), .Y(n42480) );
  CLKINVX1 U45852 ( .A(net209311), .Y(net209310) );
  NOR4X1 U45853 ( .A(n25122), .B(n25123), .C(n25124), .D(n25127), .Y(n44450)
         );
  NOR4X1 U45854 ( .A(n44449), .B(n44448), .C(n25126), .D(n25125), .Y(n44451)
         );
  XNOR2X1 U45855 ( .A(n50954), .B(n42539), .Y(n25122) );
  NOR2X1 U45856 ( .A(n44571), .B(n44465), .Y(n44466) );
  NAND3X1 U45857 ( .A(n44464), .B(n44463), .C(n44462), .Y(n44465) );
  CLKINVX1 U45858 ( .A(net210099), .Y(net171538) );
  CLKINVX1 U45859 ( .A(n10243), .Y(net171458) );
  CLKINVX1 U45860 ( .A(n10530), .Y(net171205) );
  NAND3X1 U45861 ( .A(n22879), .B(n22880), .C(n22882), .Y(n45951) );
  XNOR2X1 U45862 ( .A(n50939), .B(n41291), .Y(n23213) );
  XNOR2X1 U45863 ( .A(n50974), .B(n41291), .Y(n22346) );
  XNOR2X1 U45864 ( .A(n50961), .B(n41292), .Y(n24096) );
  XNOR2X1 U45865 ( .A(n50964), .B(n36789), .Y(n19796) );
  XNOR2X1 U45866 ( .A(n50962), .B(n36791), .Y(n19786) );
  XNOR2X1 U45867 ( .A(n50960), .B(n36792), .Y(n19736) );
  XNOR2X1 U45868 ( .A(n50938), .B(n41296), .Y(n23203) );
  XNOR2X1 U45869 ( .A(n50964), .B(n41294), .Y(n24126) );
  XNOR2X1 U45870 ( .A(n50945), .B(n41294), .Y(n23600) );
  XNOR2X1 U45871 ( .A(n50984), .B(n36789), .Y(n19543) );
  XNOR2X1 U45872 ( .A(n50940), .B(n42543), .Y(n28130) );
  XNOR2X1 U45873 ( .A(n50934), .B(n42536), .Y(n28550) );
  XNOR2X1 U45874 ( .A(n51369), .B(n42698), .Y(n28154) );
  XNOR2X1 U45875 ( .A(n51352), .B(n42701), .Y(n31553) );
  XNOR2X1 U45876 ( .A(n51153), .B(n41327), .Y(n23214) );
  XNOR2X1 U45877 ( .A(n51188), .B(n41329), .Y(n22347) );
  XNOR2X1 U45878 ( .A(n51175), .B(n41331), .Y(n24097) );
  XNOR2X1 U45879 ( .A(n51178), .B(n36720), .Y(n19797) );
  XNOR2X1 U45880 ( .A(n51176), .B(n36715), .Y(n19787) );
  XNOR2X1 U45881 ( .A(n51174), .B(n36714), .Y(n19737) );
  XNOR2X1 U45882 ( .A(n51152), .B(n41327), .Y(n23204) );
  XNOR2X1 U45883 ( .A(n51178), .B(n41328), .Y(n24127) );
  XNOR2X1 U45884 ( .A(n51159), .B(n41327), .Y(n23601) );
  XNOR2X1 U45885 ( .A(n51198), .B(n36718), .Y(n19544) );
  XNOR2X1 U45886 ( .A(n50732), .B(net219468), .Y(n24782) );
  XNOR2X1 U45887 ( .A(n51376), .B(n42641), .Y(n24868) );
  XNOR2X1 U45888 ( .A(n50735), .B(n42586), .Y(n24864) );
  XNOR2X1 U45889 ( .A(n50731), .B(net219468), .Y(n24752) );
  XNOR2X1 U45890 ( .A(n51368), .B(n42643), .Y(n28146) );
  XNOR2X1 U45891 ( .A(n50727), .B(n42587), .Y(n28142) );
  XNOR2X1 U45892 ( .A(n50729), .B(net219468), .Y(n24812) );
  XNOR2X1 U45893 ( .A(n51351), .B(n36867), .Y(n31545) );
  XNOR2X1 U45894 ( .A(n50710), .B(n36865), .Y(n31541) );
  XNOR2X1 U45895 ( .A(n50740), .B(net219434), .Y(n24992) );
  XNOR2X1 U45896 ( .A(n51380), .B(n36861), .Y(n24988) );
  XNOR2X1 U45897 ( .A(n50739), .B(n36865), .Y(n24984) );
  XNOR2X1 U45898 ( .A(n51154), .B(n42553), .Y(n28131) );
  XNOR2X1 U45899 ( .A(n51148), .B(n42548), .Y(n28551) );
  XNOR2X1 U45900 ( .A(n50752), .B(n36865), .Y(n26667) );
  XNOR2X1 U45901 ( .A(n50497), .B(n41287), .Y(n31552) );
  XNOR2X1 U45902 ( .A(n50725), .B(n36857), .Y(n23215) );
  XNOR2X1 U45903 ( .A(n50760), .B(n36858), .Y(n22348) );
  XNOR2X1 U45904 ( .A(n50747), .B(n36850), .Y(n24098) );
  XNOR2X1 U45905 ( .A(n50750), .B(n42466), .Y(n19798) );
  XNOR2X1 U45906 ( .A(n50748), .B(n42476), .Y(n19788) );
  XNOR2X1 U45907 ( .A(n50746), .B(n42465), .Y(n19738) );
  XNOR2X1 U45908 ( .A(n50724), .B(n36850), .Y(n23205) );
  XNOR2X1 U45909 ( .A(n50750), .B(n36852), .Y(n24128) );
  XNOR2X1 U45910 ( .A(n50731), .B(n36850), .Y(n23602) );
  XNOR2X1 U45911 ( .A(n50770), .B(n42465), .Y(n19545) );
  XNOR2X1 U45912 ( .A(n50950), .B(net219308), .Y(n24870) );
  XNOR2X1 U45913 ( .A(n50317), .B(n42672), .Y(n24866) );
  XNOR2X1 U45914 ( .A(n50949), .B(n42615), .Y(n24862) );
  XNOR2X1 U45915 ( .A(n50310), .B(n42712), .Y(n28152) );
  XNOR2X1 U45916 ( .A(n50309), .B(n42671), .Y(n28144) );
  XNOR2X1 U45917 ( .A(n50941), .B(n42619), .Y(n28140) );
  XNOR2X1 U45918 ( .A(n50293), .B(n42708), .Y(n31551) );
  XNOR2X1 U45919 ( .A(n50292), .B(n42670), .Y(n31543) );
  XNOR2X1 U45920 ( .A(n50924), .B(n42617), .Y(n31539) );
  XNOR2X1 U45921 ( .A(n50954), .B(net219314), .Y(n24990) );
  XNOR2X1 U45922 ( .A(n50321), .B(n42673), .Y(n24986) );
  XNOR2X1 U45923 ( .A(n50953), .B(n42613), .Y(n24982) );
  XNOR2X1 U45924 ( .A(n50967), .B(net219310), .Y(n26673) );
  XNOR2X1 U45925 ( .A(n50334), .B(n36907), .Y(n26669) );
  XNOR2X1 U45926 ( .A(n50966), .B(n42615), .Y(n26665) );
  XNOR2X1 U45927 ( .A(n51160), .B(n41281), .Y(n24781) );
  XNOR2X1 U45928 ( .A(n50521), .B(n41380), .Y(n24867) );
  XNOR2X1 U45929 ( .A(n51163), .B(n42625), .Y(n24863) );
  XNOR2X1 U45930 ( .A(n51159), .B(n41283), .Y(n24751) );
  XNOR2X1 U45931 ( .A(n50514), .B(n42725), .Y(n28153) );
  XNOR2X1 U45932 ( .A(n50513), .B(n41380), .Y(n28145) );
  XNOR2X1 U45933 ( .A(n51155), .B(n42625), .Y(n28141) );
  XNOR2X1 U45934 ( .A(n50734), .B(n42505), .Y(n24854) );
  XNOR2X1 U45935 ( .A(n51157), .B(n41281), .Y(n24811) );
  XNOR2X1 U45936 ( .A(n50496), .B(n41380), .Y(n31544) );
  XNOR2X1 U45937 ( .A(n51138), .B(n42625), .Y(n31540) );
  XNOR2X1 U45938 ( .A(n51168), .B(n41281), .Y(n24991) );
  XNOR2X1 U45939 ( .A(n50525), .B(n36905), .Y(n24987) );
  XNOR2X1 U45940 ( .A(n51167), .B(n42627), .Y(n24983) );
  XNOR2X1 U45941 ( .A(n50724), .B(n42503), .Y(n28162) );
  XNOR2X1 U45942 ( .A(n51181), .B(n41281), .Y(n26674) );
  XNOR2X1 U45943 ( .A(n50538), .B(n36905), .Y(n26670) );
  XNOR2X1 U45944 ( .A(n51180), .B(n42629), .Y(n26666) );
  XOR2X1 U45945 ( .A(n42170), .B(n36881), .Y(n28155) );
  XOR2X1 U45946 ( .A(n42171), .B(n41286), .Y(n28147) );
  XOR2X1 U45947 ( .A(n41912), .B(n42600), .Y(n28143) );
  XOR2X1 U45948 ( .A(n42161), .B(n36879), .Y(n25177) );
  XOR2X1 U45949 ( .A(n41902), .B(n36899), .Y(n25173) );
  XOR2X1 U45950 ( .A(n42162), .B(n42656), .Y(n25169) );
  XOR2X1 U45951 ( .A(n41903), .B(n42611), .Y(n25165) );
  XOR2X1 U45952 ( .A(n41928), .B(n36900), .Y(n31550) );
  XOR2X1 U45953 ( .A(n42187), .B(n36879), .Y(n31554) );
  XOR2X1 U45954 ( .A(n42188), .B(n42665), .Y(n31546) );
  XOR2X1 U45955 ( .A(n41929), .B(n42608), .Y(n31542) );
  XOR2X1 U45956 ( .A(n41932), .B(n36899), .Y(n31400) );
  XOR2X1 U45957 ( .A(n42191), .B(n36887), .Y(n31404) );
  XOR2X1 U45958 ( .A(n41914), .B(n41312), .Y(n23216) );
  XOR2X1 U45959 ( .A(n41879), .B(n41314), .Y(n22349) );
  XOR2X1 U45960 ( .A(n41889), .B(n41314), .Y(n24129) );
  XOR2X1 U45961 ( .A(n41913), .B(n42522), .Y(n28133) );
  XOR2X1 U45962 ( .A(n41888), .B(n42522), .Y(n26658) );
  XNOR2X1 U45963 ( .A(n50546), .B(n36776), .Y(n22351) );
  XNOR2X1 U45964 ( .A(n51411), .B(n36740), .Y(n19548) );
  XNOR2X1 U45965 ( .A(n51391), .B(n36743), .Y(n19801) );
  XNOR2X1 U45966 ( .A(n51395), .B(n36743), .Y(n19731) );
  XNOR2X1 U45967 ( .A(n50528), .B(n36779), .Y(n235530) );
  XNOR2X1 U45968 ( .A(n50532), .B(n36767), .Y(n19741) );
  XNOR2X1 U45969 ( .A(n51391), .B(n41303), .Y(n24131) );
  XNOR2X1 U45970 ( .A(n51375), .B(n41303), .Y(n23595) );
  XNOR2X1 U45971 ( .A(n50535), .B(n36764), .Y(n19811) );
  XNOR2X1 U45972 ( .A(n51366), .B(n41303), .Y(n23218) );
  XNOR2X1 U45973 ( .A(n50529), .B(n36777), .Y(n24162) );
  XNOR2X1 U45974 ( .A(n50528), .B(n36768), .Y(n21011) );
  XNOR2X1 U45975 ( .A(n51185), .B(n42552), .Y(n26746) );
  XNOR2X1 U45976 ( .A(n50520), .B(n42579), .Y(n24857) );
  XNOR2X1 U45977 ( .A(n50512), .B(n42583), .Y(n28135) );
  XNOR2X1 U45978 ( .A(n50506), .B(n42582), .Y(n28555) );
  CLKINVX1 U45979 ( .A(net210259), .Y(net171537) );
  XOR2X1 U45980 ( .A(n42173), .B(n36809), .Y(n23217) );
  XOR2X1 U45981 ( .A(n41898), .B(n36897), .Y(n25113) );
  XOR2X1 U45982 ( .A(n41899), .B(n36710), .Y(n25105) );
  XOR2X1 U45983 ( .A(n42151), .B(n36817), .Y(n24100) );
  XOR2X1 U45984 ( .A(n42148), .B(n42490), .Y(n19800) );
  XOR2X1 U45985 ( .A(n42148), .B(n36810), .Y(n24130) );
  XOR2X1 U45986 ( .A(n42149), .B(n42490), .Y(n19810) );
  XOR2X1 U45987 ( .A(n42128), .B(n42480), .Y(n19547) );
  XOR2X1 U45988 ( .A(n42172), .B(n41322), .Y(n28134) );
  XOR2X1 U45989 ( .A(n42147), .B(n41321), .Y(n26659) );
  NOR4X1 U45990 ( .A(n19616), .B(n19615), .C(n19614), .D(n19613), .Y(n47224)
         );
  XNOR2X1 U45991 ( .A(n50749), .B(n42466), .Y(n19808) );
  XNOR2X1 U45992 ( .A(n51177), .B(n36717), .Y(n19807) );
  NOR4X1 U45993 ( .A(n21009), .B(n21008), .C(n21007), .D(n21006), .Y(n46956)
         );
  NOR4X1 U45994 ( .A(n25204), .B(n25205), .C(n25206), .D(n25207), .Y(n44423)
         );
  NOR4X1 U45995 ( .A(n24874), .B(n24875), .C(n24876), .D(n24877), .Y(n44526)
         );
  XNOR2X1 U45996 ( .A(n50318), .B(n42708), .Y(n24874) );
  XNOR2X1 U45997 ( .A(n50522), .B(n41287), .Y(n24875) );
  XNOR2X1 U45998 ( .A(n51377), .B(n42695), .Y(n24876) );
  NOR4X1 U45999 ( .A(n24964), .B(n24965), .C(n24966), .D(n24967), .Y(n44499)
         );
  XNOR2X1 U46000 ( .A(n50315), .B(n42707), .Y(n24964) );
  XNOR2X1 U46001 ( .A(n50519), .B(n42722), .Y(n24965) );
  XNOR2X1 U46002 ( .A(n51374), .B(n42695), .Y(n24966) );
  NOR4X1 U46003 ( .A(n24754), .B(n24755), .C(n24756), .D(n24757), .Y(n44561)
         );
  XNOR2X1 U46004 ( .A(n50313), .B(n42708), .Y(n24754) );
  XNOR2X1 U46005 ( .A(n50517), .B(n41287), .Y(n24755) );
  XNOR2X1 U46006 ( .A(n51372), .B(n42697), .Y(n24756) );
  NOR4X1 U46007 ( .A(n25174), .B(n25175), .C(n25176), .D(n25177), .Y(n44432)
         );
  XNOR2X1 U46008 ( .A(n50319), .B(n42707), .Y(n25174) );
  XNOR2X1 U46009 ( .A(n50523), .B(n36709), .Y(n25175) );
  XNOR2X1 U46010 ( .A(n51378), .B(n42691), .Y(n25176) );
  NOR4X1 U46011 ( .A(n24904), .B(n24905), .C(n24906), .D(n24907), .Y(n44517)
         );
  XNOR2X1 U46012 ( .A(n50317), .B(n42707), .Y(n24904) );
  XNOR2X1 U46013 ( .A(n50521), .B(n42722), .Y(n24905) );
  XNOR2X1 U46014 ( .A(n51376), .B(n42695), .Y(n24906) );
  NOR4X1 U46015 ( .A(n24994), .B(n24995), .C(n24996), .D(n24997), .Y(n44490)
         );
  XNOR2X1 U46016 ( .A(n50322), .B(n42707), .Y(n24994) );
  XNOR2X1 U46017 ( .A(n50526), .B(n36709), .Y(n24995) );
  XNOR2X1 U46018 ( .A(n51381), .B(n42695), .Y(n24996) );
  NOR4X1 U46019 ( .A(n25024), .B(n25025), .C(n25026), .D(n25027), .Y(n44485)
         );
  XNOR2X1 U46020 ( .A(n50321), .B(n42707), .Y(n25024) );
  XNOR2X1 U46021 ( .A(n50525), .B(n36709), .Y(n25025) );
  XNOR2X1 U46022 ( .A(n51380), .B(n36871), .Y(n25026) );
  NOR4X1 U46023 ( .A(n24836), .B(n24837), .C(n24838), .D(n24839), .Y(n44534)
         );
  NOR4X1 U46024 ( .A(n25084), .B(n25085), .C(n25086), .D(n25087), .Y(n44467)
         );
  XNOR2X1 U46025 ( .A(n50326), .B(n42707), .Y(n25084) );
  XNOR2X1 U46026 ( .A(n50530), .B(n42720), .Y(n25085) );
  XNOR2X1 U46027 ( .A(n51385), .B(n42695), .Y(n25086) );
  NOR4X1 U46028 ( .A(n27068), .B(n27069), .C(n27070), .D(n27071), .Y(n44234)
         );
  XNOR2X1 U46029 ( .A(n50327), .B(n42710), .Y(n27068) );
  XNOR2X1 U46030 ( .A(n50531), .B(n42723), .Y(n27069) );
  XNOR2X1 U46031 ( .A(n51386), .B(n42697), .Y(n27070) );
  NOR4X1 U46032 ( .A(n25054), .B(n25055), .C(n25056), .D(n25057), .Y(n44476)
         );
  XNOR2X1 U46033 ( .A(n51156), .B(n41281), .Y(n28149) );
  NOR4X1 U46034 ( .A(n28118), .B(n28119), .C(n28120), .D(n28121), .Y(n43806)
         );
  NOR4X1 U46035 ( .A(n28238), .B(n28239), .C(n28240), .D(n28241), .Y(n43770)
         );
  XNOR2X1 U46036 ( .A(n50938), .B(n40039), .Y(n28238) );
  XNOR2X1 U46037 ( .A(n51152), .B(n41281), .Y(n28239) );
  XNOR2X1 U46038 ( .A(n50724), .B(net219468), .Y(n28240) );
  NOR4X1 U46039 ( .A(n28418), .B(n28419), .C(n28420), .D(n28421), .Y(n43724)
         );
  NOR4X1 U46040 ( .A(n28208), .B(n28209), .C(n28210), .D(n28211), .Y(n43779)
         );
  XNOR2X1 U46041 ( .A(n50925), .B(net219310), .Y(n31547) );
  XNOR2X1 U46042 ( .A(n51139), .B(n41283), .Y(n31548) );
  XNOR2X1 U46043 ( .A(n50711), .B(net219450), .Y(n31549) );
  NOR4X1 U46044 ( .A(n28268), .B(n28269), .C(n28270), .D(n28271), .Y(n43761)
         );
  NOR4X1 U46045 ( .A(n31577), .B(n31578), .C(n31579), .D(n31580), .Y(n43211)
         );
  NOR4X1 U46046 ( .A(n31397), .B(n31398), .C(n31399), .D(n31400), .Y(n43265)
         );
  XNOR2X1 U46047 ( .A(n50921), .B(n40039), .Y(n31397) );
  XNOR2X1 U46048 ( .A(n51135), .B(n41282), .Y(n31398) );
  XNOR2X1 U46049 ( .A(n50707), .B(net219450), .Y(n31399) );
  XNOR2X1 U46050 ( .A(n50919), .B(n36870), .Y(n31307) );
  XNOR2X1 U46051 ( .A(n51133), .B(n41281), .Y(n31308) );
  XNOR2X1 U46052 ( .A(n50705), .B(net219434), .Y(n31309) );
  NOR4X1 U46053 ( .A(n31607), .B(n31608), .C(n31609), .D(n31610), .Y(n43202)
         );
  XNOR2X1 U46054 ( .A(n50923), .B(n40039), .Y(n31607) );
  XNOR2X1 U46055 ( .A(n51137), .B(n41281), .Y(n31608) );
  XNOR2X1 U46056 ( .A(n50709), .B(net219450), .Y(n31609) );
  NOR4X1 U46057 ( .A(n28328), .B(n28329), .C(n28330), .D(n28331), .Y(n43747)
         );
  NOR4X1 U46058 ( .A(n28448), .B(n28449), .C(n28450), .D(n28451), .Y(n43715)
         );
  XNOR2X1 U46059 ( .A(n50929), .B(net219310), .Y(n28448) );
  XNOR2X1 U46060 ( .A(n51143), .B(n41282), .Y(n28449) );
  XNOR2X1 U46061 ( .A(n50715), .B(net219468), .Y(n28450) );
  NOR4X1 U46062 ( .A(n28388), .B(n28389), .C(n28390), .D(n28391), .Y(n43733)
         );
  XNOR2X1 U46063 ( .A(n50927), .B(n40039), .Y(n28388) );
  XNOR2X1 U46064 ( .A(n51141), .B(n41282), .Y(n28389) );
  XNOR2X1 U46065 ( .A(n50713), .B(net219468), .Y(n28390) );
  NOR4X1 U46066 ( .A(n31637), .B(n31638), .C(n31639), .D(n31640), .Y(n43193)
         );
  XNOR2X1 U46067 ( .A(n50924), .B(n40039), .Y(n31637) );
  XNOR2X1 U46068 ( .A(n51138), .B(n41281), .Y(n31638) );
  XNOR2X1 U46069 ( .A(n50710), .B(net219450), .Y(n31639) );
  NOR4X1 U46070 ( .A(n31277), .B(n31278), .C(n31279), .D(n31280), .Y(n43300)
         );
  XNOR2X1 U46071 ( .A(n50914), .B(net219310), .Y(n31277) );
  XNOR2X1 U46072 ( .A(n51128), .B(n41281), .Y(n31278) );
  XNOR2X1 U46073 ( .A(n50700), .B(net219460), .Y(n31279) );
  NOR4X1 U46074 ( .A(n28178), .B(n28179), .C(n28180), .D(n28181), .Y(n43788)
         );
  XNOR2X1 U46075 ( .A(n50940), .B(net219314), .Y(n28178) );
  XNOR2X1 U46076 ( .A(n51154), .B(n41281), .Y(n28179) );
  XNOR2X1 U46077 ( .A(n50726), .B(net219468), .Y(n28180) );
  NOR4X1 U46078 ( .A(n28538), .B(n28539), .C(n28540), .D(n28541), .Y(n43688)
         );
  NOR4X1 U46079 ( .A(n28508), .B(n28509), .C(n28510), .D(n28511), .Y(n43697)
         );
  NOR4X1 U46080 ( .A(n28358), .B(n28359), .C(n28360), .D(n28361), .Y(n43742)
         );
  XNOR2X1 U46081 ( .A(n50933), .B(n40039), .Y(n28358) );
  XNOR2X1 U46082 ( .A(n51147), .B(n41281), .Y(n28359) );
  XNOR2X1 U46083 ( .A(n50719), .B(net219468), .Y(n28360) );
  NOR4X1 U46084 ( .A(n28298), .B(n28299), .C(n28300), .D(n28301), .Y(n43752)
         );
  XNOR2X1 U46085 ( .A(n50931), .B(net219336), .Y(n28298) );
  XNOR2X1 U46086 ( .A(n51145), .B(n41282), .Y(n28299) );
  XNOR2X1 U46087 ( .A(n50717), .B(net219468), .Y(n28300) );
  NOR4X1 U46088 ( .A(n28478), .B(n28479), .C(n28480), .D(n28481), .Y(n43706)
         );
  NOR4X1 U46089 ( .A(n31367), .B(n31368), .C(n31369), .D(n31370), .Y(n43273)
         );
  NOR4X1 U46090 ( .A(n31187), .B(n31188), .C(n31189), .D(n31190), .Y(n43327)
         );
  XNOR2X1 U46091 ( .A(n50912), .B(net219310), .Y(n31187) );
  XNOR2X1 U46092 ( .A(n51126), .B(n41283), .Y(n31188) );
  XNOR2X1 U46093 ( .A(n50698), .B(net219434), .Y(n31189) );
  NOR4X1 U46094 ( .A(n28568), .B(n28569), .C(n28570), .D(n28571), .Y(n43681)
         );
  XNOR2X1 U46095 ( .A(n50936), .B(n40039), .Y(n28568) );
  XNOR2X1 U46096 ( .A(n51150), .B(n41281), .Y(n28569) );
  XNOR2X1 U46097 ( .A(n50722), .B(net219468), .Y(n28570) );
  NOR4X1 U46098 ( .A(n24972), .B(n24973), .C(n24974), .D(n24977), .Y(n44497)
         );
  XNOR2X1 U46099 ( .A(n50757), .B(n42506), .Y(n26747) );
  CLKINVX1 U46100 ( .A(n10726), .Y(net151726) );
  CLKINVX1 U46101 ( .A(n10863), .Y(net209250) );
  CLKINVX1 U46102 ( .A(n10725), .Y(net151728) );
  CLKINVX1 U46103 ( .A(n45727), .Y(n49501) );
  OAI21XL U46104 ( .A0(net171486), .A1(n48422), .B0(n12329), .Y(n48424) );
  AOI21X1 U46105 ( .A0(n48421), .A1(n12384), .B0(net171489), .Y(n48422) );
  OAI21XL U46106 ( .A0(n11201), .A1(net209362), .B0(n12333), .Y(n48421) );
  CLKINVX1 U46107 ( .A(n11200), .Y(net209362) );
  CLKINVX1 U46108 ( .A(n48166), .Y(n48184) );
  CLKINVX1 U46109 ( .A(net209303), .Y(net209280) );
  CLKINVX1 U46110 ( .A(n12387), .Y(net171440) );
  CLKINVX1 U46111 ( .A(n11349), .Y(net210075) );
  CLKINVX1 U46112 ( .A(n10555), .Y(net171257) );
  CLKINVX1 U46113 ( .A(n12702), .Y(n48227) );
  OAI21XL U46114 ( .A0(net151726), .A1(n48054), .B0(n10724), .Y(n48055) );
  OAI21XL U46115 ( .A0(net171546), .A1(net210132), .B0(n12970), .Y(n48053) );
  OAI2BB1X1 U46116 ( .A0N(n48222), .A1N(n12150), .B0(net209817), .Y(n48224) );
  OAI2BB1X1 U46117 ( .A0N(n48127), .A1N(n12146), .B0(n12731), .Y(n48129) );
  CLKINVX1 U46118 ( .A(n48461), .Y(n48466) );
  CLKINVX1 U46119 ( .A(n12079), .Y(net209956) );
  CLKINVX1 U46120 ( .A(n11074), .Y(net209210) );
  CLKINVX1 U46121 ( .A(n10872), .Y(net209258) );
  OAI21XL U46122 ( .A0(net209289), .A1(net209290), .B0(net209291), .Y(n48460)
         );
  AOI21X1 U46123 ( .A0(n48244), .A1(n12015), .B0(net209787), .Y(n48245) );
  CLKINVX1 U46124 ( .A(n12157), .Y(net209787) );
  AOI21X1 U46125 ( .A0(n48097), .A1(n11512), .B0(n37240), .Y(n48098) );
  OAI21XL U46126 ( .A0(net210075), .A1(n48096), .B0(n11511), .Y(n48097) );
  AOI21X1 U46127 ( .A0(n48095), .A1(n11351), .B0(net210078), .Y(n48096) );
  CLKINVX1 U46128 ( .A(n11348), .Y(net210078) );
  CLKINVX1 U46129 ( .A(n12016), .Y(net209791) );
  OAI21XL U46130 ( .A0(net171210), .A1(n48241), .B0(n12692), .Y(n48242) );
  AOI211X1 U46131 ( .A0(n47978), .A1(n47998), .B0(n47977), .C0(n47976), .Y(
        n48017) );
  OAI21XL U46132 ( .A0(n48004), .A1(n48003), .B0(n48002), .Y(n48016) );
  AOI21X1 U46133 ( .A0(n47958), .A1(n11369), .B0(n47957), .Y(n47959) );
  CLKINVX1 U46134 ( .A(n11372), .Y(net210251) );
  OAI21XL U46135 ( .A0(net151672), .A1(n47971), .B0(n11441), .Y(n47973) );
  CLKINVX1 U46136 ( .A(n48173), .Y(n48174) );
  AOI21X1 U46137 ( .A0(n47965), .A1(n11423), .B0(net210242), .Y(n47966) );
  CLKINVX1 U46138 ( .A(n11416), .Y(net210242) );
  OAI21XL U46139 ( .A0(n12951), .A1(n47964), .B0(n11422), .Y(n47965) );
  AOI21X1 U46140 ( .A0(n47963), .A1(n12954), .B0(n37205), .Y(n47964) );
  CLKINVX1 U46141 ( .A(n48179), .Y(n48180) );
  AOI21X1 U46142 ( .A0(n48219), .A1(n12723), .B0(net171257), .Y(n48220) );
  OAI21XL U46143 ( .A0(n12062), .A1(net171252), .B0(n12726), .Y(n48219) );
  OAI21XL U46144 ( .A0(net209250), .A1(n48484), .B0(n40397), .Y(n48489) );
  CLKINVX1 U46145 ( .A(n11132), .Y(net209254) );
  AOI21X1 U46146 ( .A0(n47955), .A1(n11377), .B0(net210254), .Y(n47956) );
  CLKINVX1 U46147 ( .A(n11371), .Y(net210254) );
  OAI21XL U46148 ( .A0(net210255), .A1(n47954), .B0(n11376), .Y(n47955) );
  CLKINVX1 U46149 ( .A(n11379), .Y(net210255) );
  OAI21XL U46150 ( .A0(net209367), .A1(n48416), .B0(n11209), .Y(n48417) );
  OAI21XL U46151 ( .A0(net209280), .A1(n48463), .B0(n48462), .Y(n48472) );
  NOR2X1 U46152 ( .A(n48466), .B(net209283), .Y(n48462) );
  NAND2X1 U46153 ( .A(n48018), .B(n48030), .Y(n48023) );
  AOI21X1 U46154 ( .A0(n48502), .A1(n11204), .B0(net171417), .Y(n48503) );
  CLKINVX1 U46155 ( .A(n10852), .Y(net209228) );
  NOR2BX1 U46156 ( .AN(n10727), .B(n36948), .Y(n48047) );
  AOI21X1 U46157 ( .A0(n48119), .A1(n12706), .B0(n48227), .Y(n48120) );
  CLKINVX1 U46158 ( .A(n11358), .Y(net210081) );
  NOR2X1 U46159 ( .A(n48230), .B(n48229), .Y(n48231) );
  AOI21X1 U46160 ( .A0(n47953), .A1(n12929), .B0(net210258), .Y(n47954) );
  CLKINVX1 U46161 ( .A(n11378), .Y(net210258) );
  NOR3X1 U46162 ( .A(n48080), .B(n48079), .C(n48078), .Y(n48081) );
  NOR3X1 U46163 ( .A(n48060), .B(n48059), .C(n48058), .Y(n48061) );
  NOR2X1 U46164 ( .A(n48042), .B(n48041), .Y(n48043) );
  CLKINVX1 U46165 ( .A(n48007), .Y(n48008) );
  CLKINVX1 U46166 ( .A(n48006), .Y(n48010) );
  NOR2X1 U46167 ( .A(n47991), .B(net210221), .Y(n47994) );
  NOR3X1 U46168 ( .A(n48470), .B(n48469), .C(n48468), .Y(n48471) );
  NOR3X1 U46169 ( .A(n48506), .B(n48505), .C(n48504), .Y(n48507) );
  NOR3X1 U46170 ( .A(n48487), .B(n48486), .C(n48485), .Y(n48488) );
  NAND2X1 U46171 ( .A(n12322), .B(n12385), .Y(n48485) );
  NAND2X1 U46172 ( .A(n47998), .B(n47997), .Y(n47999) );
  NAND4BBXL U46173 ( .AN(n48049), .BN(n48048), .C(n48047), .D(n48046), .Y(
        n48050) );
  NAND2X1 U46174 ( .A(n10726), .B(n12967), .Y(n48049) );
  NAND2X1 U46175 ( .A(net210142), .B(n10730), .Y(n48048) );
  NAND2X1 U46176 ( .A(n10732), .B(net210140), .Y(n48046) );
  NAND4BX1 U46177 ( .AN(n48089), .B(n48088), .C(n48087), .D(n48086), .Y(n48090) );
  NOR2X1 U46178 ( .A(net210075), .B(n48085), .Y(n48087) );
  NOR2BX1 U46179 ( .AN(n13018), .B(net210089), .Y(n48086) );
  NAND3X1 U46180 ( .A(n48122), .B(n40386), .C(n12153), .Y(n48123) );
  NAND4X1 U46181 ( .A(n48069), .B(n10706), .C(n48068), .D(n48067), .Y(n48070)
         );
  NOR2X1 U46182 ( .A(n48066), .B(n48065), .Y(n48067) );
  OAI21XL U46183 ( .A0(n48064), .A1(n48063), .B0(n48062), .Y(n48069) );
  NOR2X1 U46184 ( .A(n48213), .B(n48212), .Y(n48214) );
  NOR2X1 U46185 ( .A(n48190), .B(n48189), .Y(n48191) );
  NOR2X1 U46186 ( .A(n48195), .B(n48194), .Y(n48197) );
  NOR2X1 U46187 ( .A(n48235), .B(n48234), .Y(n48236) );
  NAND2X1 U46188 ( .A(n12156), .B(n12015), .Y(n48234) );
  CLKINVX1 U46189 ( .A(n48171), .Y(n48178) );
  NOR3X1 U46190 ( .A(n48208), .B(n48207), .C(n48206), .Y(n48209) );
  CLKINVX1 U46191 ( .A(n12708), .Y(net209969) );
  CLKINVX1 U46192 ( .A(n11351), .Y(net210089) );
  NAND2X1 U46193 ( .A(n48205), .B(n10567), .Y(n48210) );
  AOI21X1 U46194 ( .A0(n48203), .A1(n12744), .B0(net209840), .Y(n48204) );
  CLKINVX1 U46195 ( .A(n11083), .Y(n48419) );
  NAND2BX1 U46196 ( .AN(n12342), .B(net209267), .Y(n48474) );
  NAND2X1 U46197 ( .A(n11377), .B(n11372), .Y(n48079) );
  NAND3X1 U46198 ( .A(n11365), .B(n11509), .C(n11369), .Y(n48078) );
  CLKINVX1 U46199 ( .A(net210234), .Y(net210233) );
  CLKINVX1 U46200 ( .A(n10733), .Y(net210140) );
  NOR2X1 U46201 ( .A(n48162), .B(n48161), .Y(n48163) );
  NAND2X1 U46202 ( .A(n11414), .B(n11417), .Y(n48058) );
  AND2X2 U46203 ( .A(n48011), .B(n48020), .Y(n48012) );
  CLKINVX1 U46204 ( .A(n48005), .Y(n48014) );
  CLKINVX1 U46205 ( .A(n12292), .Y(net171449) );
  AOI21X1 U46206 ( .A0(n10689), .A1(n50102), .B0(n48084), .Y(n48088) );
  CLKINVX1 U46207 ( .A(n11360), .Y(n48084) );
  NAND3X1 U46208 ( .A(n48522), .B(n11058), .C(n11065), .Y(n48513) );
  NAND2X1 U46209 ( .A(net210091), .B(n11512), .Y(n48085) );
  XNOR2X1 U46210 ( .A(n50953), .B(n42539), .Y(n25092) );
  XNOR2X1 U46211 ( .A(n51167), .B(n42551), .Y(n25093) );
  XNOR2X1 U46212 ( .A(n50739), .B(n36730), .Y(n25094) );
  XNOR2X1 U46213 ( .A(n50525), .B(n42580), .Y(n25097) );
  CLKINVX1 U46214 ( .A(n11114), .Y(net209234) );
  NOR2X1 U46215 ( .A(n25138), .B(n25139), .Y(n44445) );
  XNOR2X1 U46216 ( .A(n51382), .B(n42702), .Y(n25116) );
  NOR2X1 U46217 ( .A(n25108), .B(n25109), .Y(n44453) );
  XNOR2X1 U46218 ( .A(n51381), .B(n42638), .Y(n25108) );
  XOR2X1 U46219 ( .A(n42158), .B(n42656), .Y(n25109) );
  NOR2X1 U46220 ( .A(n25146), .B(n25147), .Y(n44441) );
  CLKINVX1 U46221 ( .A(n48019), .Y(n48021) );
  OAI2BB1X1 U46222 ( .A0N(n48031), .A1N(n48030), .B0(n48029), .Y(n48035) );
  CLKINVX1 U46223 ( .A(n48028), .Y(n48031) );
  OAI2BB1X1 U46224 ( .A0N(n13015), .A1N(net171554), .B0(n12957), .Y(n47963) );
  AND2X2 U46225 ( .A(n12702), .B(n12706), .Y(n12036) );
  CLKINVX1 U46226 ( .A(n47974), .Y(n47978) );
  AND2X2 U46227 ( .A(n11204), .B(n12386), .Y(n48492) );
  NAND2X1 U46228 ( .A(n41786), .B(n41787), .Y(n44496) );
  XNOR2X1 U46229 ( .A(n42160), .B(n36873), .Y(n41786) );
  XNOR2X1 U46230 ( .A(n41901), .B(n42522), .Y(n41787) );
  XNOR2X1 U46231 ( .A(n50947), .B(n36799), .Y(n21067) );
  XNOR2X1 U46232 ( .A(n50948), .B(n36796), .Y(n21077) );
  XNOR2X1 U46233 ( .A(n50946), .B(n36799), .Y(n21057) );
  XNOR2X1 U46234 ( .A(n50945), .B(n36793), .Y(n21047) );
  XNOR2X1 U46235 ( .A(n50924), .B(n36792), .Y(n21601) );
  XNOR2X1 U46236 ( .A(n50922), .B(n41294), .Y(n22943) );
  XNOR2X1 U46237 ( .A(n50925), .B(n41294), .Y(n23173) );
  XNOR2X1 U46238 ( .A(n50920), .B(n36796), .Y(n21501) );
  XNOR2X1 U46239 ( .A(n50944), .B(n41291), .Y(n23468) );
  XNOR2X1 U46240 ( .A(n50944), .B(n36798), .Y(n21097) );
  XNOR2X1 U46241 ( .A(n50924), .B(n41297), .Y(n22963) );
  XNOR2X1 U46242 ( .A(n50927), .B(n36791), .Y(n19998) );
  XNOR2X1 U46243 ( .A(n50928), .B(n36792), .Y(n20008) );
  XNOR2X1 U46244 ( .A(n50923), .B(n42538), .Y(n31529) );
  XNOR2X1 U46245 ( .A(n50922), .B(n42538), .Y(n31619) );
  XNOR2X1 U46246 ( .A(n50919), .B(n42537), .Y(n31379) );
  XNOR2X1 U46247 ( .A(n50905), .B(n42544), .Y(n31830) );
  XNOR2X1 U46248 ( .A(n51348), .B(n42702), .Y(n31403) );
  XNOR2X1 U46249 ( .A(n51346), .B(n42702), .Y(n31313) );
  XNOR2X1 U46250 ( .A(n51142), .B(n41327), .Y(n23184) );
  XNOR2X1 U46251 ( .A(n51161), .B(n36716), .Y(n21068) );
  XNOR2X1 U46252 ( .A(n51162), .B(n36714), .Y(n21078) );
  XNOR2X1 U46253 ( .A(n51160), .B(n36721), .Y(n21058) );
  XNOR2X1 U46254 ( .A(n51159), .B(n36720), .Y(n21048) );
  XNOR2X1 U46255 ( .A(n51138), .B(n36722), .Y(n21602) );
  XNOR2X1 U46256 ( .A(n51136), .B(n41330), .Y(n22944) );
  XNOR2X1 U46257 ( .A(n51139), .B(n41331), .Y(n23174) );
  XNOR2X1 U46258 ( .A(n51134), .B(n36715), .Y(n21502) );
  XNOR2X1 U46259 ( .A(n51158), .B(n41331), .Y(n23469) );
  XNOR2X1 U46260 ( .A(n51158), .B(n36717), .Y(n21098) );
  XNOR2X1 U46261 ( .A(n51138), .B(n41331), .Y(n22964) );
  XNOR2X1 U46262 ( .A(n51141), .B(n36721), .Y(n19999) );
  XNOR2X1 U46263 ( .A(n51142), .B(n36722), .Y(n20009) );
  XNOR2X1 U46264 ( .A(n51345), .B(n42637), .Y(n31305) );
  XNOR2X1 U46265 ( .A(n50704), .B(n42588), .Y(n31301) );
  XNOR2X1 U46266 ( .A(n51137), .B(n42550), .Y(n31530) );
  XNOR2X1 U46267 ( .A(n51136), .B(n42550), .Y(n31620) );
  XNOR2X1 U46268 ( .A(n51131), .B(n42552), .Y(n31290) );
  XNOR2X1 U46269 ( .A(n51122), .B(n42552), .Y(n31771) );
  XNOR2X1 U46270 ( .A(n51336), .B(n42638), .Y(n31786) );
  XNOR2X1 U46271 ( .A(n50695), .B(n42589), .Y(n31782) );
  XNOR2X1 U46272 ( .A(n50492), .B(n42720), .Y(n31312) );
  XNOR2X1 U46273 ( .A(n50484), .B(n36709), .Y(n31793) );
  XNOR2X1 U46274 ( .A(n50733), .B(n42467), .Y(n21069) );
  XNOR2X1 U46275 ( .A(n50734), .B(n42460), .Y(n21079) );
  XNOR2X1 U46276 ( .A(n50732), .B(n42460), .Y(n21059) );
  XNOR2X1 U46277 ( .A(n50731), .B(n42459), .Y(n21049) );
  XNOR2X1 U46278 ( .A(n50710), .B(n42466), .Y(n21603) );
  XNOR2X1 U46279 ( .A(n50708), .B(n36853), .Y(n22945) );
  XNOR2X1 U46280 ( .A(n50711), .B(n36852), .Y(n23175) );
  XNOR2X1 U46281 ( .A(n50706), .B(n42459), .Y(n21503) );
  XNOR2X1 U46282 ( .A(n50730), .B(n36856), .Y(n23470) );
  XNOR2X1 U46283 ( .A(n50730), .B(n42460), .Y(n21099) );
  XNOR2X1 U46284 ( .A(n50710), .B(n36850), .Y(n22965) );
  XNOR2X1 U46285 ( .A(n50713), .B(n42467), .Y(n20000) );
  XNOR2X1 U46286 ( .A(n50714), .B(n42467), .Y(n20010) );
  XNOR2X1 U46287 ( .A(n50287), .B(n42712), .Y(n31311) );
  XNOR2X1 U46288 ( .A(n50286), .B(n42669), .Y(n31303) );
  XNOR2X1 U46289 ( .A(n50918), .B(n42617), .Y(n31299) );
  XNOR2X1 U46290 ( .A(n50292), .B(n42708), .Y(n31641) );
  XNOR2X1 U46291 ( .A(n50278), .B(n42706), .Y(n31792) );
  XNOR2X1 U46292 ( .A(n50277), .B(n42671), .Y(n31784) );
  XNOR2X1 U46293 ( .A(n50909), .B(n42614), .Y(n31780) );
  XNOR2X1 U46294 ( .A(n50491), .B(n41380), .Y(n31304) );
  XNOR2X1 U46295 ( .A(n51132), .B(n34447), .Y(n31300) );
  XNOR2X1 U46296 ( .A(n50709), .B(n42499), .Y(n31531) );
  XNOR2X1 U46297 ( .A(n50708), .B(n42499), .Y(n31621) );
  XNOR2X1 U46298 ( .A(n50705), .B(n42505), .Y(n31381) );
  XNOR2X1 U46299 ( .A(n50483), .B(n36905), .Y(n31785) );
  XNOR2X1 U46300 ( .A(n51123), .B(n42624), .Y(n31781) );
  XNOR2X1 U46301 ( .A(n50692), .B(n42508), .Y(n31862) );
  XOR2X1 U46302 ( .A(n42192), .B(n42656), .Y(n31396) );
  XOR2X1 U46303 ( .A(n41933), .B(n36819), .Y(n31392) );
  XOR2X1 U46304 ( .A(n42212), .B(n42652), .Y(n31125) );
  XOR2X1 U46305 ( .A(n41953), .B(n42606), .Y(n31121) );
  XOR2X1 U46306 ( .A(n41954), .B(n36899), .Y(n31069) );
  XOR2X1 U46307 ( .A(n42213), .B(n36889), .Y(n31073) );
  XOR2X1 U46308 ( .A(n41906), .B(n36754), .Y(n21070) );
  XOR2X1 U46309 ( .A(n41905), .B(n36756), .Y(n21080) );
  XOR2X1 U46310 ( .A(n41907), .B(n36753), .Y(n21060) );
  XOR2X1 U46311 ( .A(n41908), .B(n36756), .Y(n21050) );
  XOR2X1 U46312 ( .A(n41931), .B(n41316), .Y(n22946) );
  XOR2X1 U46313 ( .A(n41929), .B(n41313), .Y(n22966) );
  XOR2X1 U46314 ( .A(n41926), .B(n36757), .Y(n20001) );
  XOR2X1 U46315 ( .A(n41925), .B(n36761), .Y(n20011) );
  XOR2X1 U46316 ( .A(n41930), .B(n42519), .Y(n31532) );
  XOR2X1 U46317 ( .A(n41931), .B(n42519), .Y(n31622) );
  XOR2X1 U46318 ( .A(n41936), .B(n42518), .Y(n31292) );
  XOR2X1 U46319 ( .A(n41945), .B(n42520), .Y(n31773) );
  NOR4X1 U46320 ( .A(n22883), .B(n22884), .C(n22885), .D(n22886), .Y(n22882)
         );
  XNOR2X1 U46321 ( .A(n50500), .B(n36784), .Y(n23188) );
  XNOR2X1 U46322 ( .A(n51374), .B(n36741), .Y(n21072) );
  XNOR2X1 U46323 ( .A(n51375), .B(n36747), .Y(n21082) );
  XNOR2X1 U46324 ( .A(n50514), .B(n36764), .Y(n21122) );
  XNOR2X1 U46325 ( .A(n50496), .B(n36764), .Y(n21607) );
  XNOR2X1 U46326 ( .A(n51349), .B(n41301), .Y(n22948) );
  XNOR2X1 U46327 ( .A(n51342), .B(n36743), .Y(n21456) );
  XNOR2X1 U46328 ( .A(n51350), .B(n36742), .Y(n21596) );
  XNOR2X1 U46329 ( .A(n51371), .B(n36748), .Y(n21102) );
  XNOR2X1 U46330 ( .A(n50496), .B(n36780), .Y(n22968) );
  XNOR2X1 U46331 ( .A(n51343), .B(n36749), .Y(n21466) );
  XNOR2X1 U46332 ( .A(n50495), .B(n42578), .Y(n31534) );
  XNOR2X1 U46333 ( .A(n37251), .B(n42578), .Y(n31624) );
  XNOR2X1 U46334 ( .A(n50496), .B(n42578), .Y(n31564) );
  XNOR2X1 U46335 ( .A(n50492), .B(n42582), .Y(n31384) );
  XOR2X1 U46336 ( .A(n42165), .B(n42490), .Y(n21071) );
  XOR2X1 U46337 ( .A(n42164), .B(n42484), .Y(n21081) );
  XOR2X1 U46338 ( .A(n42166), .B(n42484), .Y(n21061) );
  XOR2X1 U46339 ( .A(n42167), .B(n42483), .Y(n21051) );
  XOR2X1 U46340 ( .A(n42190), .B(n36815), .Y(n22947) );
  XOR2X1 U46341 ( .A(n42187), .B(n36809), .Y(n23177) );
  XOR2X1 U46342 ( .A(n42167), .B(n36816), .Y(n23604) );
  XOR2X1 U46343 ( .A(n42188), .B(n36817), .Y(n22967) );
  XOR2X1 U46344 ( .A(n42185), .B(n42491), .Y(n20002) );
  XOR2X1 U46345 ( .A(n42189), .B(n41323), .Y(n31533) );
  XOR2X1 U46346 ( .A(n42190), .B(n41323), .Y(n31623) );
  XOR2X1 U46347 ( .A(n42195), .B(n36877), .Y(n31293) );
  XOR2X1 U46348 ( .A(n42204), .B(n41322), .Y(n31774) );
  NOR4X1 U46349 ( .A(n21464), .B(n21463), .C(n21462), .D(n21461), .Y(n46775)
         );
  NOR4X1 U46350 ( .A(n31337), .B(n31338), .C(n31339), .D(n31340), .Y(n43282)
         );
  NOR4X1 U46351 ( .A(n31517), .B(n31518), .C(n31519), .D(n31520), .Y(n43229)
         );
  NOR4X1 U46352 ( .A(n31217), .B(n31218), .C(n31219), .D(n31220), .Y(n43318)
         );
  XNOR2X1 U46353 ( .A(n50911), .B(net219310), .Y(n31217) );
  XNOR2X1 U46354 ( .A(n51125), .B(n41282), .Y(n31218) );
  XNOR2X1 U46355 ( .A(n50697), .B(net219460), .Y(n31219) );
  NOR4X1 U46356 ( .A(n31457), .B(n31458), .C(n31459), .D(n31460), .Y(n43247)
         );
  NOR4X1 U46357 ( .A(n31487), .B(n31488), .C(n31489), .D(n31490), .Y(n43238)
         );
  XNOR2X1 U46358 ( .A(n50915), .B(net219310), .Y(n31487) );
  XNOR2X1 U46359 ( .A(n51129), .B(n41283), .Y(n31488) );
  XNOR2X1 U46360 ( .A(n50701), .B(net219450), .Y(n31489) );
  NOR4X1 U46361 ( .A(n31698), .B(n31699), .C(n31700), .D(n31701), .Y(n43174)
         );
  NOR4X1 U46362 ( .A(n31788), .B(n31789), .C(n31790), .D(n31791), .Y(n43156)
         );
  XNOR2X1 U46363 ( .A(n50910), .B(net219308), .Y(n31788) );
  XNOR2X1 U46364 ( .A(n51124), .B(n41281), .Y(n31789) );
  XNOR2X1 U46365 ( .A(n50696), .B(net219434), .Y(n31790) );
  NOR4X1 U46366 ( .A(n31848), .B(n31849), .C(n31850), .D(n31851), .Y(n44583)
         );
  NOR4X1 U46367 ( .A(n31126), .B(n31127), .C(n31128), .D(n31129), .Y(n43341)
         );
  NOR4X1 U46368 ( .A(n31066), .B(n31067), .C(n31068), .D(n31069), .Y(n43358)
         );
  NOR4X1 U46369 ( .A(n31036), .B(n31037), .C(n31038), .D(n31039), .Y(n43366)
         );
  NOR4X1 U46370 ( .A(n31006), .B(n31007), .C(n31008), .D(n31009), .Y(n43375)
         );
  NOR4X1 U46371 ( .A(n31427), .B(n31428), .C(n31429), .D(n31430), .Y(n43256)
         );
  XNOR2X1 U46372 ( .A(n50917), .B(net219336), .Y(n31427) );
  XNOR2X1 U46373 ( .A(n51131), .B(n41281), .Y(n31428) );
  XNOR2X1 U46374 ( .A(n50703), .B(net219450), .Y(n31429) );
  NOR4X1 U46375 ( .A(n31247), .B(n31248), .C(n31249), .D(n31250), .Y(n43309)
         );
  XNOR2X1 U46376 ( .A(n50913), .B(n40039), .Y(n31247) );
  XNOR2X1 U46377 ( .A(n51127), .B(n41282), .Y(n31248) );
  XNOR2X1 U46378 ( .A(n50699), .B(net258207), .Y(n31249) );
  NOR4X1 U46379 ( .A(n31758), .B(n31759), .C(n31760), .D(n31761), .Y(n43165)
         );
  NOR4X1 U46380 ( .A(n31878), .B(n31879), .C(n31880), .D(n31881), .Y(n44637)
         );
  NOR4X1 U46381 ( .A(n31096), .B(n31097), .C(n31098), .D(n31099), .Y(n43349)
         );
  NOR4X1 U46382 ( .A(n31668), .B(n31669), .C(n31670), .D(n31671), .Y(net216758) );
  XNOR2X1 U46383 ( .A(n50905), .B(n36870), .Y(n31668) );
  XNOR2X1 U46384 ( .A(n51119), .B(n41282), .Y(n31669) );
  XNOR2X1 U46385 ( .A(n50691), .B(net219450), .Y(n31670) );
  NOR4X1 U46386 ( .A(n31818), .B(n31819), .C(n31820), .D(n31821), .Y(net214662) );
  NOR4X1 U46387 ( .A(n31728), .B(n31729), .C(n31730), .D(n31731), .Y(net216749) );
  NOR4X1 U46388 ( .A(n30976), .B(n30977), .C(n30978), .D(n30979), .Y(n43386)
         );
  NOR2X1 U46389 ( .A(n41735), .B(n12907), .Y(n10015) );
  CLKINVX1 U46390 ( .A(n11041), .Y(net209182) );
  CLKINVX1 U46391 ( .A(n12909), .Y(net151465) );
  AND2X2 U46392 ( .A(n11511), .B(n11512), .Y(n11342) );
  XNOR2X1 U46393 ( .A(n50907), .B(n36797), .Y(n21754) );
  XNOR2X1 U46394 ( .A(n50891), .B(n36797), .Y(n21410) );
  XNOR2X1 U46395 ( .A(n50890), .B(n41291), .Y(n22690) );
  XNOR2X1 U46396 ( .A(n50892), .B(n36789), .Y(n21420) );
  XNOR2X1 U46397 ( .A(n51121), .B(n36722), .Y(n21755) );
  XNOR2X1 U46398 ( .A(n51105), .B(n36718), .Y(n21411) );
  XNOR2X1 U46399 ( .A(n51104), .B(n36913), .Y(n22691) );
  XNOR2X1 U46400 ( .A(n51106), .B(n36716), .Y(n21421) );
  XNOR2X1 U46401 ( .A(n50693), .B(n42462), .Y(n21756) );
  XNOR2X1 U46402 ( .A(n50692), .B(n42462), .Y(n21696) );
  XNOR2X1 U46403 ( .A(n50677), .B(n42461), .Y(n21412) );
  XNOR2X1 U46404 ( .A(n50676), .B(n36858), .Y(n22692) );
  XNOR2X1 U46405 ( .A(n50678), .B(n42461), .Y(n21422) );
  XNOR2X1 U46406 ( .A(n50683), .B(n42499), .Y(n31050) );
  XOR2X1 U46407 ( .A(n42219), .B(n36887), .Y(n32156) );
  XOR2X1 U46408 ( .A(n42220), .B(n42657), .Y(n32148) );
  XOR2X1 U46409 ( .A(n41960), .B(n36899), .Y(n32152) );
  XOR2X1 U46410 ( .A(n41961), .B(n42605), .Y(n32144) );
  XOR2X1 U46411 ( .A(n41946), .B(n36756), .Y(n21757) );
  XOR2X1 U46412 ( .A(n41947), .B(n36757), .Y(n21697) );
  XOR2X1 U46413 ( .A(n41962), .B(n36761), .Y(n21413) );
  XOR2X1 U46414 ( .A(n41963), .B(n41309), .Y(n22693) );
  XOR2X1 U46415 ( .A(n41961), .B(n36755), .Y(n21423) );
  XOR2X1 U46416 ( .A(n41960), .B(n42517), .Y(n30931) );
  XNOR2X1 U46417 ( .A(n51334), .B(n41300), .Y(n22816) );
  XNOR2X1 U46418 ( .A(n51334), .B(n36742), .Y(n21759) );
  XNOR2X1 U46419 ( .A(n51333), .B(n36746), .Y(n21699) );
  XNOR2X1 U46420 ( .A(n50479), .B(n42579), .Y(n31835) );
  XOR2X1 U46421 ( .A(n42205), .B(n42487), .Y(n21758) );
  XOR2X1 U46422 ( .A(n42206), .B(n42487), .Y(n21698) );
  XOR2X1 U46423 ( .A(n42221), .B(n42485), .Y(n21414) );
  XOR2X1 U46424 ( .A(n42222), .B(n36813), .Y(n22694) );
  XOR2X1 U46425 ( .A(n42220), .B(n42485), .Y(n21424) );
  XOR2X1 U46426 ( .A(n42219), .B(n36801), .Y(n30932) );
  NOR4X1 U46427 ( .A(n21564), .B(n21563), .C(n21562), .D(n21561), .Y(n46725)
         );
  NOR4X1 U46428 ( .A(n32243), .B(n32244), .C(n32245), .D(n32246), .Y(n43055)
         );
  NOR4X1 U46429 ( .A(n32213), .B(n32214), .C(n32215), .D(n32216), .Y(n43064)
         );
  NOR4X1 U46430 ( .A(n32033), .B(n32034), .C(n32035), .D(n32036), .Y(n43127)
         );
  NOR4X1 U46431 ( .A(n32363), .B(n32364), .C(n32365), .D(n32366), .Y(n43073)
         );
  NOR4X1 U46432 ( .A(n31973), .B(n31974), .C(n31975), .D(n31976), .Y(n43137)
         );
  NOR4X1 U46433 ( .A(n32093), .B(n32094), .C(n32095), .D(n32096), .Y(n43109)
         );
  NOR4X1 U46434 ( .A(n32003), .B(n32004), .C(n32005), .D(n32006), .Y(n43132)
         );
  NOR4X1 U46435 ( .A(n31943), .B(n31944), .C(n31945), .D(n31946), .Y(n43146)
         );
  NOR4X1 U46436 ( .A(n32063), .B(n32064), .C(n32065), .D(n32066), .Y(n43118)
         );
  NOR4X1 U46437 ( .A(n32303), .B(n32304), .C(n32305), .D(n32306), .Y(n43045)
         );
  NOR4X1 U46438 ( .A(n32273), .B(n32274), .C(n32275), .D(n32276), .Y(n43050)
         );
  NOR4X1 U46439 ( .A(n31913), .B(n31914), .C(n31915), .D(n31916), .Y(n44586)
         );
  NOR4X1 U46440 ( .A(n32183), .B(n32184), .C(n32185), .D(n32186), .Y(n43083)
         );
  NOR4X1 U46441 ( .A(n32153), .B(n32154), .C(n32155), .D(n32156), .Y(n43092)
         );
  XNOR2X1 U46442 ( .A(n51320), .B(n42697), .Y(n32155) );
  NOR4X1 U46443 ( .A(n32123), .B(n32124), .C(n32125), .D(n32126), .Y(n43100)
         );
  NOR4X1 U46444 ( .A(n30856), .B(n30857), .C(n30858), .D(n30859), .Y(net216461) );
  NOR4X1 U46445 ( .A(n32329), .B(n32330), .C(n32331), .D(n32332), .Y(n43079)
         );
  NOR4X1 U46446 ( .A(n30796), .B(n30797), .C(n30798), .D(n30799), .Y(n43402)
         );
  NOR4X1 U46447 ( .A(n30766), .B(n30767), .C(n30768), .D(n30769), .Y(net216515) );
  NOR4X1 U46448 ( .A(n30946), .B(n30947), .C(n30948), .D(n30949), .Y(n43393)
         );
  NOR4X1 U46449 ( .A(n30736), .B(n30737), .C(n30738), .D(n30739), .Y(net216506) );
  NOR4X1 U46450 ( .A(n30706), .B(n30707), .C(n30708), .D(n30709), .Y(net216497) );
  NOR4X1 U46451 ( .A(n30886), .B(n30887), .C(n30888), .D(n30889), .Y(net216470) );
  CLKINVX1 U46452 ( .A(n10997), .Y(net209151) );
  AND2X2 U46453 ( .A(n11217), .B(n40395), .Y(n11009) );
  OAI221XL U46454 ( .A0(n9699), .A1(n50148), .B0(n50085), .B1(n9702), .C0(
        n9703), .Y(nxt_data_num[3]) );
  AOI221XL U46455 ( .A0(n9689), .A1(n50147), .B0(n41790), .B1(n50133), .C0(
        n9724), .Y(n9699) );
  AOI222XL U46456 ( .A0(n9704), .A1(n9705), .B0(n9706), .B1(n50148), .C0(n9679), .C1(n9707), .Y(n9703) );
  CLKINVX1 U46457 ( .A(n9721), .Y(n50085) );
  OAI222XL U46458 ( .A0(net266633), .A1(n42052), .B0(n40160), .B1(n42053),
        .C0(n40291), .C1(n42054), .Y(n13176) );
  OAI222XL U46459 ( .A0(net266633), .A1(n42311), .B0(n40160), .B1(n42312),
        .C0(n40292), .C1(n42313), .Y(n13164) );
  NOR2X1 U46460 ( .A(n39916), .B(n10661), .Y(n21608) );
  AND2X2 U46461 ( .A(n10683), .B(n10754), .Y(n21689) );
  NOR4X1 U46462 ( .A(n10223), .B(n10228), .C(n10227), .D(n22635), .Y(n9859) );
  NAND4X1 U46463 ( .A(n10806), .B(n10807), .C(n10808), .D(n22554), .Y(n9854)
         );
  NOR2X1 U46464 ( .A(net151509), .B(n10902), .Y(n22554) );
  NAND4X1 U46465 ( .A(n10903), .B(n10905), .C(n10904), .D(n22473), .Y(n9855)
         );
  NOR2BX1 U46466 ( .AN(n10706), .B(n10705), .Y(n19649) );
  NAND4X1 U46467 ( .A(n10771), .B(n10772), .C(n10776), .D(n23280), .Y(n9870)
         );
  NOR2X1 U46468 ( .A(n11228), .B(n10775), .Y(n23280) );
  NOR2X1 U46469 ( .A(net151530), .B(n10758), .Y(n21204) );
  OAI211X1 U46470 ( .A0(n9715), .A1(n50082), .B0(n43044), .C0(n43042), .Y(
        n9705) );
  AOI222XL U46471 ( .A0(net265644), .A1(n51227), .B0(n40209), .B1(n51226),
        .C0(net216978), .C1(n51225), .Y(n13118) );
  AOI222XL U46472 ( .A0(net265644), .A1(n51013), .B0(n40214), .B1(n51012),
        .C0(net216978), .C1(n51011), .Y(n13121) );
  AOI222XL U46473 ( .A0(net265644), .A1(n50799), .B0(n40214), .B1(n50798),
        .C0(net216978), .C1(n50797), .Y(n13124) );
  OAI211X1 U46474 ( .A0(n41809), .A1(n42816), .B0(n19102), .C0(n49570), .Y(
        n36540) );
  OA22X1 U46475 ( .A0(net262551), .A1(n41811), .B0(n41810), .B1(n40086), .Y(
        n19102) );
  CLKINVX1 U46476 ( .A(n19104), .Y(n49570) );
  OAI222XL U46477 ( .A0(net266402), .A1(n41806), .B0(n40174), .B1(n41807),
        .C0(n40303), .C1(n41808), .Y(n19104) );
  OA22X1 U46478 ( .A0(net262551), .A1(n41812), .B0(n41811), .B1(n40117), .Y(
        n19078) );
  CLKINVX1 U46479 ( .A(n19080), .Y(n49572) );
  OAI222XL U46480 ( .A0(net266402), .A1(n41807), .B0(n40174), .B1(n41808),
        .C0(n40303), .C1(n41809), .Y(n19080) );
  OA22X1 U46481 ( .A0(net262570), .A1(n41813), .B0(n41812), .B1(n40117), .Y(
        n19054) );
  CLKINVX1 U46482 ( .A(n19056), .Y(n49574) );
  OAI222XL U46483 ( .A0(net266402), .A1(n41808), .B0(n40174), .B1(n41809),
        .C0(n40302), .C1(n41810), .Y(n19056) );
  OAI211X1 U46484 ( .A0(n41812), .A1(n42817), .B0(n19030), .C0(n49576), .Y(
        n36516) );
  OA22X1 U46485 ( .A0(net262570), .A1(n34351), .B0(n41813), .B1(n40116), .Y(
        n19030) );
  CLKINVX1 U46486 ( .A(n19032), .Y(n49576) );
  OAI222XL U46487 ( .A0(net266402), .A1(n41809), .B0(n40174), .B1(n41810),
        .C0(n40302), .C1(n41811), .Y(n19032) );
  OA22X1 U46488 ( .A0(net262570), .A1(n41814), .B0(n34351), .B1(n40116), .Y(
        n19006) );
  CLKINVX1 U46489 ( .A(n19008), .Y(n49578) );
  OAI222XL U46490 ( .A0(net266402), .A1(n41810), .B0(n40173), .B1(n41811),
        .C0(n40302), .C1(n41812), .Y(n19008) );
  OA22X1 U46491 ( .A0(net262589), .A1(n41815), .B0(n41814), .B1(n40115), .Y(
        n18982) );
  CLKINVX1 U46492 ( .A(n18984), .Y(n49580) );
  OAI222XL U46493 ( .A0(net266402), .A1(n41811), .B0(n40173), .B1(n41812),
        .C0(n40302), .C1(n41813), .Y(n18984) );
  OAI211X1 U46494 ( .A0(n41814), .A1(n42818), .B0(n18958), .C0(n49582), .Y(
        n36492) );
  OA22X1 U46495 ( .A0(net262589), .A1(n41816), .B0(n41815), .B1(n40115), .Y(
        n18958) );
  CLKINVX1 U46496 ( .A(n18960), .Y(n49582) );
  OAI222XL U46497 ( .A0(net266402), .A1(n41812), .B0(n40173), .B1(n41813),
        .C0(n40302), .C1(n34351), .Y(n18960) );
  OA22X1 U46498 ( .A0(net262608), .A1(n41817), .B0(n41816), .B1(n40114), .Y(
        n18934) );
  CLKINVX1 U46499 ( .A(n18936), .Y(n49584) );
  OAI222XL U46500 ( .A0(net266402), .A1(n41813), .B0(n40173), .B1(n34351),
        .C0(n40302), .C1(n41814), .Y(n18936) );
  OA22X1 U46501 ( .A0(net262608), .A1(n41818), .B0(n41817), .B1(n40114), .Y(
        n18910) );
  CLKINVX1 U46502 ( .A(n18912), .Y(n49586) );
  OAI222XL U46503 ( .A0(net266423), .A1(n34351), .B0(n40173), .B1(n41814),
        .C0(n40302), .C1(n41815), .Y(n18912) );
  OA22X1 U46504 ( .A0(net262627), .A1(n41819), .B0(n41818), .B1(n40113), .Y(
        n18886) );
  CLKINVX1 U46505 ( .A(n18888), .Y(n49588) );
  OAI222XL U46506 ( .A0(net266423), .A1(n41814), .B0(n40173), .B1(n41815),
        .C0(n40302), .C1(n41816), .Y(n18888) );
  OAI211X1 U46507 ( .A0(n41818), .A1(n42819), .B0(n18862), .C0(n49590), .Y(
        n36460) );
  OA22X1 U46508 ( .A0(net262627), .A1(n41820), .B0(n41819), .B1(n40113), .Y(
        n18862) );
  CLKINVX1 U46509 ( .A(n18864), .Y(n49590) );
  OAI222XL U46510 ( .A0(net266423), .A1(n41815), .B0(n40173), .B1(n41816),
        .C0(n40302), .C1(n41817), .Y(n18864) );
  OA22X1 U46511 ( .A0(net262646), .A1(n41821), .B0(n41820), .B1(n40112), .Y(
        n18838) );
  CLKINVX1 U46512 ( .A(n18840), .Y(n49592) );
  OAI222XL U46513 ( .A0(net266423), .A1(n41816), .B0(n40173), .B1(n41817),
        .C0(n40301), .C1(n41818), .Y(n18840) );
  OA22X1 U46514 ( .A0(net262646), .A1(n41822), .B0(n41821), .B1(n40112), .Y(
        n18814) );
  CLKINVX1 U46515 ( .A(n18816), .Y(n49594) );
  OAI222XL U46516 ( .A0(net266423), .A1(n41817), .B0(n40172), .B1(n41818),
        .C0(n40301), .C1(n41819), .Y(n18816) );
  OAI211X1 U46517 ( .A0(n41821), .A1(n42820), .B0(n18790), .C0(n49596), .Y(
        n36436) );
  OA22X1 U46518 ( .A0(net262456), .A1(n41823), .B0(n41822), .B1(n40129), .Y(
        n18790) );
  CLKINVX1 U46519 ( .A(n18792), .Y(n49596) );
  OAI222XL U46520 ( .A0(net266423), .A1(n41818), .B0(n40172), .B1(n41819),
        .C0(n40301), .C1(n41820), .Y(n18792) );
  OA22X1 U46521 ( .A0(net262399), .A1(n41824), .B0(n41823), .B1(n40123), .Y(
        n18766) );
  CLKINVX1 U46522 ( .A(n18768), .Y(n49598) );
  OAI222XL U46523 ( .A0(net266423), .A1(n41819), .B0(n40172), .B1(n41820),
        .C0(n40301), .C1(n41821), .Y(n18768) );
  OA22X1 U46524 ( .A0(net262399), .A1(n41825), .B0(n41824), .B1(n40122), .Y(
        n18742) );
  CLKINVX1 U46525 ( .A(n18744), .Y(n49600) );
  OAI222XL U46526 ( .A0(net266423), .A1(n41820), .B0(n40172), .B1(n41821),
        .C0(n40301), .C1(n41822), .Y(n18744) );
  OA22X1 U46527 ( .A0(net262418), .A1(n41826), .B0(n41825), .B1(n40122), .Y(
        n18718) );
  CLKINVX1 U46528 ( .A(n18720), .Y(n49602) );
  OAI222XL U46529 ( .A0(net266423), .A1(n41821), .B0(n40172), .B1(n41822),
        .C0(n40301), .C1(n41823), .Y(n18720) );
  OAI211X1 U46530 ( .A0(n41825), .A1(n42821), .B0(n18694), .C0(n49604), .Y(
        n36404) );
  OA22X1 U46531 ( .A0(net262418), .A1(n41827), .B0(n41826), .B1(n40121), .Y(
        n18694) );
  CLKINVX1 U46532 ( .A(n18696), .Y(n49604) );
  OAI222XL U46533 ( .A0(net266423), .A1(n41822), .B0(n40172), .B1(n41823),
        .C0(n40301), .C1(n41824), .Y(n18696) );
  OA22X1 U46534 ( .A0(net262418), .A1(n41828), .B0(n41827), .B1(n40121), .Y(
        n18670) );
  CLKINVX1 U46535 ( .A(n18672), .Y(n49606) );
  OAI222XL U46536 ( .A0(net266444), .A1(n41823), .B0(n40172), .B1(n41824),
        .C0(n40301), .C1(n41825), .Y(n18672) );
  OA22X1 U46537 ( .A0(net262437), .A1(n41829), .B0(n41828), .B1(n40120), .Y(
        n18646) );
  CLKINVX1 U46538 ( .A(n18648), .Y(n49608) );
  OAI222XL U46539 ( .A0(net266444), .A1(n41824), .B0(n40172), .B1(n41825),
        .C0(n40301), .C1(n41826), .Y(n18648) );
  OAI211X1 U46540 ( .A0(n41828), .A1(n42822), .B0(n18622), .C0(n49610), .Y(
        n36380) );
  OA22X1 U46541 ( .A0(net262437), .A1(n41830), .B0(n41829), .B1(n40120), .Y(
        n18622) );
  CLKINVX1 U46542 ( .A(n18624), .Y(n49610) );
  OAI222XL U46543 ( .A0(net266444), .A1(n41825), .B0(n40172), .B1(n41826),
        .C0(n40300), .C1(n41827), .Y(n18624) );
  OA22X1 U46544 ( .A0(net262456), .A1(n41831), .B0(n41830), .B1(net218914),
        .Y(n18598) );
  CLKINVX1 U46545 ( .A(n18600), .Y(n49612) );
  OAI222XL U46546 ( .A0(net266444), .A1(n41826), .B0(n40171), .B1(n41827),
        .C0(n40300), .C1(n41828), .Y(n18600) );
  OA22X1 U46547 ( .A0(net262456), .A1(n41832), .B0(n41831), .B1(net218866),
        .Y(n18574) );
  CLKINVX1 U46548 ( .A(n18576), .Y(n49614) );
  OAI222XL U46549 ( .A0(net266444), .A1(n41827), .B0(n40171), .B1(n41828),
        .C0(n40300), .C1(n41829), .Y(n18576) );
  OA22X1 U46550 ( .A0(net262475), .A1(n41833), .B0(n41832), .B1(n40119), .Y(
        n18550) );
  CLKINVX1 U46551 ( .A(n18552), .Y(n49616) );
  OAI222XL U46552 ( .A0(net266444), .A1(n41828), .B0(n40171), .B1(n41829),
        .C0(n40300), .C1(n41830), .Y(n18552) );
  OAI211X1 U46553 ( .A0(n41832), .A1(n42823), .B0(n18526), .C0(n49618), .Y(
        n36348) );
  OA22X1 U46554 ( .A0(net262475), .A1(n41834), .B0(n41833), .B1(n40119), .Y(
        n18526) );
  CLKINVX1 U46555 ( .A(n18528), .Y(n49618) );
  OAI222XL U46556 ( .A0(net266444), .A1(n41829), .B0(n40171), .B1(n41830),
        .C0(n40300), .C1(n41831), .Y(n18528) );
  OA22X1 U46557 ( .A0(net218494), .A1(n41835), .B0(n41834), .B1(net218752),
        .Y(n18502) );
  CLKINVX1 U46558 ( .A(n18504), .Y(n49620) );
  OAI222XL U46559 ( .A0(net266444), .A1(n41830), .B0(n40171), .B1(n41831),
        .C0(n40300), .C1(n41832), .Y(n18504) );
  OA22X1 U46560 ( .A0(net218420), .A1(n41836), .B0(n41835), .B1(net218658),
        .Y(n18478) );
  CLKINVX1 U46561 ( .A(n18480), .Y(n49622) );
  OAI222XL U46562 ( .A0(net266444), .A1(n41831), .B0(n40171), .B1(n41832),
        .C0(n40300), .C1(n41833), .Y(n18480) );
  OAI211X1 U46563 ( .A0(n41835), .A1(n42824), .B0(n18454), .C0(n49624), .Y(
        n36324) );
  OA22X1 U46564 ( .A0(net262513), .A1(n41837), .B0(n41836), .B1(n40118), .Y(
        n18454) );
  CLKINVX1 U46565 ( .A(n18456), .Y(n49624) );
  OAI222XL U46566 ( .A0(net266444), .A1(n41832), .B0(n40171), .B1(n41833),
        .C0(n40300), .C1(n41834), .Y(n18456) );
  OA22X1 U46567 ( .A0(net262513), .A1(n41838), .B0(n41837), .B1(n40118), .Y(
        n18430) );
  CLKINVX1 U46568 ( .A(n18432), .Y(n49626) );
  OAI222XL U46569 ( .A0(net266465), .A1(n41833), .B0(n40171), .B1(n41834),
        .C0(n40300), .C1(n41835), .Y(n18432) );
  OA22X1 U46570 ( .A0(net262855), .A1(n41839), .B0(n41838), .B1(n40103), .Y(
        n18406) );
  CLKINVX1 U46571 ( .A(n18408), .Y(n49628) );
  OAI222XL U46572 ( .A0(net266465), .A1(n41834), .B0(n40170), .B1(n41835),
        .C0(n40299), .C1(n41836), .Y(n18408) );
  OAI211X1 U46573 ( .A0(n41838), .A1(n42825), .B0(n18382), .C0(n49630), .Y(
        n36300) );
  OA22X1 U46574 ( .A0(net262798), .A1(n41840), .B0(n41839), .B1(n40106), .Y(
        n18382) );
  CLKINVX1 U46575 ( .A(n18384), .Y(n49630) );
  OAI222XL U46576 ( .A0(net266465), .A1(n41835), .B0(n40170), .B1(n41836),
        .C0(n40299), .C1(n41837), .Y(n18384) );
  OA22X1 U46577 ( .A0(net262798), .A1(n41841), .B0(n41840), .B1(n40105), .Y(
        n18358) );
  CLKINVX1 U46578 ( .A(n18360), .Y(n49632) );
  OAI222XL U46579 ( .A0(net266465), .A1(n41836), .B0(n40170), .B1(n41837),
        .C0(n40299), .C1(n41838), .Y(n18360) );
  OA22X1 U46580 ( .A0(net262817), .A1(n41842), .B0(n41841), .B1(n40105), .Y(
        n18334) );
  CLKINVX1 U46581 ( .A(n18336), .Y(n49634) );
  OAI222XL U46582 ( .A0(net266465), .A1(n41837), .B0(n40170), .B1(n41838),
        .C0(n40299), .C1(n41839), .Y(n18336) );
  OA22X1 U46583 ( .A0(net262817), .A1(n41843), .B0(n41842), .B1(net218790),
        .Y(n18310) );
  CLKINVX1 U46584 ( .A(n18312), .Y(n49636) );
  OAI222XL U46585 ( .A0(net266465), .A1(n41838), .B0(n40170), .B1(n41839),
        .C0(n40299), .C1(n41840), .Y(n18312) );
  OA22X1 U46586 ( .A0(net262836), .A1(n41844), .B0(n41843), .B1(net218902),
        .Y(n18286) );
  CLKINVX1 U46587 ( .A(n18288), .Y(n49638) );
  OAI222XL U46588 ( .A0(net266465), .A1(n41839), .B0(n40170), .B1(n41840),
        .C0(n40299), .C1(n41841), .Y(n18288) );
  OA22X1 U46589 ( .A0(net262836), .A1(n41845), .B0(n41844), .B1(n40104), .Y(
        n18262) );
  CLKINVX1 U46590 ( .A(n18264), .Y(n49640) );
  OAI222XL U46591 ( .A0(net266465), .A1(n41840), .B0(n40170), .B1(n41841),
        .C0(n40299), .C1(n41842), .Y(n18264) );
  OA22X1 U46592 ( .A0(net262855), .A1(n41846), .B0(n41845), .B1(n40104), .Y(
        n18238) );
  CLKINVX1 U46593 ( .A(n18240), .Y(n49642) );
  OAI222XL U46594 ( .A0(net266465), .A1(n41841), .B0(n40170), .B1(n41842),
        .C0(n40299), .C1(n41843), .Y(n18240) );
  OA22X1 U46595 ( .A0(net262855), .A1(n41847), .B0(n41846), .B1(n40103), .Y(
        n18214) );
  CLKINVX1 U46596 ( .A(n18216), .Y(n49644) );
  OAI222XL U46597 ( .A0(net266465), .A1(n41842), .B0(n40169), .B1(n41843),
        .C0(n40299), .C1(n41844), .Y(n18216) );
  OA22X1 U46598 ( .A0(net262874), .A1(n41848), .B0(n41847), .B1(n40103), .Y(
        n18190) );
  CLKINVX1 U46599 ( .A(n18192), .Y(n49646) );
  OAI222XL U46600 ( .A0(net266486), .A1(n41843), .B0(n40169), .B1(n41844),
        .C0(n40298), .C1(n41845), .Y(n18192) );
  OA22X1 U46601 ( .A0(net262874), .A1(n41849), .B0(n41848), .B1(n40102), .Y(
        n18166) );
  CLKINVX1 U46602 ( .A(n18168), .Y(n49648) );
  OAI222XL U46603 ( .A0(net266486), .A1(n41844), .B0(n40169), .B1(n41845),
        .C0(n40298), .C1(n41846), .Y(n18168) );
  OAI211X1 U46604 ( .A0(n41848), .A1(n42831), .B0(n18142), .C0(n49650), .Y(
        n36220) );
  OA22X1 U46605 ( .A0(net262893), .A1(n41850), .B0(n41849), .B1(n40102), .Y(
        n18142) );
  CLKINVX1 U46606 ( .A(n18144), .Y(n49650) );
  OAI222XL U46607 ( .A0(net266486), .A1(n41845), .B0(n40169), .B1(n41846),
        .C0(n40298), .C1(n41847), .Y(n18144) );
  OAI211X1 U46608 ( .A0(n41849), .A1(n42800), .B0(n18118), .C0(n49652), .Y(
        n36212) );
  OA22X1 U46609 ( .A0(net262893), .A1(n41851), .B0(n41850), .B1(n40132), .Y(
        n18118) );
  CLKINVX1 U46610 ( .A(n18120), .Y(n49652) );
  OAI222XL U46611 ( .A0(net266486), .A1(n41846), .B0(n40169), .B1(n41847),
        .C0(n40298), .C1(n41848), .Y(n18120) );
  OA22X1 U46612 ( .A0(net262893), .A1(n41852), .B0(n41851), .B1(n40072), .Y(
        n18094) );
  CLKINVX1 U46613 ( .A(n18096), .Y(n49654) );
  OAI222XL U46614 ( .A0(net266486), .A1(n41847), .B0(n40169), .B1(n41848),
        .C0(n40298), .C1(n41849), .Y(n18096) );
  OA22X1 U46615 ( .A0(net262912), .A1(n41853), .B0(n41852), .B1(n40101), .Y(
        n18070) );
  CLKINVX1 U46616 ( .A(n18072), .Y(n49656) );
  OAI222XL U46617 ( .A0(net266486), .A1(n41848), .B0(n40169), .B1(n41849),
        .C0(n40298), .C1(n41850), .Y(n18072) );
  OA22X1 U46618 ( .A0(net262912), .A1(n41854), .B0(n41853), .B1(n40101), .Y(
        n18046) );
  CLKINVX1 U46619 ( .A(n18048), .Y(n49658) );
  OAI222XL U46620 ( .A0(net266486), .A1(n41849), .B0(n40169), .B1(n41850),
        .C0(n40298), .C1(n41851), .Y(n18048) );
  OA22X1 U46621 ( .A0(net262665), .A1(n41855), .B0(n41854), .B1(n40066), .Y(
        n18022) );
  CLKINVX1 U46622 ( .A(n18024), .Y(n49660) );
  OAI222XL U46623 ( .A0(net266486), .A1(n41850), .B0(n40169), .B1(n41851),
        .C0(n40298), .C1(n41852), .Y(n18024) );
  OA22X1 U46624 ( .A0(net262665), .A1(n41856), .B0(n41855), .B1(n40061), .Y(
        n17998) );
  CLKINVX1 U46625 ( .A(n18000), .Y(n49662) );
  OAI222XL U46626 ( .A0(net266486), .A1(n41851), .B0(n40168), .B1(n41852),
        .C0(n40297), .C1(n41853), .Y(n18000) );
  OAI211X1 U46627 ( .A0(n41855), .A1(n42806), .B0(n17974), .C0(n49664), .Y(
        n36164) );
  OA22X1 U46628 ( .A0(net262665), .A1(n41857), .B0(n41856), .B1(n40111), .Y(
        n17974) );
  CLKINVX1 U46629 ( .A(n17976), .Y(n49664) );
  OAI222XL U46630 ( .A0(net266486), .A1(n41852), .B0(n40168), .B1(n41853),
        .C0(n40297), .C1(n41854), .Y(n17976) );
  OA22X1 U46631 ( .A0(net262798), .A1(n41858), .B0(n41857), .B1(n40111), .Y(
        n17950) );
  CLKINVX1 U46632 ( .A(n17952), .Y(n49666) );
  OAI222XL U46633 ( .A0(net266507), .A1(n41853), .B0(n40168), .B1(n41854),
        .C0(n40297), .C1(n41855), .Y(n17952) );
  OAI211X1 U46634 ( .A0(n41857), .A1(n42809), .B0(n17926), .C0(n49668), .Y(
        n36148) );
  OA22X1 U46635 ( .A0(net218416), .A1(n41859), .B0(n41858), .B1(n40110), .Y(
        n17926) );
  CLKINVX1 U46636 ( .A(n17928), .Y(n49668) );
  OAI222XL U46637 ( .A0(net266507), .A1(n41854), .B0(n40168), .B1(n41855),
        .C0(n40297), .C1(n41856), .Y(n17928) );
  OA22X1 U46638 ( .A0(net262703), .A1(n41860), .B0(n41859), .B1(n40110), .Y(
        n17902) );
  CLKINVX1 U46639 ( .A(n17904), .Y(n49670) );
  OAI222XL U46640 ( .A0(net266507), .A1(n41855), .B0(n40168), .B1(n41856),
        .C0(n40297), .C1(n41857), .Y(n17904) );
  OA22X1 U46641 ( .A0(net262703), .A1(n41861), .B0(n41860), .B1(n40109), .Y(
        n17878) );
  CLKINVX1 U46642 ( .A(n17880), .Y(n49672) );
  OAI222XL U46643 ( .A0(net266507), .A1(n41856), .B0(n40168), .B1(n41857),
        .C0(n40297), .C1(n41858), .Y(n17880) );
  OAI211X1 U46644 ( .A0(n41860), .A1(n42812), .B0(n17854), .C0(n49674), .Y(
        n36124) );
  OA22X1 U46645 ( .A0(net262722), .A1(n41862), .B0(n41861), .B1(n40109), .Y(
        n17854) );
  CLKINVX1 U46646 ( .A(n17856), .Y(n49674) );
  OAI222XL U46647 ( .A0(net266507), .A1(n41857), .B0(n40168), .B1(n41858),
        .C0(n40297), .C1(n41859), .Y(n17856) );
  OA22X1 U46648 ( .A0(net262722), .A1(n41863), .B0(n41862), .B1(net218840),
        .Y(n17830) );
  CLKINVX1 U46649 ( .A(n17832), .Y(n49676) );
  OAI222XL U46650 ( .A0(net266507), .A1(n41858), .B0(n40168), .B1(n41859),
        .C0(n40297), .C1(n41860), .Y(n17832) );
  OAI211X1 U46651 ( .A0(n41862), .A1(n42815), .B0(n17806), .C0(n49678), .Y(
        n36108) );
  OA22X1 U46652 ( .A0(net262741), .A1(n41864), .B0(n41863), .B1(n40058), .Y(
        n17806) );
  CLKINVX1 U46653 ( .A(n17808), .Y(n49678) );
  OAI222XL U46654 ( .A0(net266507), .A1(n41859), .B0(n40167), .B1(n41860),
        .C0(n40297), .C1(n41861), .Y(n17808) );
  OAI211X1 U46655 ( .A0(n41863), .A1(n42848), .B0(n17782), .C0(n49680), .Y(
        n36100) );
  OA22X1 U46656 ( .A0(net262741), .A1(n41865), .B0(n41864), .B1(n40108), .Y(
        n17782) );
  CLKINVX1 U46657 ( .A(n17784), .Y(n49680) );
  OAI222XL U46658 ( .A0(net266507), .A1(n41860), .B0(n40167), .B1(n41861),
        .C0(n40296), .C1(n41862), .Y(n17784) );
  OAI211X1 U46659 ( .A0(n41864), .A1(n42849), .B0(n17758), .C0(n49682), .Y(
        n36092) );
  OA22X1 U46660 ( .A0(net262741), .A1(n41866), .B0(n41865), .B1(n40108), .Y(
        n17758) );
  CLKINVX1 U46661 ( .A(n17760), .Y(n49682) );
  OAI222XL U46662 ( .A0(net266507), .A1(n41861), .B0(n40167), .B1(n41862),
        .C0(n40296), .C1(n41863), .Y(n17760) );
  OAI211X1 U46663 ( .A0(n41865), .A1(n42850), .B0(n17734), .C0(n49684), .Y(
        n36084) );
  OA22X1 U46664 ( .A0(net263349), .A1(n41867), .B0(n41866), .B1(net218628),
        .Y(n17734) );
  CLKINVX1 U46665 ( .A(n17736), .Y(n49684) );
  OAI222XL U46666 ( .A0(net266507), .A1(n41862), .B0(n40167), .B1(n41863),
        .C0(n40296), .C1(n41864), .Y(n17736) );
  OAI211X1 U46667 ( .A0(n41866), .A1(n42851), .B0(n17710), .C0(n49686), .Y(
        n36076) );
  OA22X1 U46668 ( .A0(net263444), .A1(n41868), .B0(n41867), .B1(net218632),
        .Y(n17710) );
  CLKINVX1 U46669 ( .A(n17712), .Y(n49686) );
  OAI222XL U46670 ( .A0(net266528), .A1(n41863), .B0(n40167), .B1(n41864),
        .C0(n40296), .C1(n41865), .Y(n17712) );
  OA22X1 U46671 ( .A0(net262779), .A1(n41869), .B0(n41868), .B1(n40107), .Y(
        n17686) );
  CLKINVX1 U46672 ( .A(n17688), .Y(n49688) );
  OAI222XL U46673 ( .A0(net266528), .A1(n41864), .B0(n40167), .B1(n41865),
        .C0(n40296), .C1(n41866), .Y(n17688) );
  OA22X1 U46674 ( .A0(net262779), .A1(n41870), .B0(n41869), .B1(n40107), .Y(
        n17662) );
  CLKINVX1 U46675 ( .A(n17664), .Y(n49690) );
  OAI222XL U46676 ( .A0(net266318), .A1(n41865), .B0(n40178), .B1(n41866),
        .C0(n40296), .C1(n41867), .Y(n17664) );
  OAI211X1 U46677 ( .A0(n41869), .A1(n42855), .B0(n17638), .C0(n49692), .Y(
        n36052) );
  OA22X1 U46678 ( .A0(net262038), .A1(n41871), .B0(n41870), .B1(n40141), .Y(
        n17638) );
  CLKINVX1 U46679 ( .A(n17640), .Y(n49692) );
  OAI222XL U46680 ( .A0(net266318), .A1(n41866), .B0(n40178), .B1(n41867),
        .C0(n40296), .C1(n41868), .Y(n17640) );
  OA22X1 U46681 ( .A0(net261981), .A1(n41872), .B0(n41871), .B1(n40144), .Y(
        n17614) );
  CLKINVX1 U46682 ( .A(n17616), .Y(n49694) );
  OAI222XL U46683 ( .A0(net266318), .A1(n41867), .B0(n40179), .B1(n41868),
        .C0(n40296), .C1(n41869), .Y(n17616) );
  OA22X1 U46684 ( .A0(net262000), .A1(n41873), .B0(n41872), .B1(n40143), .Y(
        n17590) );
  CLKINVX1 U46685 ( .A(n17592), .Y(n49696) );
  OAI222XL U46686 ( .A0(net266318), .A1(n41868), .B0(n40179), .B1(n41869),
        .C0(n40296), .C1(n41870), .Y(n17592) );
  OA22X1 U46687 ( .A0(net262000), .A1(n41874), .B0(n41873), .B1(n40143), .Y(
        n17566) );
  CLKINVX1 U46688 ( .A(n17568), .Y(n49698) );
  OAI222XL U46689 ( .A0(net266297), .A1(n41869), .B0(n40179), .B1(n41870),
        .C0(n40295), .C1(n41871), .Y(n17568) );
  OA22X1 U46690 ( .A0(net262019), .A1(n41875), .B0(n41874), .B1(net218834),
        .Y(n17542) );
  CLKINVX1 U46691 ( .A(n17544), .Y(n49700) );
  OAI222XL U46692 ( .A0(net266297), .A1(n41870), .B0(n40179), .B1(n41871),
        .C0(n40295), .C1(n41872), .Y(n17544) );
  OA22X1 U46693 ( .A0(net262019), .A1(n41876), .B0(n41875), .B1(net218830),
        .Y(n17518) );
  CLKINVX1 U46694 ( .A(n17520), .Y(n49702) );
  OAI222XL U46695 ( .A0(net266297), .A1(n41871), .B0(n40179), .B1(n41872),
        .C0(n40295), .C1(n41873), .Y(n17520) );
  OAI211X1 U46696 ( .A0(n41875), .A1(n42862), .B0(n17494), .C0(n49704), .Y(
        n36004) );
  OA22X1 U46697 ( .A0(net262038), .A1(n41877), .B0(n41876), .B1(n40142), .Y(
        n17494) );
  CLKINVX1 U46698 ( .A(n17496), .Y(n49704) );
  OAI222XL U46699 ( .A0(net266297), .A1(n41872), .B0(n40179), .B1(n41873),
        .C0(n40295), .C1(n41874), .Y(n17496) );
  OA22X1 U46700 ( .A0(net262038), .A1(n41878), .B0(n41877), .B1(n40142), .Y(
        n17470) );
  CLKINVX1 U46701 ( .A(n17472), .Y(n49706) );
  OAI222XL U46702 ( .A0(net266297), .A1(n41873), .B0(n40179), .B1(n41874),
        .C0(n40295), .C1(n41875), .Y(n17472) );
  OAI211X1 U46703 ( .A0(n41877), .A1(n42832), .B0(n17446), .C0(n49708), .Y(
        n35988) );
  OA22X1 U46704 ( .A0(net262057), .A1(n41879), .B0(n41878), .B1(n40141), .Y(
        n17446) );
  CLKINVX1 U46705 ( .A(n17448), .Y(n49708) );
  OAI222XL U46706 ( .A0(net266297), .A1(n41874), .B0(n40179), .B1(n41875),
        .C0(n40295), .C1(n41876), .Y(n17448) );
  OAI211X1 U46707 ( .A0(n41878), .A1(n42833), .B0(n17422), .C0(n49710), .Y(
        n35980) );
  OA22X1 U46708 ( .A0(net262057), .A1(n41880), .B0(n41879), .B1(n40141), .Y(
        n17422) );
  CLKINVX1 U46709 ( .A(n17424), .Y(n49710) );
  OAI222XL U46710 ( .A0(net266297), .A1(n41875), .B0(n40180), .B1(n41876),
        .C0(n40295), .C1(n41877), .Y(n17424) );
  OAI211X1 U46711 ( .A0(n41879), .A1(n42834), .B0(n17398), .C0(n49712), .Y(
        n35972) );
  OA22X1 U46712 ( .A0(net262057), .A1(n41881), .B0(n41880), .B1(n40140), .Y(
        n17398) );
  CLKINVX1 U46713 ( .A(n17400), .Y(n49712) );
  OAI222XL U46714 ( .A0(net266297), .A1(n41876), .B0(n40180), .B1(n41877),
        .C0(n40295), .C1(n41878), .Y(n17400) );
  OAI211X1 U46715 ( .A0(n41880), .A1(n42835), .B0(n17374), .C0(n49714), .Y(
        n35964) );
  OA22X1 U46716 ( .A0(net263235), .A1(n41882), .B0(n41881), .B1(n40140), .Y(
        n17374) );
  CLKINVX1 U46717 ( .A(n17376), .Y(n49714) );
  OAI222XL U46718 ( .A0(net266297), .A1(n41877), .B0(n40180), .B1(n41878),
        .C0(n40295), .C1(n41879), .Y(n17376) );
  OAI211X1 U46719 ( .A0(n41881), .A1(n42836), .B0(n17350), .C0(n49716), .Y(
        n35956) );
  OA22X1 U46720 ( .A0(net263235), .A1(n41883), .B0(n41882), .B1(n40088), .Y(
        n17350) );
  CLKINVX1 U46721 ( .A(n17352), .Y(n49716) );
  OAI222XL U46722 ( .A0(net266297), .A1(n41878), .B0(n40180), .B1(n41879),
        .C0(n40294), .C1(n41880), .Y(n17352) );
  OAI211X1 U46723 ( .A0(n41882), .A1(n42837), .B0(n17326), .C0(n49718), .Y(
        n35948) );
  OA22X1 U46724 ( .A0(net262095), .A1(n41884), .B0(n41883), .B1(n40088), .Y(
        n17326) );
  CLKINVX1 U46725 ( .A(n17328), .Y(n49718) );
  OAI222XL U46726 ( .A0(net266276), .A1(n41879), .B0(n40180), .B1(n41880),
        .C0(n40294), .C1(n41881), .Y(n17328) );
  OAI211X1 U46727 ( .A0(n41883), .A1(n42839), .B0(n17302), .C0(n49720), .Y(
        n35940) );
  OA22X1 U46728 ( .A0(net262095), .A1(n41885), .B0(n41884), .B1(n40139), .Y(
        n17302) );
  CLKINVX1 U46729 ( .A(n17304), .Y(n49720) );
  OAI222XL U46730 ( .A0(net266276), .A1(n41880), .B0(n40180), .B1(n41881),
        .C0(n40294), .C1(n41882), .Y(n17304) );
  OAI211X1 U46731 ( .A0(n41884), .A1(n42840), .B0(n17278), .C0(n49722), .Y(
        n35932) );
  OA22X1 U46732 ( .A0(net262114), .A1(n41886), .B0(n41885), .B1(n40139), .Y(
        n17278) );
  CLKINVX1 U46733 ( .A(n17280), .Y(n49722) );
  OAI222XL U46734 ( .A0(net266276), .A1(n41881), .B0(n40180), .B1(n41882),
        .C0(n40294), .C1(n41883), .Y(n17280) );
  OAI211X1 U46735 ( .A0(n41885), .A1(n42841), .B0(n17254), .C0(n49724), .Y(
        n35924) );
  CLKINVX1 U46736 ( .A(n17256), .Y(n49724) );
  OAI222XL U46737 ( .A0(net266276), .A1(n41882), .B0(n40180), .B1(n41883),
        .C0(n40294), .C1(n41884), .Y(n17256) );
  OAI211X1 U46738 ( .A0(n41886), .A1(n42842), .B0(n17230), .C0(n49726), .Y(
        n35916) );
  CLKINVX1 U46739 ( .A(n17232), .Y(n49726) );
  OAI222XL U46740 ( .A0(net266276), .A1(n41883), .B0(n40181), .B1(n41884),
        .C0(n40294), .C1(n41885), .Y(n17232) );
  OAI211X1 U46741 ( .A0(n41887), .A1(n42843), .B0(n17206), .C0(n49728), .Y(
        n35908) );
  OA22X1 U46742 ( .A0(net261867), .A1(n41889), .B0(n41888), .B1(n40151), .Y(
        n17206) );
  CLKINVX1 U46743 ( .A(n17208), .Y(n49728) );
  OAI222XL U46744 ( .A0(net266276), .A1(n41884), .B0(n40181), .B1(n41885),
        .C0(n40294), .C1(n41886), .Y(n17208) );
  OAI211X1 U46745 ( .A0(n41888), .A1(n42844), .B0(n17182), .C0(n49730), .Y(
        n35900) );
  OA22X1 U46746 ( .A0(net261867), .A1(n41890), .B0(n41889), .B1(n40151), .Y(
        n17182) );
  CLKINVX1 U46747 ( .A(n17184), .Y(n49730) );
  OAI222XL U46748 ( .A0(net266276), .A1(n41885), .B0(n40181), .B1(n41886),
        .C0(n40294), .C1(n41887), .Y(n17184) );
  OA22X1 U46749 ( .A0(net261886), .A1(n41891), .B0(n41890), .B1(n40150), .Y(
        n17158) );
  CLKINVX1 U46750 ( .A(n17160), .Y(n49732) );
  OAI222XL U46751 ( .A0(net266276), .A1(n41886), .B0(n40181), .B1(n41887),
        .C0(n40294), .C1(n41888), .Y(n17160) );
  OA22X1 U46752 ( .A0(net261886), .A1(n41892), .B0(n41891), .B1(n40150), .Y(
        n17134) );
  CLKINVX1 U46753 ( .A(n17136), .Y(n49734) );
  OAI222XL U46754 ( .A0(net266276), .A1(n41887), .B0(n40181), .B1(n41888),
        .C0(n40293), .C1(n41889), .Y(n17136) );
  OAI211X1 U46755 ( .A0(n41891), .A1(n42751), .B0(n17110), .C0(n49736), .Y(
        n35876) );
  OA22X1 U46756 ( .A0(net261905), .A1(n41893), .B0(n41892), .B1(n40149), .Y(
        n17110) );
  CLKINVX1 U46757 ( .A(n17112), .Y(n49736) );
  OAI222XL U46758 ( .A0(net266276), .A1(n41888), .B0(n40181), .B1(n41889),
        .C0(n40293), .C1(n41890), .Y(n17112) );
  OA22X1 U46759 ( .A0(net261905), .A1(n41894), .B0(n41893), .B1(n40149), .Y(
        n17086) );
  CLKINVX1 U46760 ( .A(n17088), .Y(n49738) );
  OAI222XL U46761 ( .A0(net266255), .A1(n41889), .B0(n40181), .B1(n41890),
        .C0(n40293), .C1(n41891), .Y(n17088) );
  OA22X1 U46762 ( .A0(net261905), .A1(n41895), .B0(n41894), .B1(n40148), .Y(
        n17062) );
  CLKINVX1 U46763 ( .A(n17064), .Y(n49740) );
  OAI222XL U46764 ( .A0(net266255), .A1(n41890), .B0(n40181), .B1(n41891),
        .C0(n40293), .C1(n41892), .Y(n17064) );
  OAI211X1 U46765 ( .A0(n41894), .A1(n42754), .B0(n17038), .C0(n49742), .Y(
        n35852) );
  OA22X1 U46766 ( .A0(net261924), .A1(n41896), .B0(n41895), .B1(n40148), .Y(
        n17038) );
  CLKINVX1 U46767 ( .A(n17040), .Y(n49742) );
  OAI222XL U46768 ( .A0(net266255), .A1(n41891), .B0(n40181), .B1(n41892),
        .C0(n40293), .C1(n41893), .Y(n17040) );
  OA22X1 U46769 ( .A0(net261924), .A1(n41897), .B0(n41896), .B1(n40147), .Y(
        n17014) );
  CLKINVX1 U46770 ( .A(n17016), .Y(n49744) );
  OAI222XL U46771 ( .A0(net266255), .A1(n41892), .B0(n40182), .B1(n41893),
        .C0(n40293), .C1(n41894), .Y(n17016) );
  OAI211X1 U46772 ( .A0(n41896), .A1(n42757), .B0(n16990), .C0(n49746), .Y(
        n35836) );
  OA22X1 U46773 ( .A0(net261943), .A1(n41898), .B0(n41897), .B1(n40147), .Y(
        n16990) );
  CLKINVX1 U46774 ( .A(n16992), .Y(n49746) );
  OAI222XL U46775 ( .A0(net266255), .A1(n41893), .B0(n40182), .B1(n41894),
        .C0(n40293), .C1(n41895), .Y(n16992) );
  OAI211X1 U46776 ( .A0(n41897), .A1(n42758), .B0(n16966), .C0(n49748), .Y(
        n35828) );
  OA22X1 U46777 ( .A0(net261943), .A1(n41899), .B0(n41898), .B1(n40146), .Y(
        n16966) );
  CLKINVX1 U46778 ( .A(n16968), .Y(n49748) );
  OAI222XL U46779 ( .A0(net266255), .A1(n41894), .B0(n40182), .B1(n41895),
        .C0(n40293), .C1(n41896), .Y(n16968) );
  OAI211X1 U46780 ( .A0(n41898), .A1(n42759), .B0(n16942), .C0(n49750), .Y(
        n35820) );
  OA22X1 U46781 ( .A0(net218464), .A1(n41900), .B0(n41899), .B1(n40146), .Y(
        n16942) );
  CLKINVX1 U46782 ( .A(n16944), .Y(n49750) );
  OAI222XL U46783 ( .A0(net266255), .A1(n41895), .B0(n40182), .B1(n41896),
        .C0(n40293), .C1(n41897), .Y(n16944) );
  OAI211X1 U46784 ( .A0(n41899), .A1(n42760), .B0(n16918), .C0(n49752), .Y(
        n35812) );
  OA22X1 U46785 ( .A0(net218386), .A1(n41901), .B0(n41900), .B1(n40145), .Y(
        n16918) );
  CLKINVX1 U46786 ( .A(n16920), .Y(n49752) );
  OAI222XL U46787 ( .A0(net266255), .A1(n41896), .B0(n40182), .B1(n41897),
        .C0(n40292), .C1(n41898), .Y(n16920) );
  OAI211X1 U46788 ( .A0(n41900), .A1(n42761), .B0(n16894), .C0(n49754), .Y(
        n35804) );
  OA22X1 U46789 ( .A0(net261981), .A1(n41902), .B0(n41901), .B1(n40145), .Y(
        n16894) );
  CLKINVX1 U46790 ( .A(n16896), .Y(n49754) );
  OAI222XL U46791 ( .A0(net266318), .A1(n41897), .B0(n40180), .B1(n41898),
        .C0(n40311), .C1(n41899), .Y(n16896) );
  OA22X1 U46792 ( .A0(net262247), .A1(n41903), .B0(n41902), .B1(n40130), .Y(
        n16870) );
  CLKINVX1 U46793 ( .A(n16872), .Y(n49756) );
  OAI222XL U46794 ( .A0(net266318), .A1(n41898), .B0(n40178), .B1(n41899),
        .C0(net217128), .C1(n41900), .Y(n16872) );
  OA22X1 U46795 ( .A0(net262266), .A1(n41904), .B0(n41903), .B1(n40130), .Y(
        n16846) );
  CLKINVX1 U46796 ( .A(n16848), .Y(n49758) );
  OAI222XL U46797 ( .A0(net266318), .A1(n41899), .B0(n40178), .B1(n41900),
        .C0(net217166), .C1(n41901), .Y(n16848) );
  OA22X1 U46798 ( .A0(net262266), .A1(n41905), .B0(n41904), .B1(n40129), .Y(
        n16822) );
  CLKINVX1 U46799 ( .A(n16824), .Y(n49760) );
  OAI222XL U46800 ( .A0(net266318), .A1(n41900), .B0(n40178), .B1(n41901),
        .C0(net217244), .C1(n41902), .Y(n16824) );
  OAI211X1 U46801 ( .A0(n41904), .A1(n42766), .B0(n16798), .C0(n49762), .Y(
        n35772) );
  OA22X1 U46802 ( .A0(net262285), .A1(n41906), .B0(n41905), .B1(n40129), .Y(
        n16798) );
  CLKINVX1 U46803 ( .A(n16800), .Y(n49762) );
  OAI222XL U46804 ( .A0(net266318), .A1(n41901), .B0(n40178), .B1(n41902),
        .C0(net217140), .C1(n41903), .Y(n16800) );
  OAI211X1 U46805 ( .A0(n41905), .A1(n42736), .B0(n16774), .C0(n49764), .Y(
        n35764) );
  OA22X1 U46806 ( .A0(net262285), .A1(n41907), .B0(n41906), .B1(n40094), .Y(
        n16774) );
  CLKINVX1 U46807 ( .A(n16776), .Y(n49764) );
  OAI222XL U46808 ( .A0(net266318), .A1(n41902), .B0(n40178), .B1(n41903),
        .C0(net217138), .C1(n41904), .Y(n16776) );
  OA22X1 U46809 ( .A0(net262285), .A1(n41908), .B0(n41907), .B1(n40078), .Y(
        n16750) );
  CLKINVX1 U46810 ( .A(n16752), .Y(n49766) );
  OAI222XL U46811 ( .A0(net266339), .A1(n41903), .B0(n40178), .B1(n41904),
        .C0(net217146), .C1(n41905), .Y(n16752) );
  OA22X1 U46812 ( .A0(net262304), .A1(n41909), .B0(n41908), .B1(n40128), .Y(
        n16726) );
  CLKINVX1 U46813 ( .A(n16728), .Y(n49768) );
  OAI222XL U46814 ( .A0(net266339), .A1(n41904), .B0(n40178), .B1(n41905),
        .C0(net217154), .C1(n41906), .Y(n16728) );
  OA22X1 U46815 ( .A0(net262304), .A1(n41910), .B0(n41909), .B1(n40128), .Y(
        n16702) );
  CLKINVX1 U46816 ( .A(n16704), .Y(n49770) );
  OAI222XL U46817 ( .A0(net266339), .A1(n41905), .B0(n40177), .B1(n41906),
        .C0(n40309), .C1(n41907), .Y(n16704) );
  OA22X1 U46818 ( .A0(net262323), .A1(n41911), .B0(n41910), .B1(n40127), .Y(
        n16678) );
  CLKINVX1 U46819 ( .A(n16680), .Y(n49772) );
  OAI222XL U46820 ( .A0(net266339), .A1(n41906), .B0(n40177), .B1(n41907),
        .C0(n40309), .C1(n41908), .Y(n16680) );
  OAI211X1 U46821 ( .A0(n41910), .A1(n42741), .B0(n16654), .C0(n49774), .Y(
        n35724) );
  OA22X1 U46822 ( .A0(net262323), .A1(n41912), .B0(n41911), .B1(n40127), .Y(
        n16654) );
  CLKINVX1 U46823 ( .A(n16656), .Y(n49774) );
  OAI222XL U46824 ( .A0(net266339), .A1(n41907), .B0(n40177), .B1(n41908),
        .C0(n40309), .C1(n41909), .Y(n16656) );
  OAI211X1 U46825 ( .A0(n41911), .A1(n42742), .B0(n16630), .C0(n49776), .Y(
        n35716) );
  OA22X1 U46826 ( .A0(net262342), .A1(n41913), .B0(n41912), .B1(n40126), .Y(
        n16630) );
  CLKINVX1 U46827 ( .A(n16632), .Y(n49776) );
  OAI222XL U46828 ( .A0(net266339), .A1(n41908), .B0(n40177), .B1(n41909),
        .C0(n40309), .C1(n41910), .Y(n16632) );
  OAI211X1 U46829 ( .A0(n41912), .A1(n42743), .B0(n16606), .C0(n49778), .Y(
        n35708) );
  OA22X1 U46830 ( .A0(net262342), .A1(n41914), .B0(n41913), .B1(n40126), .Y(
        n16606) );
  CLKINVX1 U46831 ( .A(n16608), .Y(n49778) );
  OAI222XL U46832 ( .A0(net266339), .A1(n41909), .B0(n40177), .B1(n41910),
        .C0(n40309), .C1(n41911), .Y(n16608) );
  OAI211X1 U46833 ( .A0(n41913), .A1(n42744), .B0(n16582), .C0(n49780), .Y(
        n35700) );
  OA22X1 U46834 ( .A0(net262361), .A1(n41915), .B0(n41914), .B1(n40125), .Y(
        n16582) );
  CLKINVX1 U46835 ( .A(n16584), .Y(n49780) );
  OAI222XL U46836 ( .A0(net266339), .A1(n41910), .B0(n40177), .B1(n41911),
        .C0(n40309), .C1(n41912), .Y(n16584) );
  OA22X1 U46837 ( .A0(net262361), .A1(n41916), .B0(n41915), .B1(n40125), .Y(
        n16558) );
  CLKINVX1 U46838 ( .A(n16560), .Y(n49782) );
  OAI222XL U46839 ( .A0(net266339), .A1(n41911), .B0(n40177), .B1(n41912),
        .C0(n40309), .C1(n41913), .Y(n16560) );
  OA22X1 U46840 ( .A0(net262361), .A1(n41917), .B0(n41916), .B1(n40124), .Y(
        n16534) );
  CLKINVX1 U46841 ( .A(n16536), .Y(n49784) );
  OAI222XL U46842 ( .A0(net266339), .A1(n41912), .B0(n40177), .B1(n41913),
        .C0(n40309), .C1(n41914), .Y(n16536) );
  OA22X1 U46843 ( .A0(net262380), .A1(n41918), .B0(n41917), .B1(n40124), .Y(
        n16510) );
  CLKINVX1 U46844 ( .A(n16512), .Y(n49786) );
  OAI222XL U46845 ( .A0(net266360), .A1(n41913), .B0(n40176), .B1(n41914),
        .C0(n40309), .C1(n41915), .Y(n16512) );
  OA22X1 U46846 ( .A0(net262114), .A1(n41919), .B0(n41918), .B1(n40138), .Y(
        n16486) );
  CLKINVX1 U46847 ( .A(n16488), .Y(n49788) );
  OAI222XL U46848 ( .A0(net266360), .A1(n41914), .B0(n40176), .B1(n41915),
        .C0(n40310), .C1(n41916), .Y(n16488) );
  OA22X1 U46849 ( .A0(net262133), .A1(n41920), .B0(n41919), .B1(n40138), .Y(
        n16462) );
  CLKINVX1 U46850 ( .A(n16464), .Y(n49790) );
  OAI222XL U46851 ( .A0(net266360), .A1(n41915), .B0(n40176), .B1(n41916),
        .C0(n40310), .C1(n41917), .Y(n16464) );
  OA22X1 U46852 ( .A0(net262133), .A1(n41921), .B0(n41920), .B1(n40137), .Y(
        n16438) );
  CLKINVX1 U46853 ( .A(n16440), .Y(n49792) );
  OAI222XL U46854 ( .A0(net266360), .A1(n41916), .B0(n40176), .B1(n41917),
        .C0(n40310), .C1(n41918), .Y(n16440) );
  OA22X1 U46855 ( .A0(net262133), .A1(n41922), .B0(n41921), .B1(n40137), .Y(
        n16414) );
  CLKINVX1 U46856 ( .A(n16416), .Y(n49794) );
  OAI222XL U46857 ( .A0(net266360), .A1(n41917), .B0(n40176), .B1(n41918),
        .C0(n40310), .C1(n41919), .Y(n16416) );
  OAI211X1 U46858 ( .A0(n41921), .A1(n42785), .B0(n16390), .C0(n49796), .Y(
        n35636) );
  OA22X1 U46859 ( .A0(net262152), .A1(n41923), .B0(n41922), .B1(n40136), .Y(
        n16390) );
  CLKINVX1 U46860 ( .A(n16392), .Y(n49796) );
  OAI222XL U46861 ( .A0(net266360), .A1(n41918), .B0(n40176), .B1(n41919),
        .C0(n40310), .C1(n41920), .Y(n16392) );
  OAI211X1 U46862 ( .A0(n41922), .A1(n42787), .B0(n16366), .C0(n49798), .Y(
        n35628) );
  OA22X1 U46863 ( .A0(net262152), .A1(n41924), .B0(n41923), .B1(n40136), .Y(
        n16366) );
  CLKINVX1 U46864 ( .A(n16368), .Y(n49798) );
  OAI222XL U46865 ( .A0(net266360), .A1(n41919), .B0(n40176), .B1(n41920),
        .C0(n40310), .C1(n41921), .Y(n16368) );
  OAI211X1 U46866 ( .A0(n41923), .A1(n42788), .B0(n16342), .C0(n49800), .Y(
        n35620) );
  OA22X1 U46867 ( .A0(net262171), .A1(n41925), .B0(n41924), .B1(n40135), .Y(
        n16342) );
  CLKINVX1 U46868 ( .A(n16344), .Y(n49800) );
  OAI222XL U46869 ( .A0(net266360), .A1(n41920), .B0(n40176), .B1(n41921),
        .C0(n40310), .C1(n41922), .Y(n16344) );
  OA22X1 U46870 ( .A0(net262171), .A1(n41926), .B0(n41925), .B1(n40135), .Y(
        n16318) );
  CLKINVX1 U46871 ( .A(n16320), .Y(n49802) );
  OAI222XL U46872 ( .A0(net266360), .A1(n41921), .B0(n40176), .B1(n41922),
        .C0(n40310), .C1(n41923), .Y(n16320) );
  OA22X1 U46873 ( .A0(net262190), .A1(n41927), .B0(n41926), .B1(n40134), .Y(
        n16294) );
  CLKINVX1 U46874 ( .A(n16296), .Y(n49804) );
  OAI222XL U46875 ( .A0(net266360), .A1(n41922), .B0(n40175), .B1(n41923),
        .C0(n40311), .C1(n41924), .Y(n16296) );
  OA22X1 U46876 ( .A0(net262190), .A1(n41928), .B0(n41927), .B1(n40134), .Y(
        n16270) );
  CLKINVX1 U46877 ( .A(n16272), .Y(n49806) );
  OAI222XL U46878 ( .A0(net266381), .A1(n41923), .B0(n40175), .B1(n41924),
        .C0(n40310), .C1(n41925), .Y(n16272) );
  OA22X1 U46879 ( .A0(net262209), .A1(n41929), .B0(n41928), .B1(n40133), .Y(
        n16246) );
  CLKINVX1 U46880 ( .A(n16248), .Y(n49808) );
  OAI222XL U46881 ( .A0(net266381), .A1(n41924), .B0(n40175), .B1(n41925),
        .C0(n40311), .C1(n41926), .Y(n16248) );
  OA22X1 U46882 ( .A0(net262209), .A1(n41930), .B0(n41929), .B1(n40133), .Y(
        n16222) );
  CLKINVX1 U46883 ( .A(n16224), .Y(n49810) );
  OAI222XL U46884 ( .A0(net266381), .A1(n41925), .B0(n40175), .B1(n41926),
        .C0(n40311), .C1(n41927), .Y(n16224) );
  OA22X1 U46885 ( .A0(net262228), .A1(n41931), .B0(n41930), .B1(n40132), .Y(
        n16198) );
  CLKINVX1 U46886 ( .A(n16200), .Y(n49812) );
  OAI222XL U46887 ( .A0(net266381), .A1(n41926), .B0(n40175), .B1(n41927),
        .C0(n40311), .C1(n41928), .Y(n16200) );
  OA22X1 U46888 ( .A0(net262228), .A1(n41932), .B0(n41931), .B1(n40132), .Y(
        n16174) );
  CLKINVX1 U46889 ( .A(n16176), .Y(n49814) );
  OAI222XL U46890 ( .A0(net266381), .A1(n41927), .B0(n40175), .B1(n41928),
        .C0(n40311), .C1(n41929), .Y(n16176) );
  OA22X1 U46891 ( .A0(net262228), .A1(n41933), .B0(n41932), .B1(n40131), .Y(
        n16150) );
  CLKINVX1 U46892 ( .A(n16152), .Y(n49816) );
  OAI222XL U46893 ( .A0(net266381), .A1(n41928), .B0(n40175), .B1(n41929),
        .C0(n40311), .C1(n41930), .Y(n16152) );
  OA22X1 U46894 ( .A0(net262247), .A1(n41934), .B0(n41933), .B1(n40131), .Y(
        n16126) );
  CLKINVX1 U46895 ( .A(n16128), .Y(n49818) );
  OAI222XL U46896 ( .A0(net266381), .A1(n41929), .B0(n40175), .B1(n41930),
        .C0(n40311), .C1(n41931), .Y(n16128) );
  OA22X1 U46897 ( .A0(net263672), .A1(n41935), .B0(n41934), .B1(net218878),
        .Y(n16102) );
  CLKINVX1 U46898 ( .A(n16104), .Y(n49820) );
  OAI222XL U46899 ( .A0(net266738), .A1(n41930), .B0(n40174), .B1(n41931),
        .C0(n40311), .C1(n41932), .Y(n16104) );
  OAI211X1 U46900 ( .A0(n41934), .A1(n42768), .B0(n16078), .C0(n49822), .Y(
        n35532) );
  OA22X1 U46901 ( .A0(net263615), .A1(n41936), .B0(n41935), .B1(n40061), .Y(
        n16078) );
  CLKINVX1 U46902 ( .A(n16080), .Y(n49822) );
  OAI222XL U46903 ( .A0(net266654), .A1(n41931), .B0(n40159), .B1(n41932),
        .C0(n40312), .C1(n41933), .Y(n16080) );
  OA22X1 U46904 ( .A0(net263615), .A1(n41937), .B0(n41936), .B1(n40060), .Y(
        n16054) );
  CLKINVX1 U46905 ( .A(n16056), .Y(n49824) );
  OAI222XL U46906 ( .A0(net266654), .A1(n41932), .B0(n40159), .B1(n41933),
        .C0(n40311), .C1(n41934), .Y(n16056) );
  OA22X1 U46907 ( .A0(net263634), .A1(n41938), .B0(n41937), .B1(n40060), .Y(
        n16030) );
  CLKINVX1 U46908 ( .A(n16032), .Y(n49826) );
  OAI222XL U46909 ( .A0(net266675), .A1(n41933), .B0(n40159), .B1(n41934),
        .C0(n40312), .C1(n41935), .Y(n16032) );
  OA22X1 U46910 ( .A0(net263634), .A1(n41939), .B0(n41938), .B1(n40059), .Y(
        n16006) );
  CLKINVX1 U46911 ( .A(n16008), .Y(n49828) );
  OAI222XL U46912 ( .A0(net266675), .A1(n41934), .B0(n40159), .B1(n41935),
        .C0(n40312), .C1(n41936), .Y(n16008) );
  OA22X1 U46913 ( .A0(net263634), .A1(n41940), .B0(n41939), .B1(n40059), .Y(
        n15982) );
  CLKINVX1 U46914 ( .A(n15984), .Y(n49830) );
  OAI222XL U46915 ( .A0(net266675), .A1(n41935), .B0(n40159), .B1(n41936),
        .C0(n40312), .C1(n41937), .Y(n15984) );
  OA22X1 U46916 ( .A0(net263653), .A1(n41941), .B0(n41940), .B1(n40058), .Y(
        n15958) );
  CLKINVX1 U46917 ( .A(n15960), .Y(n49832) );
  OAI222XL U46918 ( .A0(net266675), .A1(n41936), .B0(n40158), .B1(n41937),
        .C0(n40312), .C1(n41938), .Y(n15960) );
  OA22X1 U46919 ( .A0(net263653), .A1(n41942), .B0(n41941), .B1(n40058), .Y(
        n15934) );
  CLKINVX1 U46920 ( .A(n15936), .Y(n49834) );
  OAI222XL U46921 ( .A0(net266675), .A1(n41937), .B0(n40158), .B1(n41938),
        .C0(n40312), .C1(n41939), .Y(n15936) );
  OA22X1 U46922 ( .A0(net263672), .A1(n41943), .B0(n41942), .B1(net218796),
        .Y(n15910) );
  CLKINVX1 U46923 ( .A(n15912), .Y(n49836) );
  OAI222XL U46924 ( .A0(net266675), .A1(n41938), .B0(n40158), .B1(n41939),
        .C0(n40312), .C1(n41940), .Y(n15912) );
  OAI211X1 U46925 ( .A0(n41942), .A1(n42777), .B0(n15886), .C0(n49838), .Y(
        n35468) );
  OA22X1 U46926 ( .A0(net263672), .A1(n41944), .B0(n41943), .B1(n40142), .Y(
        n15886) );
  CLKINVX1 U46927 ( .A(n15888), .Y(n49838) );
  OAI222XL U46928 ( .A0(net266675), .A1(n41939), .B0(n40158), .B1(n41940),
        .C0(n40312), .C1(n41941), .Y(n15888) );
  OA22X1 U46929 ( .A0(net263691), .A1(n41945), .B0(n41944), .B1(n40057), .Y(
        n15862) );
  CLKINVX1 U46930 ( .A(n15864), .Y(n49840) );
  OAI222XL U46931 ( .A0(net266675), .A1(n41940), .B0(n40158), .B1(n41941),
        .C0(n40313), .C1(n41942), .Y(n15864) );
  OA22X1 U46932 ( .A0(net263691), .A1(n41946), .B0(n41945), .B1(n40057), .Y(
        n15838) );
  CLKINVX1 U46933 ( .A(n15840), .Y(n49842) );
  OAI222XL U46934 ( .A0(net266675), .A1(n41941), .B0(n40158), .B1(n41942),
        .C0(n40312), .C1(n41943), .Y(n15840) );
  OAI211X1 U46935 ( .A0(n41945), .A1(n42781), .B0(n15814), .C0(n49844), .Y(
        n35444) );
  OA22X1 U46936 ( .A0(net263710), .A1(n41947), .B0(n41946), .B1(n40056), .Y(
        n15814) );
  CLKINVX1 U46937 ( .A(n15816), .Y(n49844) );
  OAI222XL U46938 ( .A0(net266675), .A1(n41942), .B0(n40158), .B1(n41943),
        .C0(n40310), .C1(n41944), .Y(n15816) );
  OA22X1 U46939 ( .A0(net263710), .A1(n41948), .B0(n41947), .B1(n40056), .Y(
        n15790) );
  CLKINVX1 U46940 ( .A(n15792), .Y(n49846) );
  OAI222XL U46941 ( .A0(net266696), .A1(n41943), .B0(n40158), .B1(n41944),
        .C0(n40308), .C1(n41945), .Y(n15792) );
  OA22X1 U46942 ( .A0(net218464), .A1(n41949), .B0(n41948), .B1(n40055), .Y(
        n15766) );
  CLKINVX1 U46943 ( .A(n15768), .Y(n49848) );
  OAI222XL U46944 ( .A0(net266696), .A1(n41944), .B0(n40157), .B1(n41945),
        .C0(n40308), .C1(n41946), .Y(n15768) );
  OA22X1 U46945 ( .A0(net218530), .A1(n41950), .B0(n41949), .B1(n40055), .Y(
        n15742) );
  CLKINVX1 U46946 ( .A(n15744), .Y(n49850) );
  OAI222XL U46947 ( .A0(net266696), .A1(n41945), .B0(n40157), .B1(n41946),
        .C0(n40308), .C1(n41947), .Y(n15744) );
  OA22X1 U46948 ( .A0(net263463), .A1(n41951), .B0(n41950), .B1(n40069), .Y(
        n15718) );
  CLKINVX1 U46949 ( .A(n15720), .Y(n49852) );
  OAI222XL U46950 ( .A0(net266696), .A1(n41946), .B0(n40157), .B1(n41947),
        .C0(n40308), .C1(n41948), .Y(n15720) );
  OA22X1 U46951 ( .A0(net218428), .A1(n41952), .B0(n41951), .B1(n40069), .Y(
        n15694) );
  CLKINVX1 U46952 ( .A(n15696), .Y(n49854) );
  OAI222XL U46953 ( .A0(net266696), .A1(n41947), .B0(n40157), .B1(n41948),
        .C0(n40308), .C1(n41949), .Y(n15696) );
  OA22X1 U46954 ( .A0(net218430), .A1(n41953), .B0(n41952), .B1(n40068), .Y(
        n15670) );
  CLKINVX1 U46955 ( .A(n15672), .Y(n49856) );
  OAI222XL U46956 ( .A0(net266696), .A1(n41948), .B0(n40157), .B1(n41949),
        .C0(n40308), .C1(n41950), .Y(n15672) );
  OA22X1 U46957 ( .A0(net263501), .A1(n41954), .B0(n41953), .B1(n40068), .Y(
        n15646) );
  CLKINVX1 U46958 ( .A(n15648), .Y(n49858) );
  OAI222XL U46959 ( .A0(net266696), .A1(n41949), .B0(n40157), .B1(n41950),
        .C0(n40308), .C1(n41951), .Y(n15648) );
  OA22X1 U46960 ( .A0(net263501), .A1(n41955), .B0(n41954), .B1(n40067), .Y(
        n15622) );
  CLKINVX1 U46961 ( .A(n15624), .Y(n49860) );
  OAI222XL U46962 ( .A0(net266696), .A1(n41950), .B0(n40157), .B1(n41951),
        .C0(n40308), .C1(n41952), .Y(n15624) );
  OAI211X1 U46963 ( .A0(n41954), .A1(n42952), .B0(n15598), .C0(n49862), .Y(
        n35372) );
  OA22X1 U46964 ( .A0(net263501), .A1(n41956), .B0(n41955), .B1(n40067), .Y(
        n15598) );
  CLKINVX1 U46965 ( .A(n15600), .Y(n49862) );
  OAI222XL U46966 ( .A0(net266696), .A1(n41951), .B0(n40157), .B1(n41952),
        .C0(n40308), .C1(n41953), .Y(n15600) );
  OA22X1 U46967 ( .A0(net218524), .A1(n41957), .B0(n41956), .B1(n40066), .Y(
        n15574) );
  CLKINVX1 U46968 ( .A(n15576), .Y(n49864) );
  OAI222XL U46969 ( .A0(net266696), .A1(n41952), .B0(n40157), .B1(n41953),
        .C0(n40307), .C1(n41954), .Y(n15576) );
  OA22X1 U46970 ( .A0(net218536), .A1(n41958), .B0(n41957), .B1(n40066), .Y(
        n15550) );
  CLKINVX1 U46971 ( .A(n15552), .Y(n49866) );
  OAI222XL U46972 ( .A0(net266717), .A1(n41953), .B0(n40156), .B1(n41954),
        .C0(n40307), .C1(n41955), .Y(n15552) );
  OA22X1 U46973 ( .A0(net263539), .A1(n41959), .B0(n41958), .B1(n40065), .Y(
        n15526) );
  CLKINVX1 U46974 ( .A(n15528), .Y(n49868) );
  OAI222XL U46975 ( .A0(net266717), .A1(n41954), .B0(n40156), .B1(n41955),
        .C0(n40307), .C1(n41956), .Y(n15528) );
  OA22X1 U46976 ( .A0(net263539), .A1(n41960), .B0(n41959), .B1(n40065), .Y(
        n15502) );
  CLKINVX1 U46977 ( .A(n15504), .Y(n49870) );
  OAI222XL U46978 ( .A0(net266717), .A1(n41955), .B0(n40156), .B1(n41956),
        .C0(n40307), .C1(n41957), .Y(n15504) );
  OAI211X1 U46979 ( .A0(n41959), .A1(n42958), .B0(n15478), .C0(n49872), .Y(
        n35332) );
  OA22X1 U46980 ( .A0(net263558), .A1(n41961), .B0(n41960), .B1(n40064), .Y(
        n15478) );
  OAI222XL U46981 ( .A0(net266717), .A1(n41956), .B0(n40156), .B1(n41957),
        .C0(n40307), .C1(n41958), .Y(n15480) );
  OAI211X1 U46982 ( .A0(n41960), .A1(n42959), .B0(n15454), .C0(n49874), .Y(
        n35324) );
  OA22X1 U46983 ( .A0(net263558), .A1(n41962), .B0(n41961), .B1(n40064), .Y(
        n15454) );
  OAI222XL U46984 ( .A0(net266717), .A1(n41957), .B0(n40156), .B1(n41958),
        .C0(n40307), .C1(n41959), .Y(n15456) );
  OAI211X1 U46985 ( .A0(n41961), .A1(n42928), .B0(n15430), .C0(n49876), .Y(
        n35316) );
  OA22X1 U46986 ( .A0(net263577), .A1(n41963), .B0(n41962), .B1(n40063), .Y(
        n15430) );
  OAI222XL U46987 ( .A0(net266717), .A1(n41958), .B0(n40156), .B1(n41959),
        .C0(n40307), .C1(n41960), .Y(n15432) );
  OAI211X1 U46988 ( .A0(n41962), .A1(n42929), .B0(n15406), .C0(n49878), .Y(
        n35308) );
  OA22X1 U46989 ( .A0(net263577), .A1(n41964), .B0(n41963), .B1(n40063), .Y(
        n15406) );
  OAI222XL U46990 ( .A0(net266717), .A1(n41959), .B0(n40156), .B1(n41960),
        .C0(n40307), .C1(n41961), .Y(n15408) );
  OAI211X1 U46991 ( .A0(n41963), .A1(n42930), .B0(n15382), .C0(n49880), .Y(
        n35300) );
  OA22X1 U46992 ( .A0(net263577), .A1(n41965), .B0(n41964), .B1(n40062), .Y(
        n15382) );
  OAI222XL U46993 ( .A0(net266717), .A1(n41960), .B0(n40156), .B1(n41961),
        .C0(n40307), .C1(n41962), .Y(n15384) );
  OAI211X1 U46994 ( .A0(n41964), .A1(n42931), .B0(n15358), .C0(n49882), .Y(
        n35292) );
  OA22X1 U46995 ( .A0(net263596), .A1(n41966), .B0(n41965), .B1(n40062), .Y(
        n15358) );
  OAI222XL U46996 ( .A0(net266717), .A1(n41961), .B0(n40155), .B1(n41962),
        .C0(n40306), .C1(n41963), .Y(n15360) );
  OAI211X1 U46997 ( .A0(n41965), .A1(n42932), .B0(n15334), .C0(n49884), .Y(
        n35284) );
  OA22X1 U46998 ( .A0(net263881), .A1(n41967), .B0(n41966), .B1(n40046), .Y(
        n15334) );
  OAI222XL U46999 ( .A0(net266717), .A1(n41962), .B0(n40155), .B1(n41963),
        .C0(n40306), .C1(n41964), .Y(n15336) );
  OAI211X1 U47000 ( .A0(n41966), .A1(n42933), .B0(n15310), .C0(n49886), .Y(
        n35276) );
  OA22X1 U47001 ( .A0(net263881), .A1(n41968), .B0(n41967), .B1(n40046), .Y(
        n15310) );
  OAI222XL U47002 ( .A0(net266738), .A1(n41963), .B0(n40155), .B1(n41964),
        .C0(n40306), .C1(n41965), .Y(n15312) );
  OAI211X1 U47003 ( .A0(n41967), .A1(n42935), .B0(n15286), .C0(n49888), .Y(
        n35268) );
  OA22X1 U47004 ( .A0(net263881), .A1(n41969), .B0(n41968), .B1(n40045), .Y(
        n15286) );
  OAI222XL U47005 ( .A0(net266738), .A1(n41964), .B0(n40155), .B1(n41965),
        .C0(n40306), .C1(n41966), .Y(n15288) );
  OAI211X1 U47006 ( .A0(n41968), .A1(n42936), .B0(n15262), .C0(n49890), .Y(
        n35260) );
  OA22X1 U47007 ( .A0(net263900), .A1(n41970), .B0(n41969), .B1(n40045), .Y(
        n15262) );
  OAI222XL U47008 ( .A0(net266738), .A1(n41965), .B0(n40155), .B1(n41966),
        .C0(n40306), .C1(n41967), .Y(n15264) );
  OAI211X1 U47009 ( .A0(n41969), .A1(n42937), .B0(n15238), .C0(n49892), .Y(
        n35252) );
  OA22X1 U47010 ( .A0(net263900), .A1(n41971), .B0(n41970), .B1(n40044), .Y(
        n15238) );
  OAI222XL U47011 ( .A0(net266738), .A1(n41966), .B0(n40155), .B1(n41967),
        .C0(n40306), .C1(n41968), .Y(n15240) );
  OAI211X1 U47012 ( .A0(n41970), .A1(n42938), .B0(n15214), .C0(n49894), .Y(
        n35244) );
  OA22X1 U47013 ( .A0(net263919), .A1(n41972), .B0(n41971), .B1(n40044), .Y(
        n15214) );
  OAI222XL U47014 ( .A0(net266738), .A1(n41967), .B0(n40155), .B1(n41968),
        .C0(n40306), .C1(n41969), .Y(n15216) );
  OAI211X1 U47015 ( .A0(n41971), .A1(n42939), .B0(n15190), .C0(n49896), .Y(
        n35236) );
  OA22X1 U47016 ( .A0(net263919), .A1(n41973), .B0(n41972), .B1(n40043), .Y(
        n15190) );
  OAI222XL U47017 ( .A0(net266738), .A1(n41968), .B0(n40155), .B1(n41969),
        .C0(n40306), .C1(n41970), .Y(n15192) );
  OAI211X1 U47018 ( .A0(n41972), .A1(n42940), .B0(n15166), .C0(n49898), .Y(
        n35228) );
  OA22X1 U47019 ( .A0(net263862), .A1(n41974), .B0(n41973), .B1(n40043), .Y(
        n15166) );
  OAI222XL U47020 ( .A0(net266738), .A1(n41969), .B0(n40155), .B1(n41970),
        .C0(n40306), .C1(n41971), .Y(n15168) );
  OAI211X1 U47021 ( .A0(n41973), .A1(n42942), .B0(n15142), .C0(n49900), .Y(
        n35220) );
  OA22X1 U47022 ( .A0(net262817), .A1(n41975), .B0(n41974), .B1(n40064), .Y(
        n15142) );
  OAI222XL U47023 ( .A0(net266738), .A1(n41970), .B0(n40154), .B1(n41971),
        .C0(n40305), .C1(n41972), .Y(n15144) );
  OAI211X1 U47024 ( .A0(n41974), .A1(n42943), .B0(n15118), .C0(n49902), .Y(
        n35212) );
  OA22X1 U47025 ( .A0(net263957), .A1(n41976), .B0(n41975), .B1(n40064), .Y(
        n15118) );
  OAI222XL U47026 ( .A0(net266738), .A1(n41971), .B0(n40154), .B1(n41972),
        .C0(n40305), .C1(n41973), .Y(n15120) );
  OAI211X1 U47027 ( .A0(n41975), .A1(n42976), .B0(n15094), .C0(n49904), .Y(
        n35204) );
  OA22X1 U47028 ( .A0(net263957), .A1(n41977), .B0(n41976), .B1(n40042), .Y(
        n15094) );
  OAI222XL U47029 ( .A0(net266759), .A1(n41972), .B0(n40154), .B1(n41973),
        .C0(n40305), .C1(n41974), .Y(n15096) );
  OAI211X1 U47030 ( .A0(n41976), .A1(n42977), .B0(n15070), .C0(n49906), .Y(
        n35196) );
  OA22X1 U47031 ( .A0(net263957), .A1(n41978), .B0(n41977), .B1(n40042), .Y(
        n15070) );
  OAI222XL U47032 ( .A0(net266759), .A1(n41973), .B0(n40154), .B1(n41974),
        .C0(n40305), .C1(n41975), .Y(n15072) );
  OAI211X1 U47033 ( .A0(n41977), .A1(n42978), .B0(n15046), .C0(n49908), .Y(
        n35188) );
  OA22X1 U47034 ( .A0(net263976), .A1(n41979), .B0(n41978), .B1(n40041), .Y(
        n15046) );
  OAI222XL U47035 ( .A0(net266759), .A1(n41974), .B0(n40154), .B1(n41975),
        .C0(n40305), .C1(n41976), .Y(n15048) );
  OAI211X1 U47036 ( .A0(n41978), .A1(n42980), .B0(n15022), .C0(n49910), .Y(
        n35180) );
  OA22X1 U47037 ( .A0(net263976), .A1(n41980), .B0(n41979), .B1(n40041), .Y(
        n15022) );
  OAI222XL U47038 ( .A0(net266759), .A1(n41975), .B0(n40154), .B1(n41976),
        .C0(n40305), .C1(n41977), .Y(n15024) );
  OAI211X1 U47039 ( .A0(n41979), .A1(n42981), .B0(n14998), .C0(n49912), .Y(
        n35172) );
  OA22X1 U47040 ( .A0(net263995), .A1(n41981), .B0(n41980), .B1(n40040), .Y(
        n14998) );
  OAI222XL U47041 ( .A0(net266759), .A1(n41976), .B0(n40154), .B1(n41977),
        .C0(n40305), .C1(n41978), .Y(n15000) );
  OAI211X1 U47042 ( .A0(n41980), .A1(n42982), .B0(n14974), .C0(n49914), .Y(
        n35164) );
  OA22X1 U47043 ( .A0(net263995), .A1(n41982), .B0(n41981), .B1(n40040), .Y(
        n14974) );
  OAI222XL U47044 ( .A0(net266759), .A1(n41977), .B0(n40154), .B1(n41978),
        .C0(n40305), .C1(n41979), .Y(n14976) );
  OAI211X1 U47045 ( .A0(n41981), .A1(n42983), .B0(n14950), .C0(n49916), .Y(
        n35156) );
  OA22X1 U47046 ( .A0(net218388), .A1(n41983), .B0(n41982), .B1(n40054), .Y(
        n14950) );
  OAI222XL U47047 ( .A0(net266759), .A1(n41978), .B0(n40153), .B1(n41979),
        .C0(n40305), .C1(n41980), .Y(n14952) );
  OAI211X1 U47048 ( .A0(n41982), .A1(n42984), .B0(n14926), .C0(n49918), .Y(
        n35148) );
  OA22X1 U47049 ( .A0(net263748), .A1(n41984), .B0(n41983), .B1(n40054), .Y(
        n14926) );
  OAI222XL U47050 ( .A0(net266759), .A1(n41979), .B0(n40153), .B1(n41980),
        .C0(n40304), .C1(n41981), .Y(n14928) );
  OAI211X1 U47051 ( .A0(n41983), .A1(n42985), .B0(n14902), .C0(n49920), .Y(
        n35140) );
  OA22X1 U47052 ( .A0(net263748), .A1(n41985), .B0(n41984), .B1(n40053), .Y(
        n14902) );
  OAI222XL U47053 ( .A0(net266759), .A1(n41980), .B0(n40153), .B1(n41981),
        .C0(n40304), .C1(n41982), .Y(n14904) );
  OAI211X1 U47054 ( .A0(n41984), .A1(n42986), .B0(n14878), .C0(n49922), .Y(
        n35132) );
  OA22X1 U47055 ( .A0(net263767), .A1(n41986), .B0(n41985), .B1(n40053), .Y(
        n14878) );
  OAI222XL U47056 ( .A0(net266759), .A1(n41981), .B0(n40153), .B1(n41982),
        .C0(n40304), .C1(n41983), .Y(n14880) );
  OAI211X1 U47057 ( .A0(n41985), .A1(n42988), .B0(n14854), .C0(n49924), .Y(
        n35124) );
  OA22X1 U47058 ( .A0(net263767), .A1(n41987), .B0(n41986), .B1(n40052), .Y(
        n14854) );
  OAI222XL U47059 ( .A0(net266759), .A1(n41982), .B0(n40153), .B1(n41983),
        .C0(n40304), .C1(n41984), .Y(n14856) );
  OAI211X1 U47060 ( .A0(n41986), .A1(n42989), .B0(n14830), .C0(n49926), .Y(
        n35116) );
  OA22X1 U47061 ( .A0(net218476), .A1(n41988), .B0(n41987), .B1(n40052), .Y(
        n14830) );
  OAI222XL U47062 ( .A0(net266780), .A1(n41983), .B0(n40153), .B1(n41984),
        .C0(n40304), .C1(n41985), .Y(n14832) );
  OAI211X1 U47063 ( .A0(n41987), .A1(n42990), .B0(n14806), .C0(n49928), .Y(
        n35108) );
  OA22X1 U47064 ( .A0(net218374), .A1(n41989), .B0(n41988), .B1(n40051), .Y(
        n14806) );
  OAI222XL U47065 ( .A0(net266780), .A1(n41984), .B0(n40153), .B1(n41985),
        .C0(n40304), .C1(n41986), .Y(n14808) );
  OAI211X1 U47066 ( .A0(n41988), .A1(n42967), .B0(n14782), .C0(n49930), .Y(
        n35100) );
  OA22X1 U47067 ( .A0(net263805), .A1(n41990), .B0(n41989), .B1(n40051), .Y(
        n14782) );
  OAI222XL U47068 ( .A0(net266780), .A1(n41985), .B0(n40153), .B1(n41986),
        .C0(n40304), .C1(n41987), .Y(n14784) );
  OAI211X1 U47069 ( .A0(n41989), .A1(n42960), .B0(n14758), .C0(n49932), .Y(
        n35092) );
  OA22X1 U47070 ( .A0(net263805), .A1(n41991), .B0(n41990), .B1(n40050), .Y(
        n14758) );
  OAI222XL U47071 ( .A0(net266780), .A1(n41986), .B0(n40153), .B1(n41987),
        .C0(n40304), .C1(n41988), .Y(n14760) );
  OAI211X1 U47072 ( .A0(n41990), .A1(n42961), .B0(n14734), .C0(n49934), .Y(
        n35084) );
  OA22X1 U47073 ( .A0(net263824), .A1(n41992), .B0(n41991), .B1(n40050), .Y(
        n14734) );
  OAI222XL U47074 ( .A0(net266780), .A1(n41987), .B0(n40152), .B1(n41988),
        .C0(n40304), .C1(n41989), .Y(n14736) );
  OAI211X1 U47075 ( .A0(n41991), .A1(n42962), .B0(n14710), .C0(n49936), .Y(
        n35076) );
  OA22X1 U47076 ( .A0(net263824), .A1(n41993), .B0(n41992), .B1(n40049), .Y(
        n14710) );
  OAI222XL U47077 ( .A0(net266780), .A1(n41988), .B0(n40152), .B1(n41989),
        .C0(n40303), .C1(n41990), .Y(n14712) );
  OAI211X1 U47078 ( .A0(n41992), .A1(n42963), .B0(n14686), .C0(n49938), .Y(
        n35068) );
  OA22X1 U47079 ( .A0(net263824), .A1(n41994), .B0(n41993), .B1(n40049), .Y(
        n14686) );
  OAI222XL U47080 ( .A0(net266780), .A1(n41989), .B0(n40152), .B1(n41990),
        .C0(n40303), .C1(n41991), .Y(n14688) );
  OAI211X1 U47081 ( .A0(n41993), .A1(n42964), .B0(n14662), .C0(n49940), .Y(
        n35060) );
  OA22X1 U47082 ( .A0(net263843), .A1(n41995), .B0(n41994), .B1(n40048), .Y(
        n14662) );
  OAI222XL U47083 ( .A0(net266780), .A1(n41990), .B0(n40152), .B1(n41991),
        .C0(n40303), .C1(n41992), .Y(n14664) );
  OAI211X1 U47084 ( .A0(n41994), .A1(n42966), .B0(n14638), .C0(n49942), .Y(
        n35052) );
  OA22X1 U47085 ( .A0(net263843), .A1(n41996), .B0(n41995), .B1(n40048), .Y(
        n14638) );
  OAI222XL U47086 ( .A0(net266780), .A1(n41991), .B0(n40152), .B1(n41992),
        .C0(n40289), .C1(n41993), .Y(n14640) );
  OAI211X1 U47087 ( .A0(n41995), .A1(n42967), .B0(n14614), .C0(n49944), .Y(
        n35044) );
  OA22X1 U47088 ( .A0(net263862), .A1(n41997), .B0(n41996), .B1(n40047), .Y(
        n14614) );
  OAI222XL U47089 ( .A0(net266780), .A1(n41992), .B0(n40152), .B1(n41993),
        .C0(n40288), .C1(n41994), .Y(n14616) );
  OAI211X1 U47090 ( .A0(n41996), .A1(n42968), .B0(n14590), .C0(n49946), .Y(
        n35036) );
  OA22X1 U47091 ( .A0(net263862), .A1(n41998), .B0(n41997), .B1(n40047), .Y(
        n14590) );
  OAI222XL U47092 ( .A0(net221954), .A1(n41993), .B0(n40152), .B1(n41994),
        .C0(n40288), .C1(n41995), .Y(n14592) );
  OAI211X1 U47093 ( .A0(n41997), .A1(n42969), .B0(n14566), .C0(n49948), .Y(
        n35028) );
  OA22X1 U47094 ( .A0(net263064), .A1(n41999), .B0(n41998), .B1(n40092), .Y(
        n14566) );
  OAI222XL U47095 ( .A0(net266780), .A1(n41994), .B0(n40152), .B1(n41995),
        .C0(n40288), .C1(n41996), .Y(n14568) );
  OAI211X1 U47096 ( .A0(n41998), .A1(n42970), .B0(n14542), .C0(n49950), .Y(
        n35020) );
  OA22X1 U47097 ( .A0(net263064), .A1(n42000), .B0(n41999), .B1(n40092), .Y(
        n14542) );
  CLKINVX1 U47098 ( .A(n14544), .Y(n49950) );
  OAI222XL U47099 ( .A0(net266780), .A1(n41995), .B0(net218220), .B1(n41996),
        .C0(n40288), .C1(n41997), .Y(n14544) );
  OAI211X1 U47100 ( .A0(n41999), .A1(n42971), .B0(n14518), .C0(n49952), .Y(
        n35012) );
  OA22X1 U47101 ( .A0(net263083), .A1(n42001), .B0(n42000), .B1(n40091), .Y(
        n14518) );
  OAI222XL U47102 ( .A0(net266528), .A1(n41996), .B0(n40167), .B1(n41997),
        .C0(n40288), .C1(n41998), .Y(n14520) );
  OAI211X1 U47103 ( .A0(n42000), .A1(n42973), .B0(n14494), .C0(n49954), .Y(
        n35004) );
  OA22X1 U47104 ( .A0(net263083), .A1(n42002), .B0(n42001), .B1(n40091), .Y(
        n14494) );
  OAI222XL U47105 ( .A0(net266528), .A1(n41997), .B0(n40167), .B1(n41998),
        .C0(n40288), .C1(n41999), .Y(n14496) );
  OAI211X1 U47106 ( .A0(n42001), .A1(n42974), .B0(n14470), .C0(n49956), .Y(
        n34996) );
  OA22X1 U47107 ( .A0(net263102), .A1(n42003), .B0(n42002), .B1(n40090), .Y(
        n14470) );
  OAI222XL U47108 ( .A0(net266528), .A1(n41998), .B0(n40166), .B1(n41999),
        .C0(n40288), .C1(n42000), .Y(n14472) );
  OAI211X1 U47109 ( .A0(n42002), .A1(n42975), .B0(n14446), .C0(n49958), .Y(
        n34988) );
  OA22X1 U47110 ( .A0(net263102), .A1(n42004), .B0(n42003), .B1(n40090), .Y(
        n14446) );
  OAI222XL U47111 ( .A0(net266528), .A1(n41999), .B0(n40166), .B1(n42000),
        .C0(n40288), .C1(n42001), .Y(n14448) );
  OAI211X1 U47112 ( .A0(n42003), .A1(n42895), .B0(n14422), .C0(n49960), .Y(
        n34980) );
  OA22X1 U47113 ( .A0(net263121), .A1(n42005), .B0(n42004), .B1(n40089), .Y(
        n14422) );
  OAI222XL U47114 ( .A0(net266528), .A1(n42000), .B0(n40166), .B1(n42001),
        .C0(n40288), .C1(n42002), .Y(n14424) );
  OAI211X1 U47115 ( .A0(n42004), .A1(n42880), .B0(n14398), .C0(n49962), .Y(
        n34972) );
  OA22X1 U47116 ( .A0(net263121), .A1(n42006), .B0(n42005), .B1(n40089), .Y(
        n14398) );
  OAI222XL U47117 ( .A0(net266528), .A1(n42001), .B0(n40166), .B1(n42002),
        .C0(n40287), .C1(n42003), .Y(n14400) );
  OAI211X1 U47118 ( .A0(n42005), .A1(n42881), .B0(n14374), .C0(n49964), .Y(
        n34964) );
  OA22X1 U47119 ( .A0(net263121), .A1(n42007), .B0(n42006), .B1(n40088), .Y(
        n14374) );
  OAI222XL U47120 ( .A0(net266528), .A1(n42002), .B0(n40166), .B1(n42003),
        .C0(n40287), .C1(n42004), .Y(n14376) );
  OAI211X1 U47121 ( .A0(n42006), .A1(n42882), .B0(n14350), .C0(n49966), .Y(
        n34956) );
  OA22X1 U47122 ( .A0(net263140), .A1(n42008), .B0(n42007), .B1(n40088), .Y(
        n14350) );
  OAI222XL U47123 ( .A0(net266528), .A1(n42003), .B0(n40166), .B1(n42004),
        .C0(n40287), .C1(n42005), .Y(n14352) );
  OAI211X1 U47124 ( .A0(n42007), .A1(n42883), .B0(n14326), .C0(n49968), .Y(
        n34948) );
  OA22X1 U47125 ( .A0(net263140), .A1(n42009), .B0(n42008), .B1(n40087), .Y(
        n14326) );
  OAI222XL U47126 ( .A0(net266549), .A1(n42004), .B0(n40166), .B1(n42005),
        .C0(n40287), .C1(n42006), .Y(n14328) );
  OAI211X1 U47127 ( .A0(n42008), .A1(n42885), .B0(n14302), .C0(n49970), .Y(
        n34940) );
  OA22X1 U47128 ( .A0(net263159), .A1(n42010), .B0(n42009), .B1(n40087), .Y(
        n14302) );
  OAI222XL U47129 ( .A0(net266549), .A1(n42005), .B0(n40166), .B1(n42006),
        .C0(n40287), .C1(n42007), .Y(n14304) );
  OAI211X1 U47130 ( .A0(n42009), .A1(n42886), .B0(n14278), .C0(n49972), .Y(
        n34932) );
  OA22X1 U47131 ( .A0(net263159), .A1(n42011), .B0(n42010), .B1(n40086), .Y(
        n14278) );
  OAI222XL U47132 ( .A0(net266549), .A1(n42006), .B0(n40166), .B1(n42007),
        .C0(n40287), .C1(n42008), .Y(n14280) );
  OAI211X1 U47133 ( .A0(n42010), .A1(n42887), .B0(n14254), .C0(n49974), .Y(
        n34924) );
  OA22X1 U47134 ( .A0(net263178), .A1(n42012), .B0(n42011), .B1(n40086), .Y(
        n14254) );
  OAI222XL U47135 ( .A0(net266549), .A1(n42007), .B0(n40165), .B1(n42008),
        .C0(n40287), .C1(n42009), .Y(n14256) );
  OAI211X1 U47136 ( .A0(n42011), .A1(n42888), .B0(n14230), .C0(n49976), .Y(
        n34916) );
  OA22X1 U47137 ( .A0(net263178), .A1(n42013), .B0(n42012), .B1(n40085), .Y(
        n14230) );
  OAI222XL U47138 ( .A0(net266549), .A1(n42008), .B0(n40165), .B1(n42009),
        .C0(n40287), .C1(n42010), .Y(n14232) );
  OAI211X1 U47139 ( .A0(n42012), .A1(n42889), .B0(n14206), .C0(n49978), .Y(
        n34908) );
  OA22X1 U47140 ( .A0(net218556), .A1(n42014), .B0(n42013), .B1(n40085), .Y(
        n14206) );
  OAI222XL U47141 ( .A0(net266549), .A1(n42009), .B0(n40165), .B1(n42010),
        .C0(n40286), .C1(n42011), .Y(n14208) );
  OAI211X1 U47142 ( .A0(n42013), .A1(n42890), .B0(n14182), .C0(n49980), .Y(
        n34900) );
  OA22X1 U47143 ( .A0(net262931), .A1(n42015), .B0(n42014), .B1(n40100), .Y(
        n14182) );
  OAI222XL U47144 ( .A0(net266549), .A1(n42010), .B0(n40165), .B1(n42011),
        .C0(n40286), .C1(n42012), .Y(n14184) );
  OAI211X1 U47145 ( .A0(n42014), .A1(n42892), .B0(n14158), .C0(n49982), .Y(
        n34892) );
  OA22X1 U47146 ( .A0(net262931), .A1(n42016), .B0(n42015), .B1(n40100), .Y(
        n14158) );
  OAI222XL U47147 ( .A0(net266549), .A1(n42011), .B0(n40165), .B1(n42012),
        .C0(n40287), .C1(n42013), .Y(n14160) );
  OAI211X1 U47148 ( .A0(n42015), .A1(n42893), .B0(n14134), .C0(n49984), .Y(
        n34884) );
  OA22X1 U47149 ( .A0(net262950), .A1(n42017), .B0(n42016), .B1(n40099), .Y(
        n14134) );
  OAI222XL U47150 ( .A0(net266549), .A1(n42012), .B0(n40165), .B1(n42013),
        .C0(n40286), .C1(n42014), .Y(n14136) );
  OAI211X1 U47151 ( .A0(n42016), .A1(n42894), .B0(n14110), .C0(n49986), .Y(
        n34876) );
  OA22X1 U47152 ( .A0(net262950), .A1(n42018), .B0(n42017), .B1(n40099), .Y(
        n14110) );
  OAI222XL U47153 ( .A0(net266549), .A1(n42013), .B0(n40165), .B1(n42014),
        .C0(n40286), .C1(n42015), .Y(n14112) );
  OAI211X1 U47154 ( .A0(n42017), .A1(n42895), .B0(n14086), .C0(n49988), .Y(
        n34868) );
  OA22X1 U47155 ( .A0(net262969), .A1(n42019), .B0(n42018), .B1(n40098), .Y(
        n14086) );
  OAI222XL U47156 ( .A0(net266570), .A1(n42014), .B0(n40165), .B1(n42015),
        .C0(n40286), .C1(n42016), .Y(n14088) );
  OAI211X1 U47157 ( .A0(n42018), .A1(n42864), .B0(n14062), .C0(n49990), .Y(
        n34860) );
  OA22X1 U47158 ( .A0(net262969), .A1(n42020), .B0(n42019), .B1(n40098), .Y(
        n14062) );
  OAI222XL U47159 ( .A0(net266570), .A1(n42015), .B0(n40164), .B1(n42016),
        .C0(n40286), .C1(n42017), .Y(n14064) );
  OAI211X1 U47160 ( .A0(n42019), .A1(n42865), .B0(n14038), .C0(n49992), .Y(
        n34852) );
  OA22X1 U47161 ( .A0(net262969), .A1(n42021), .B0(n42020), .B1(n40097), .Y(
        n14038) );
  OAI222XL U47162 ( .A0(net266570), .A1(n42016), .B0(n40164), .B1(n42017),
        .C0(n40286), .C1(n42018), .Y(n14040) );
  OAI211X1 U47163 ( .A0(n42020), .A1(n42866), .B0(n14014), .C0(n49994), .Y(
        n34844) );
  OA22X1 U47164 ( .A0(net262988), .A1(n42022), .B0(n42021), .B1(n40097), .Y(
        n14014) );
  OAI222XL U47165 ( .A0(net266570), .A1(n42017), .B0(n40164), .B1(n42018),
        .C0(n40286), .C1(n42019), .Y(n14016) );
  OAI211X1 U47166 ( .A0(n42021), .A1(n42867), .B0(n13990), .C0(n49996), .Y(
        n34836) );
  OA22X1 U47167 ( .A0(net262988), .A1(n42023), .B0(n42022), .B1(n40096), .Y(
        n13990) );
  OAI222XL U47168 ( .A0(net266570), .A1(n42018), .B0(n40164), .B1(n42019),
        .C0(net217178), .C1(n42020), .Y(n13992) );
  OAI211X1 U47169 ( .A0(n42022), .A1(n42869), .B0(n13966), .C0(n49998), .Y(
        n34828) );
  OA22X1 U47170 ( .A0(net263007), .A1(n42024), .B0(n42023), .B1(n40096), .Y(
        n13966) );
  OAI222XL U47171 ( .A0(net266570), .A1(n42019), .B0(n40164), .B1(n42020),
        .C0(net217178), .C1(n42021), .Y(n13968) );
  OAI211X1 U47172 ( .A0(n42023), .A1(n42870), .B0(n13942), .C0(n50000), .Y(
        n34820) );
  OA22X1 U47173 ( .A0(net263007), .A1(n42025), .B0(n42024), .B1(n40095), .Y(
        n13942) );
  OAI222XL U47174 ( .A0(net266570), .A1(n42020), .B0(n40164), .B1(n42021),
        .C0(net217178), .C1(n42022), .Y(n13944) );
  OAI211X1 U47175 ( .A0(n42024), .A1(n42871), .B0(n13918), .C0(n50002), .Y(
        n34812) );
  OA22X1 U47176 ( .A0(net263026), .A1(n42026), .B0(n42025), .B1(n40095), .Y(
        n13918) );
  OAI222XL U47177 ( .A0(net266570), .A1(n42021), .B0(n40164), .B1(n42022),
        .C0(net217178), .C1(n42023), .Y(n13920) );
  OAI211X1 U47178 ( .A0(n42025), .A1(n42872), .B0(n13894), .C0(n50004), .Y(
        n34804) );
  OA22X1 U47179 ( .A0(net263026), .A1(n42027), .B0(n42026), .B1(n40094), .Y(
        n13894) );
  OAI222XL U47180 ( .A0(net266570), .A1(n42022), .B0(n40164), .B1(n42023),
        .C0(net217178), .C1(n42024), .Y(n13896) );
  OAI211X1 U47181 ( .A0(n42026), .A1(n42873), .B0(n13870), .C0(n50006), .Y(
        n34796) );
  OA22X1 U47182 ( .A0(net263045), .A1(n42028), .B0(n42027), .B1(n40094), .Y(
        n13870) );
  OAI222XL U47183 ( .A0(net266570), .A1(n42023), .B0(n40164), .B1(n42024),
        .C0(net217178), .C1(n42025), .Y(n13872) );
  OAI211X1 U47184 ( .A0(n42027), .A1(n42874), .B0(n13846), .C0(n50008), .Y(
        n34788) );
  OA22X1 U47185 ( .A0(net263045), .A1(n42029), .B0(n42028), .B1(n40093), .Y(
        n13846) );
  OAI222XL U47186 ( .A0(net266591), .A1(n42024), .B0(n40163), .B1(n42025),
        .C0(net217178), .C1(n42026), .Y(n13848) );
  OAI211X1 U47187 ( .A0(n42028), .A1(n42876), .B0(n13822), .C0(n50010), .Y(
        n34780) );
  OA22X1 U47188 ( .A0(net263064), .A1(n42030), .B0(n42029), .B1(n40093), .Y(
        n13822) );
  OAI222XL U47189 ( .A0(net266591), .A1(n42025), .B0(n40163), .B1(n42026),
        .C0(net217178), .C1(n42027), .Y(n13824) );
  OAI211X1 U47190 ( .A0(n42029), .A1(n42877), .B0(n13798), .C0(n50012), .Y(
        n34772) );
  OA22X1 U47191 ( .A0(net263330), .A1(n42031), .B0(n42030), .B1(n40077), .Y(
        n13798) );
  OAI222XL U47192 ( .A0(net266591), .A1(n42026), .B0(n40163), .B1(n42027),
        .C0(n40289), .C1(n42028), .Y(n13800) );
  OAI211X1 U47193 ( .A0(n42030), .A1(n42878), .B0(n13774), .C0(n50014), .Y(
        n34764) );
  OA22X1 U47194 ( .A0(net263349), .A1(n42032), .B0(n42031), .B1(n40077), .Y(
        n13774) );
  OAI222XL U47195 ( .A0(net266591), .A1(n42027), .B0(n40163), .B1(n42028),
        .C0(n40289), .C1(n42029), .Y(n13776) );
  OAI211X1 U47196 ( .A0(n42031), .A1(n42879), .B0(n13750), .C0(n50016), .Y(
        n34756) );
  OA22X1 U47197 ( .A0(net263349), .A1(n42033), .B0(n42032), .B1(n40076), .Y(
        n13750) );
  OAI222XL U47198 ( .A0(net266654), .A1(n42028), .B0(n40163), .B1(n42029),
        .C0(n40289), .C1(n42030), .Y(n13752) );
  OAI211X1 U47199 ( .A0(n42032), .A1(n42912), .B0(n13726), .C0(n50018), .Y(
        n34748) );
  OA22X1 U47200 ( .A0(net263349), .A1(n42034), .B0(n42033), .B1(n40076), .Y(
        n13726) );
  OAI222XL U47201 ( .A0(net266591), .A1(n42029), .B0(n40159), .B1(n42030),
        .C0(n40289), .C1(n42031), .Y(n13728) );
  OAI211X1 U47202 ( .A0(n42033), .A1(n42913), .B0(n13702), .C0(n50020), .Y(
        n34740) );
  OA22X1 U47203 ( .A0(net263368), .A1(n42035), .B0(n42034), .B1(n40075), .Y(
        n13702) );
  OAI222XL U47204 ( .A0(net266591), .A1(n42030), .B0(n40163), .B1(n42031),
        .C0(n40289), .C1(n42032), .Y(n13704) );
  OAI211X1 U47205 ( .A0(n42034), .A1(n42914), .B0(n13678), .C0(n50022), .Y(
        n34732) );
  OA22X1 U47206 ( .A0(net263368), .A1(n42036), .B0(n42035), .B1(n40075), .Y(
        n13678) );
  OAI222XL U47207 ( .A0(net266591), .A1(n42031), .B0(n40163), .B1(n42032),
        .C0(n40289), .C1(n42033), .Y(n13680) );
  OAI211X1 U47208 ( .A0(n42035), .A1(n42916), .B0(n13654), .C0(n50024), .Y(
        n34724) );
  OA22X1 U47209 ( .A0(net263387), .A1(n42037), .B0(n42036), .B1(n40074), .Y(
        n13654) );
  OAI222XL U47210 ( .A0(net266591), .A1(n42032), .B0(n40162), .B1(n42033),
        .C0(n40289), .C1(n42034), .Y(n13656) );
  OAI211X1 U47211 ( .A0(n42036), .A1(n42917), .B0(n13630), .C0(n50026), .Y(
        n34716) );
  OA22X1 U47212 ( .A0(net263387), .A1(n42038), .B0(n42037), .B1(n40074), .Y(
        n13630) );
  OAI222XL U47213 ( .A0(net266591), .A1(n42033), .B0(n40162), .B1(n42034),
        .C0(n40289), .C1(n42035), .Y(n13632) );
  OAI211X1 U47214 ( .A0(n42037), .A1(n42918), .B0(n13606), .C0(n50028), .Y(
        n34708) );
  OA22X1 U47215 ( .A0(net263406), .A1(n42039), .B0(n42038), .B1(n40073), .Y(
        n13606) );
  OAI222XL U47216 ( .A0(net266612), .A1(n42034), .B0(n40162), .B1(n42035),
        .C0(n40289), .C1(n42036), .Y(n13608) );
  OAI211X1 U47217 ( .A0(n42038), .A1(n42919), .B0(n13582), .C0(n50030), .Y(
        n34700) );
  OA22X1 U47218 ( .A0(net263406), .A1(n42040), .B0(n42039), .B1(n40073), .Y(
        n13582) );
  OAI222XL U47219 ( .A0(net266612), .A1(n42035), .B0(n40162), .B1(n42036),
        .C0(n40290), .C1(n42037), .Y(n13584) );
  OAI211X1 U47220 ( .A0(n42039), .A1(n42920), .B0(n13558), .C0(n50032), .Y(
        n34692) );
  OA22X1 U47221 ( .A0(net218412), .A1(n42041), .B0(n42040), .B1(n40072), .Y(
        n13558) );
  OAI222XL U47222 ( .A0(net266612), .A1(n42036), .B0(n40162), .B1(n42037),
        .C0(n40290), .C1(n42038), .Y(n13560) );
  OAI211X1 U47223 ( .A0(n42040), .A1(n42921), .B0(n13534), .C0(n50034), .Y(
        n34684) );
  OA22X1 U47224 ( .A0(net218488), .A1(n42042), .B0(n42041), .B1(n40072), .Y(
        n13534) );
  OAI222XL U47225 ( .A0(net266612), .A1(n42037), .B0(n40162), .B1(n42038),
        .C0(n40290), .C1(n42039), .Y(n13536) );
  OAI211X1 U47226 ( .A0(n42041), .A1(n42923), .B0(n13510), .C0(n50036), .Y(
        n34676) );
  OA22X1 U47227 ( .A0(net263444), .A1(n42043), .B0(n42042), .B1(n40071), .Y(
        n13510) );
  OAI222XL U47228 ( .A0(net266612), .A1(n42038), .B0(n40162), .B1(n42039),
        .C0(n40290), .C1(n42040), .Y(n13512) );
  OAI211X1 U47229 ( .A0(n42042), .A1(n42924), .B0(n13486), .C0(n50038), .Y(
        n34668) );
  OA22X1 U47230 ( .A0(net263444), .A1(n42044), .B0(n42043), .B1(n40071), .Y(
        n13486) );
  OAI222XL U47231 ( .A0(net266612), .A1(n42039), .B0(n40162), .B1(n42040),
        .C0(n40290), .C1(n42041), .Y(n13488) );
  OAI211X1 U47232 ( .A0(n42043), .A1(n42925), .B0(n13462), .C0(n50040), .Y(
        n34660) );
  OA22X1 U47233 ( .A0(net263444), .A1(n42045), .B0(n42044), .B1(n40070), .Y(
        n13462) );
  OAI222XL U47234 ( .A0(net266612), .A1(n42040), .B0(n40162), .B1(n42041),
        .C0(n40290), .C1(n42042), .Y(n13464) );
  OAI211X1 U47235 ( .A0(n42044), .A1(n42926), .B0(n13438), .C0(n50042), .Y(
        n34652) );
  OA22X1 U47236 ( .A0(net263463), .A1(n42046), .B0(n42045), .B1(n40070), .Y(
        n13438) );
  OAI222XL U47237 ( .A0(net266612), .A1(n42041), .B0(n40161), .B1(n42042),
        .C0(n40290), .C1(n42043), .Y(n13440) );
  OAI211X1 U47238 ( .A0(n42045), .A1(n42927), .B0(n13414), .C0(n50044), .Y(
        n34644) );
  OA22X1 U47239 ( .A0(net218414), .A1(n42047), .B0(n42046), .B1(n40084), .Y(
        n13414) );
  OAI222XL U47240 ( .A0(net266612), .A1(n42042), .B0(n40161), .B1(n42043),
        .C0(n40290), .C1(n42044), .Y(n13416) );
  OAI211X1 U47241 ( .A0(n42046), .A1(n42896), .B0(n13390), .C0(n50046), .Y(
        n34636) );
  OA22X1 U47242 ( .A0(net263216), .A1(n42048), .B0(n42047), .B1(n40084), .Y(
        n13390) );
  OAI222XL U47243 ( .A0(net266612), .A1(n42043), .B0(n40161), .B1(n42044),
        .C0(n40290), .C1(n42045), .Y(n13392) );
  OAI211X1 U47244 ( .A0(n42047), .A1(n42897), .B0(n13366), .C0(n50048), .Y(
        n34628) );
  OA22X1 U47245 ( .A0(net263216), .A1(n42049), .B0(n42048), .B1(n40083), .Y(
        n13366) );
  OAI222XL U47246 ( .A0(net266633), .A1(n42044), .B0(n40161), .B1(n42045),
        .C0(n40291), .C1(n42046), .Y(n13368) );
  OAI211X1 U47247 ( .A0(n42048), .A1(n42898), .B0(n13342), .C0(n50050), .Y(
        n34620) );
  OA22X1 U47248 ( .A0(net263216), .A1(n42050), .B0(n42049), .B1(n40083), .Y(
        n13342) );
  OAI222XL U47249 ( .A0(net266633), .A1(n42045), .B0(n40161), .B1(n42046),
        .C0(n40291), .C1(n42047), .Y(n13344) );
  OAI211X1 U47250 ( .A0(n42049), .A1(n42899), .B0(n13318), .C0(n50052), .Y(
        n34612) );
  OA22X1 U47251 ( .A0(net263235), .A1(n42051), .B0(n42050), .B1(n40082), .Y(
        n13318) );
  OAI222XL U47252 ( .A0(net266633), .A1(n42046), .B0(n40161), .B1(n42047),
        .C0(n40291), .C1(n42048), .Y(n13320) );
  OAI211X1 U47253 ( .A0(n42050), .A1(n42901), .B0(n13294), .C0(n50054), .Y(
        n34604) );
  OA22X1 U47254 ( .A0(net263235), .A1(n42052), .B0(n42051), .B1(n40082), .Y(
        n13294) );
  OAI222XL U47255 ( .A0(net266633), .A1(n42047), .B0(n40161), .B1(n42048),
        .C0(n40291), .C1(n42049), .Y(n13296) );
  OAI211X1 U47256 ( .A0(n42051), .A1(n42902), .B0(n13270), .C0(n50056), .Y(
        n34596) );
  OA22X1 U47257 ( .A0(net263254), .A1(n42053), .B0(n42052), .B1(n40081), .Y(
        n13270) );
  OAI222XL U47258 ( .A0(net266633), .A1(n42048), .B0(n40161), .B1(n42049),
        .C0(n40291), .C1(n42050), .Y(n13272) );
  OAI211X1 U47259 ( .A0(n42052), .A1(n42903), .B0(n13246), .C0(n50058), .Y(
        n34588) );
  OA22X1 U47260 ( .A0(net263254), .A1(n42054), .B0(n42053), .B1(n40081), .Y(
        n13246) );
  OAI222XL U47261 ( .A0(net266633), .A1(n42049), .B0(n40160), .B1(n42050),
        .C0(n40291), .C1(n42051), .Y(n13248) );
  OAI211X1 U47262 ( .A0(n42053), .A1(n42904), .B0(n13222), .C0(n50060), .Y(
        n34580) );
  OA22X1 U47263 ( .A0(net218300), .A1(n42055), .B0(n42054), .B1(n40080), .Y(
        n13222) );
  OAI222XL U47264 ( .A0(net266633), .A1(n42050), .B0(n40160), .B1(n42051),
        .C0(n40291), .C1(n42052), .Y(n13224) );
  OAI211X1 U47265 ( .A0(n42054), .A1(n42905), .B0(n13198), .C0(n50062), .Y(
        n34572) );
  OA22X1 U47266 ( .A0(net218314), .A1(n42056), .B0(n42055), .B1(n40080), .Y(
        n13198) );
  OAI222XL U47267 ( .A0(net266633), .A1(n42051), .B0(n40160), .B1(n42052),
        .C0(n40291), .C1(n42053), .Y(n13200) );
  OAI211X1 U47268 ( .A0(n42055), .A1(n42906), .B0(n13174), .C0(n50064), .Y(
        n34564) );
  OA22X1 U47269 ( .A0(net263292), .A1(n36897), .B0(n42056), .B1(n40079), .Y(
        n13174) );
  OAI211X1 U47270 ( .A0(n42056), .A1(n42908), .B0(n13150), .C0(n50066), .Y(
        n34556) );
  OAI222XL U47271 ( .A0(net266633), .A1(n42053), .B0(n40160), .B1(n42054),
        .C0(n40292), .C1(n42055), .Y(n13152) );
  OAI222XL U47272 ( .A0(net266654), .A1(n42054), .B0(n40160), .B1(n42055),
        .C0(n40292), .C1(n42056), .Y(n13128) );
  OAI222XL U47273 ( .A0(net266654), .A1(n42055), .B0(n40160), .B1(n42056),
        .C0(n40292), .C1(n36892), .Y(n13104) );
  OAI222XL U47274 ( .A0(net266654), .A1(n42056), .B0(n40160), .B1(n36891),
        .C0(n40292), .C1(n42609), .Y(n13078) );
  AOI222XL U47275 ( .A0(net265644), .A1(n50585), .B0(n40214), .B1(n50584),
        .C0(net216978), .C1(n50583), .Y(n13130) );
  AOI222XL U47276 ( .A0(net265720), .A1(n50382), .B0(n40266), .B1(n50381),
        .C0(net216978), .C1(n50380), .Y(n13109) );
  AOI222XL U47277 ( .A0(net265644), .A1(n50167), .B0(n40203), .B1(n50166),
        .C0(net216970), .C1(n50165), .Y(n13112) );
  OA22X1 U47278 ( .A0(net262551), .A1(n42069), .B0(n42068), .B1(n40063), .Y(
        n19090) );
  CLKINVX1 U47279 ( .A(n19092), .Y(n49571) );
  OAI222XL U47280 ( .A0(net266402), .A1(n42064), .B0(n40174), .B1(n42065),
        .C0(n40303), .C1(n42066), .Y(n19092) );
  OA22X1 U47281 ( .A0(net262551), .A1(n42070), .B0(n42069), .B1(n40117), .Y(
        n19066) );
  CLKINVX1 U47282 ( .A(n19068), .Y(n49573) );
  OAI222XL U47283 ( .A0(net266402), .A1(n42065), .B0(n40174), .B1(n42066),
        .C0(n40302), .C1(n42067), .Y(n19068) );
  OA22X1 U47284 ( .A0(net262570), .A1(n42071), .B0(n42070), .B1(n40117), .Y(
        n19042) );
  CLKINVX1 U47285 ( .A(n19044), .Y(n49575) );
  OAI222XL U47286 ( .A0(net266402), .A1(n42066), .B0(n40174), .B1(n42067),
        .C0(n40302), .C1(n42068), .Y(n19044) );
  OA22X1 U47287 ( .A0(net262570), .A1(n42072), .B0(n42071), .B1(n40116), .Y(
        n19018) );
  CLKINVX1 U47288 ( .A(n19020), .Y(n49577) );
  OAI222XL U47289 ( .A0(net266402), .A1(n42067), .B0(n40173), .B1(n42068),
        .C0(n40302), .C1(n42069), .Y(n19020) );
  OA22X1 U47290 ( .A0(net262589), .A1(n42073), .B0(n42072), .B1(n40116), .Y(
        n18994) );
  CLKINVX1 U47291 ( .A(n18996), .Y(n49579) );
  OAI222XL U47292 ( .A0(net266402), .A1(n42068), .B0(n40173), .B1(n42069),
        .C0(n40302), .C1(n42070), .Y(n18996) );
  OA22X1 U47293 ( .A0(net262589), .A1(n42074), .B0(n42073), .B1(n40115), .Y(
        n18970) );
  CLKINVX1 U47294 ( .A(n18972), .Y(n49581) );
  OAI222XL U47295 ( .A0(net266402), .A1(n42069), .B0(n40173), .B1(n42070),
        .C0(n40302), .C1(n42071), .Y(n18972) );
  OA22X1 U47296 ( .A0(net262608), .A1(n42075), .B0(n42074), .B1(n40115), .Y(
        n18946) );
  CLKINVX1 U47297 ( .A(n18948), .Y(n49583) );
  OAI222XL U47298 ( .A0(net266402), .A1(n42070), .B0(n40173), .B1(n42071),
        .C0(n40302), .C1(n42072), .Y(n18948) );
  OA22X1 U47299 ( .A0(net262608), .A1(n42076), .B0(n42075), .B1(n40114), .Y(
        n18922) );
  CLKINVX1 U47300 ( .A(n18924), .Y(n49585) );
  OAI222XL U47301 ( .A0(net266402), .A1(n42071), .B0(n40173), .B1(n42072),
        .C0(n40302), .C1(n42073), .Y(n18924) );
  OA22X1 U47302 ( .A0(net262608), .A1(n42077), .B0(n42076), .B1(n40114), .Y(
        n18898) );
  CLKINVX1 U47303 ( .A(n18900), .Y(n49587) );
  OAI222XL U47304 ( .A0(net266423), .A1(n42072), .B0(n40173), .B1(n42073),
        .C0(n40302), .C1(n42074), .Y(n18900) );
  OA22X1 U47305 ( .A0(net262627), .A1(n42078), .B0(n42077), .B1(n40113), .Y(
        n18874) );
  CLKINVX1 U47306 ( .A(n18876), .Y(n49589) );
  OAI222XL U47307 ( .A0(net266423), .A1(n42073), .B0(n40173), .B1(n42074),
        .C0(n40302), .C1(n42075), .Y(n18876) );
  OA22X1 U47308 ( .A0(net262627), .A1(n42079), .B0(n42078), .B1(n40113), .Y(
        n18850) );
  CLKINVX1 U47309 ( .A(n18852), .Y(n49591) );
  OAI222XL U47310 ( .A0(net266423), .A1(n42074), .B0(n40173), .B1(n42075),
        .C0(n40301), .C1(n42076), .Y(n18852) );
  OA22X1 U47311 ( .A0(net262646), .A1(n42080), .B0(n42079), .B1(n40112), .Y(
        n18826) );
  CLKINVX1 U47312 ( .A(n18828), .Y(n49593) );
  OAI222XL U47313 ( .A0(net266423), .A1(n42075), .B0(n40173), .B1(n42076),
        .C0(n40301), .C1(n42077), .Y(n18828) );
  OA22X1 U47314 ( .A0(net262646), .A1(n42081), .B0(n42080), .B1(n40112), .Y(
        n18802) );
  CLKINVX1 U47315 ( .A(n18804), .Y(n49595) );
  OAI222XL U47316 ( .A0(net266423), .A1(n42076), .B0(n40172), .B1(n42077),
        .C0(n40301), .C1(n42078), .Y(n18804) );
  OA22X1 U47317 ( .A0(net262380), .A1(n42082), .B0(n42081), .B1(n40123), .Y(
        n18778) );
  CLKINVX1 U47318 ( .A(n18780), .Y(n49597) );
  OAI222XL U47319 ( .A0(net266423), .A1(n42077), .B0(n40172), .B1(n42078),
        .C0(n40301), .C1(n42079), .Y(n18780) );
  OA22X1 U47320 ( .A0(net262399), .A1(n42083), .B0(n42082), .B1(n40123), .Y(
        n18754) );
  CLKINVX1 U47321 ( .A(n18756), .Y(n49599) );
  OAI222XL U47322 ( .A0(net266423), .A1(n42078), .B0(n40172), .B1(n42079),
        .C0(n40301), .C1(n42080), .Y(n18756) );
  OA22X1 U47323 ( .A0(net262399), .A1(n42084), .B0(n42083), .B1(n40122), .Y(
        n18730) );
  CLKINVX1 U47324 ( .A(n18732), .Y(n49601) );
  OAI222XL U47325 ( .A0(net266423), .A1(n42079), .B0(n40172), .B1(n42080),
        .C0(n40301), .C1(n42081), .Y(n18732) );
  OA22X1 U47326 ( .A0(net262418), .A1(n42085), .B0(n42084), .B1(n40122), .Y(
        n18706) );
  CLKINVX1 U47327 ( .A(n18708), .Y(n49603) );
  OAI222XL U47328 ( .A0(net266423), .A1(n42080), .B0(n40172), .B1(n42081),
        .C0(n40301), .C1(n42082), .Y(n18708) );
  OA22X1 U47329 ( .A0(net262418), .A1(n42086), .B0(n42085), .B1(n40121), .Y(
        n18682) );
  CLKINVX1 U47330 ( .A(n18684), .Y(n49605) );
  OAI222XL U47331 ( .A0(net266423), .A1(n42081), .B0(n40172), .B1(n42082),
        .C0(n40301), .C1(n42083), .Y(n18684) );
  OA22X1 U47332 ( .A0(net262437), .A1(n42087), .B0(n42086), .B1(n40121), .Y(
        n18658) );
  CLKINVX1 U47333 ( .A(n18660), .Y(n49607) );
  OAI222XL U47334 ( .A0(net266444), .A1(n42082), .B0(n40172), .B1(n42083),
        .C0(n40301), .C1(n42084), .Y(n18660) );
  OA22X1 U47335 ( .A0(net262437), .A1(n42088), .B0(n42087), .B1(n40120), .Y(
        n18634) );
  CLKINVX1 U47336 ( .A(n18636), .Y(n49609) );
  OAI222XL U47337 ( .A0(net266444), .A1(n42083), .B0(n40172), .B1(n42084),
        .C0(n40300), .C1(n42085), .Y(n18636) );
  OA22X1 U47338 ( .A0(net262456), .A1(n42089), .B0(n42088), .B1(n40120), .Y(
        n18610) );
  CLKINVX1 U47339 ( .A(n18612), .Y(n49611) );
  OAI222XL U47340 ( .A0(net266444), .A1(n42084), .B0(n40171), .B1(n42085),
        .C0(n40300), .C1(n42086), .Y(n18612) );
  OA22X1 U47341 ( .A0(net262456), .A1(n42090), .B0(n42089), .B1(net218940),
        .Y(n18586) );
  CLKINVX1 U47342 ( .A(n18588), .Y(n49613) );
  OAI222XL U47343 ( .A0(net266444), .A1(n42085), .B0(n40171), .B1(n42086),
        .C0(n40300), .C1(n42087), .Y(n18588) );
  OA22X1 U47344 ( .A0(net262475), .A1(n42091), .B0(n42090), .B1(n40119), .Y(
        n18562) );
  CLKINVX1 U47345 ( .A(n18564), .Y(n49615) );
  OAI222XL U47346 ( .A0(net266444), .A1(n42086), .B0(n40171), .B1(n42087),
        .C0(n40300), .C1(n42088), .Y(n18564) );
  OA22X1 U47347 ( .A0(net262475), .A1(n42092), .B0(n42091), .B1(n40119), .Y(
        n18538) );
  CLKINVX1 U47348 ( .A(n18540), .Y(n49617) );
  OAI222XL U47349 ( .A0(net266444), .A1(n42087), .B0(n40171), .B1(n42088),
        .C0(n40300), .C1(n42089), .Y(n18540) );
  OA22X1 U47350 ( .A0(net262475), .A1(n42093), .B0(n42092), .B1(net218912),
        .Y(n18514) );
  CLKINVX1 U47351 ( .A(n18516), .Y(n49619) );
  OAI222XL U47352 ( .A0(net266444), .A1(n42088), .B0(n40171), .B1(n42089),
        .C0(n40300), .C1(n42090), .Y(n18516) );
  OA22X1 U47353 ( .A0(net218338), .A1(n42094), .B0(n42093), .B1(net218912),
        .Y(n18490) );
  CLKINVX1 U47354 ( .A(n18492), .Y(n49621) );
  OAI222XL U47355 ( .A0(net266444), .A1(n42089), .B0(n40171), .B1(n42090),
        .C0(n40300), .C1(n42091), .Y(n18492) );
  OA22X1 U47356 ( .A0(net218564), .A1(n42095), .B0(n42094), .B1(n40118), .Y(
        n18466) );
  CLKINVX1 U47357 ( .A(n18468), .Y(n49623) );
  OAI222XL U47358 ( .A0(net266444), .A1(n42090), .B0(n40171), .B1(n42091),
        .C0(n40300), .C1(n42092), .Y(n18468) );
  OA22X1 U47359 ( .A0(net262513), .A1(n42096), .B0(n42095), .B1(n40118), .Y(
        n18442) );
  CLKINVX1 U47360 ( .A(n18444), .Y(n49625) );
  OAI222XL U47361 ( .A0(net266465), .A1(n42091), .B0(n40171), .B1(n42092),
        .C0(n40300), .C1(n42093), .Y(n18444) );
  OA22X1 U47362 ( .A0(net262513), .A1(n42097), .B0(n42096), .B1(n40091), .Y(
        n18418) );
  CLKINVX1 U47363 ( .A(n18420), .Y(n49627) );
  OAI222XL U47364 ( .A0(net266465), .A1(n42092), .B0(n40170), .B1(n42093),
        .C0(n40299), .C1(n42094), .Y(n18420) );
  OA22X1 U47365 ( .A0(net262798), .A1(n42098), .B0(n42097), .B1(n40106), .Y(
        n18394) );
  CLKINVX1 U47366 ( .A(n18396), .Y(n49629) );
  OAI222XL U47367 ( .A0(net266465), .A1(n42093), .B0(n40170), .B1(n42094),
        .C0(n40299), .C1(n42095), .Y(n18396) );
  OA22X1 U47368 ( .A0(net262798), .A1(n42099), .B0(n42098), .B1(n40106), .Y(
        n18370) );
  CLKINVX1 U47369 ( .A(n18372), .Y(n49631) );
  OAI222XL U47370 ( .A0(net266465), .A1(n42094), .B0(n40170), .B1(n42095),
        .C0(n40299), .C1(n42096), .Y(n18372) );
  OA22X1 U47371 ( .A0(net262817), .A1(n42100), .B0(n42099), .B1(n40105), .Y(
        n18346) );
  CLKINVX1 U47372 ( .A(n18348), .Y(n49633) );
  OAI222XL U47373 ( .A0(net266465), .A1(n42095), .B0(n40170), .B1(n42096),
        .C0(n40299), .C1(n42097), .Y(n18348) );
  OA22X1 U47374 ( .A0(net262817), .A1(n42101), .B0(n42100), .B1(n40105), .Y(
        n18322) );
  CLKINVX1 U47375 ( .A(n18324), .Y(n49635) );
  OAI222XL U47376 ( .A0(net266465), .A1(n42096), .B0(n40170), .B1(n42097),
        .C0(n40299), .C1(n42098), .Y(n18324) );
  OA22X1 U47377 ( .A0(net262836), .A1(n42102), .B0(n42101), .B1(net218632),
        .Y(n18298) );
  CLKINVX1 U47378 ( .A(n18300), .Y(n49637) );
  OAI222XL U47379 ( .A0(net266465), .A1(n42097), .B0(n40170), .B1(n42098),
        .C0(n40299), .C1(n42099), .Y(n18300) );
  OA22X1 U47380 ( .A0(net262836), .A1(n42103), .B0(n42102), .B1(net218628),
        .Y(n18274) );
  CLKINVX1 U47381 ( .A(n18276), .Y(n49639) );
  OAI222XL U47382 ( .A0(net266465), .A1(n42098), .B0(n40170), .B1(n42099),
        .C0(n40299), .C1(n42100), .Y(n18276) );
  OA22X1 U47383 ( .A0(net262836), .A1(n42104), .B0(n42103), .B1(n40104), .Y(
        n18250) );
  CLKINVX1 U47384 ( .A(n18252), .Y(n49641) );
  OAI222XL U47385 ( .A0(net266465), .A1(n42099), .B0(n40170), .B1(n42100),
        .C0(n40299), .C1(n42101), .Y(n18252) );
  OA22X1 U47386 ( .A0(net262855), .A1(n42105), .B0(n42104), .B1(n40104), .Y(
        n18226) );
  CLKINVX1 U47387 ( .A(n18228), .Y(n49643) );
  OAI222XL U47388 ( .A0(net266465), .A1(n42100), .B0(n40170), .B1(n42101),
        .C0(n40299), .C1(n42102), .Y(n18228) );
  OA22X1 U47389 ( .A0(net262855), .A1(n42106), .B0(n42105), .B1(n40103), .Y(
        n18202) );
  CLKINVX1 U47390 ( .A(n18204), .Y(n49645) );
  OAI222XL U47391 ( .A0(net266486), .A1(n42101), .B0(n40169), .B1(n42102),
        .C0(n40298), .C1(n42103), .Y(n18204) );
  OA22X1 U47392 ( .A0(net262874), .A1(n42107), .B0(n42106), .B1(n40102), .Y(
        n18178) );
  CLKINVX1 U47393 ( .A(n18180), .Y(n49647) );
  OAI222XL U47394 ( .A0(net266486), .A1(n42102), .B0(n40169), .B1(n42103),
        .C0(n40298), .C1(n42104), .Y(n18180) );
  OAI211X1 U47395 ( .A0(n42106), .A1(n42830), .B0(n18154), .C0(n49649), .Y(
        n36224) );
  OA22X1 U47396 ( .A0(net262874), .A1(n42108), .B0(n42107), .B1(n40102), .Y(
        n18154) );
  CLKINVX1 U47397 ( .A(n18156), .Y(n49649) );
  OAI222XL U47398 ( .A0(net266486), .A1(n42103), .B0(n40169), .B1(n42104),
        .C0(n40298), .C1(n42105), .Y(n18156) );
  OAI211X1 U47399 ( .A0(n42107), .A1(n42799), .B0(n18130), .C0(n49651), .Y(
        n36216) );
  OA22X1 U47400 ( .A0(net262893), .A1(n42109), .B0(n42108), .B1(n40123), .Y(
        n18130) );
  CLKINVX1 U47401 ( .A(n18132), .Y(n49651) );
  OAI222XL U47402 ( .A0(net266486), .A1(n42104), .B0(n40169), .B1(n42105),
        .C0(n40298), .C1(n42106), .Y(n18132) );
  OA22X1 U47403 ( .A0(net262893), .A1(n42110), .B0(n42109), .B1(net218796),
        .Y(n18106) );
  CLKINVX1 U47404 ( .A(n18108), .Y(n49653) );
  OAI222XL U47405 ( .A0(net266486), .A1(n42105), .B0(n40169), .B1(n42106),
        .C0(n40298), .C1(n42107), .Y(n18108) );
  OA22X1 U47406 ( .A0(net262912), .A1(n42111), .B0(n42110), .B1(n40101), .Y(
        n18082) );
  CLKINVX1 U47407 ( .A(n18084), .Y(n49655) );
  OAI222XL U47408 ( .A0(net266486), .A1(n42106), .B0(n40169), .B1(n42107),
        .C0(n40298), .C1(n42108), .Y(n18084) );
  OA22X1 U47409 ( .A0(net262912), .A1(n42112), .B0(n42111), .B1(n40101), .Y(
        n18058) );
  CLKINVX1 U47410 ( .A(n18060), .Y(n49657) );
  OAI222XL U47411 ( .A0(net266486), .A1(n42107), .B0(n40169), .B1(n42108),
        .C0(n40298), .C1(n42109), .Y(n18060) );
  OA22X1 U47412 ( .A0(net262931), .A1(n42113), .B0(n42112), .B1(n40100), .Y(
        n18034) );
  CLKINVX1 U47413 ( .A(n18036), .Y(n49659) );
  OAI222XL U47414 ( .A0(net266486), .A1(n42108), .B0(n40169), .B1(n42109),
        .C0(n40298), .C1(n42110), .Y(n18036) );
  OA22X1 U47415 ( .A0(net262665), .A1(n42114), .B0(n42113), .B1(n40067), .Y(
        n18010) );
  CLKINVX1 U47416 ( .A(n18012), .Y(n49661) );
  OAI222XL U47417 ( .A0(net266486), .A1(n42109), .B0(n40168), .B1(n42110),
        .C0(n40298), .C1(n42111), .Y(n18012) );
  OA22X1 U47418 ( .A0(net262665), .A1(n42115), .B0(n42114), .B1(n40111), .Y(
        n17986) );
  CLKINVX1 U47419 ( .A(n17988), .Y(n49663) );
  OAI222XL U47420 ( .A0(net266486), .A1(n42110), .B0(n40168), .B1(n42111),
        .C0(n40297), .C1(n42112), .Y(n17988) );
  OAI211X1 U47421 ( .A0(n42114), .A1(n42807), .B0(n17962), .C0(n49665), .Y(
        n36160) );
  OA22X1 U47422 ( .A0(net263406), .A1(n42116), .B0(n42115), .B1(n40111), .Y(
        n17962) );
  CLKINVX1 U47423 ( .A(n17964), .Y(n49665) );
  OAI222XL U47424 ( .A0(net266507), .A1(n42111), .B0(n40168), .B1(n42112),
        .C0(n40297), .C1(n42113), .Y(n17964) );
  OA22X1 U47425 ( .A0(net218344), .A1(n42117), .B0(n42116), .B1(n40110), .Y(
        n17938) );
  CLKINVX1 U47426 ( .A(n17940), .Y(n49667) );
  OAI222XL U47427 ( .A0(net266507), .A1(n42112), .B0(n40168), .B1(n42113),
        .C0(n40297), .C1(n42114), .Y(n17940) );
  OA22X1 U47428 ( .A0(net262703), .A1(n42118), .B0(n42117), .B1(n40110), .Y(
        n17914) );
  CLKINVX1 U47429 ( .A(n17916), .Y(n49669) );
  OAI222XL U47430 ( .A0(net266507), .A1(n42113), .B0(n40168), .B1(n42114),
        .C0(n40297), .C1(n42115), .Y(n17916) );
  OA22X1 U47431 ( .A0(net262703), .A1(n42119), .B0(n42118), .B1(n40109), .Y(
        n17890) );
  CLKINVX1 U47432 ( .A(n17892), .Y(n49671) );
  OAI222XL U47433 ( .A0(net266507), .A1(n42114), .B0(n40168), .B1(n42115),
        .C0(n40297), .C1(n42116), .Y(n17892) );
  OA22X1 U47434 ( .A0(net262703), .A1(n42120), .B0(n42119), .B1(n40109), .Y(
        n17866) );
  CLKINVX1 U47435 ( .A(n17868), .Y(n49673) );
  OAI222XL U47436 ( .A0(net266507), .A1(n42115), .B0(n40168), .B1(n42116),
        .C0(n40297), .C1(n42117), .Y(n17868) );
  OA22X1 U47437 ( .A0(net262722), .A1(n42121), .B0(n42120), .B1(net218750),
        .Y(n17842) );
  CLKINVX1 U47438 ( .A(n17844), .Y(n49675) );
  OAI222XL U47439 ( .A0(net266507), .A1(n42116), .B0(n40168), .B1(n42117),
        .C0(n40297), .C1(n42118), .Y(n17844) );
  OA22X1 U47440 ( .A0(net262722), .A1(n42122), .B0(n42121), .B1(net218838),
        .Y(n17818) );
  CLKINVX1 U47441 ( .A(n17820), .Y(n49677) );
  OAI222XL U47442 ( .A0(net266507), .A1(n42117), .B0(n40168), .B1(n42118),
        .C0(n40297), .C1(n42119), .Y(n17820) );
  OA22X1 U47443 ( .A0(net262741), .A1(n42123), .B0(n42122), .B1(n40108), .Y(
        n17794) );
  CLKINVX1 U47444 ( .A(n17796), .Y(n49679) );
  OAI222XL U47445 ( .A0(net266507), .A1(n42118), .B0(n40167), .B1(n42119),
        .C0(n40297), .C1(n42120), .Y(n17796) );
  OA22X1 U47446 ( .A0(net262741), .A1(n42124), .B0(n42123), .B1(n40108), .Y(
        n17770) );
  CLKINVX1 U47447 ( .A(n17772), .Y(n49681) );
  OAI222XL U47448 ( .A0(net266507), .A1(n42119), .B0(n40167), .B1(n42120),
        .C0(n40296), .C1(n42121), .Y(n17772) );
  OA22X1 U47449 ( .A0(net218506), .A1(n42125), .B0(n42124), .B1(net218628),
        .Y(n17746) );
  CLKINVX1 U47450 ( .A(n17748), .Y(n49683) );
  OAI222XL U47451 ( .A0(net266507), .A1(n42120), .B0(n40167), .B1(n42121),
        .C0(n40296), .C1(n42122), .Y(n17748) );
  OA22X1 U47452 ( .A0(net218442), .A1(n42126), .B0(n42125), .B1(n40068), .Y(
        n17722) );
  CLKINVX1 U47453 ( .A(n17724), .Y(n49685) );
  OAI222XL U47454 ( .A0(net266528), .A1(n42121), .B0(n40167), .B1(n42122),
        .C0(n40296), .C1(n42123), .Y(n17724) );
  OA22X1 U47455 ( .A0(net262779), .A1(n42127), .B0(n42126), .B1(n40107), .Y(
        n17698) );
  CLKINVX1 U47456 ( .A(n17700), .Y(n49687) );
  OAI222XL U47457 ( .A0(net266528), .A1(n42122), .B0(n40167), .B1(n42123),
        .C0(n40296), .C1(n42124), .Y(n17700) );
  OA22X1 U47458 ( .A0(net262779), .A1(n42128), .B0(n42127), .B1(n40107), .Y(
        n17674) );
  CLKINVX1 U47459 ( .A(n17676), .Y(n49689) );
  OAI222XL U47460 ( .A0(net266318), .A1(n42123), .B0(n40167), .B1(n42124),
        .C0(n40296), .C1(n42125), .Y(n17676) );
  OA22X1 U47461 ( .A0(net262779), .A1(n42129), .B0(n42128), .B1(n40106), .Y(
        n17650) );
  CLKINVX1 U47462 ( .A(n17652), .Y(n49691) );
  OAI222XL U47463 ( .A0(net266318), .A1(n42124), .B0(n40178), .B1(n42125),
        .C0(n40296), .C1(n42126), .Y(n17652) );
  OA22X1 U47464 ( .A0(net261981), .A1(n42130), .B0(n42129), .B1(n40144), .Y(
        n17626) );
  CLKINVX1 U47465 ( .A(n17628), .Y(n49693) );
  OAI222XL U47466 ( .A0(net266318), .A1(n42125), .B0(n40179), .B1(n42126),
        .C0(n40296), .C1(n42127), .Y(n17628) );
  OA22X1 U47467 ( .A0(net262000), .A1(n42131), .B0(n42130), .B1(n40144), .Y(
        n17602) );
  CLKINVX1 U47468 ( .A(n17604), .Y(n49695) );
  OAI222XL U47469 ( .A0(net266318), .A1(n42126), .B0(n40179), .B1(n42127),
        .C0(n40296), .C1(n42128), .Y(n17604) );
  OA22X1 U47470 ( .A0(net262000), .A1(n42132), .B0(n42131), .B1(n40143), .Y(
        n17578) );
  CLKINVX1 U47471 ( .A(n17580), .Y(n49697) );
  OAI222XL U47472 ( .A0(net266297), .A1(n42127), .B0(n40179), .B1(n42128),
        .C0(n40296), .C1(n42129), .Y(n17580) );
  OA22X1 U47473 ( .A0(net262000), .A1(n42133), .B0(n42132), .B1(n40143), .Y(
        n17554) );
  CLKINVX1 U47474 ( .A(n17556), .Y(n49699) );
  OAI222XL U47475 ( .A0(net266297), .A1(n42128), .B0(n40179), .B1(n42129),
        .C0(n40295), .C1(n42130), .Y(n17556) );
  OA22X1 U47476 ( .A0(net262019), .A1(n42134), .B0(n42133), .B1(n40068), .Y(
        n17530) );
  CLKINVX1 U47477 ( .A(n17532), .Y(n49701) );
  OAI222XL U47478 ( .A0(net266297), .A1(n42129), .B0(n40179), .B1(n42130),
        .C0(n40295), .C1(n42131), .Y(n17532) );
  OA22X1 U47479 ( .A0(net262019), .A1(n42135), .B0(n42134), .B1(n40068), .Y(
        n17506) );
  CLKINVX1 U47480 ( .A(n17508), .Y(n49703) );
  OAI222XL U47481 ( .A0(net266297), .A1(n42130), .B0(n40179), .B1(n42131),
        .C0(n40295), .C1(n42132), .Y(n17508) );
  OA22X1 U47482 ( .A0(net262038), .A1(n42136), .B0(n42135), .B1(n40142), .Y(
        n17482) );
  CLKINVX1 U47483 ( .A(n17484), .Y(n49705) );
  OAI222XL U47484 ( .A0(net266297), .A1(n42131), .B0(n40179), .B1(n42132),
        .C0(n40295), .C1(n42133), .Y(n17484) );
  OA22X1 U47485 ( .A0(net262038), .A1(n42137), .B0(n42136), .B1(n40142), .Y(
        n17458) );
  CLKINVX1 U47486 ( .A(n17460), .Y(n49707) );
  OAI222XL U47487 ( .A0(net266297), .A1(n42132), .B0(n40179), .B1(n42133),
        .C0(n40295), .C1(n42134), .Y(n17460) );
  OA22X1 U47488 ( .A0(net262057), .A1(n42138), .B0(n42137), .B1(n40141), .Y(
        n17434) );
  CLKINVX1 U47489 ( .A(n17436), .Y(n49709) );
  OAI222XL U47490 ( .A0(net266297), .A1(n42133), .B0(n40179), .B1(n42134),
        .C0(n40295), .C1(n42135), .Y(n17436) );
  OA22X1 U47491 ( .A0(net262057), .A1(n42139), .B0(n42138), .B1(n40140), .Y(
        n17410) );
  CLKINVX1 U47492 ( .A(n17412), .Y(n49711) );
  OAI222XL U47493 ( .A0(net266528), .A1(n42134), .B0(n40180), .B1(n42135),
        .C0(n40295), .C1(n42136), .Y(n17412) );
  OA22X1 U47494 ( .A0(net218308), .A1(n42140), .B0(n42139), .B1(n40140), .Y(
        n17386) );
  CLKINVX1 U47495 ( .A(n17388), .Y(n49713) );
  OAI222XL U47496 ( .A0(net266297), .A1(n42135), .B0(n40180), .B1(n42136),
        .C0(n40295), .C1(n42137), .Y(n17388) );
  OA22X1 U47497 ( .A0(net218406), .A1(n42141), .B0(n42140), .B1(n40087), .Y(
        n17362) );
  CLKINVX1 U47498 ( .A(n17364), .Y(n49715) );
  OAI222XL U47499 ( .A0(net266297), .A1(n42136), .B0(n40180), .B1(n42137),
        .C0(n40295), .C1(n42138), .Y(n17364) );
  OA22X1 U47500 ( .A0(net262095), .A1(n42142), .B0(n42141), .B1(n40068), .Y(
        n17338) );
  CLKINVX1 U47501 ( .A(n17340), .Y(n49717) );
  OAI222XL U47502 ( .A0(net266297), .A1(n42137), .B0(n40180), .B1(n42138),
        .C0(n40294), .C1(n42139), .Y(n17340) );
  OAI211X1 U47503 ( .A0(n42141), .A1(n42838), .B0(n17314), .C0(n49719), .Y(
        n35944) );
  OA22X1 U47504 ( .A0(net262095), .A1(n42143), .B0(n42142), .B1(n40139), .Y(
        n17314) );
  CLKINVX1 U47505 ( .A(n17316), .Y(n49719) );
  OAI222XL U47506 ( .A0(net266276), .A1(n42138), .B0(n40180), .B1(n42139),
        .C0(n40294), .C1(n42140), .Y(n17316) );
  OA22X1 U47507 ( .A0(net262095), .A1(n42144), .B0(n42143), .B1(n40139), .Y(
        n17290) );
  CLKINVX1 U47508 ( .A(n17292), .Y(n49721) );
  OAI222XL U47509 ( .A0(net266276), .A1(n42139), .B0(n40180), .B1(n42140),
        .C0(n40294), .C1(n42141), .Y(n17292) );
  OA22X1 U47510 ( .A0(net262114), .A1(n42145), .B0(n42144), .B1(n40138), .Y(
        n17266) );
  CLKINVX1 U47511 ( .A(n17268), .Y(n49723) );
  OAI222XL U47512 ( .A0(net266276), .A1(n42140), .B0(n40180), .B1(n42141),
        .C0(n40294), .C1(n42142), .Y(n17268) );
  CLKINVX1 U47513 ( .A(n17244), .Y(n49725) );
  OAI222XL U47514 ( .A0(net266276), .A1(n42141), .B0(n40180), .B1(n42142),
        .C0(n40294), .C1(n42143), .Y(n17244) );
  OA22X1 U47515 ( .A0(net261867), .A1(n42147), .B0(n42146), .B1(n40151), .Y(
        n17218) );
  CLKINVX1 U47516 ( .A(n17220), .Y(n49727) );
  OAI222XL U47517 ( .A0(net266276), .A1(n42142), .B0(n40181), .B1(n42143),
        .C0(n40294), .C1(n42144), .Y(n17220) );
  OA22X1 U47518 ( .A0(net261867), .A1(n42148), .B0(n42147), .B1(n40151), .Y(
        n17194) );
  CLKINVX1 U47519 ( .A(n17196), .Y(n49729) );
  OAI222XL U47520 ( .A0(net266276), .A1(n42143), .B0(n40181), .B1(n42144),
        .C0(n40294), .C1(n42145), .Y(n17196) );
  OA22X1 U47521 ( .A0(net261867), .A1(n42149), .B0(n42148), .B1(n40150), .Y(
        n17170) );
  CLKINVX1 U47522 ( .A(n17172), .Y(n49731) );
  OAI222XL U47523 ( .A0(net266276), .A1(n42144), .B0(n40181), .B1(n42145),
        .C0(n40294), .C1(n42146), .Y(n17172) );
  OA22X1 U47524 ( .A0(net261886), .A1(n42150), .B0(n42149), .B1(n40150), .Y(
        n17146) );
  CLKINVX1 U47525 ( .A(n17148), .Y(n49733) );
  OAI222XL U47526 ( .A0(net266276), .A1(n42145), .B0(n40181), .B1(n42146),
        .C0(n40294), .C1(n42147), .Y(n17148) );
  OA22X1 U47527 ( .A0(net261886), .A1(n42151), .B0(n42150), .B1(n40149), .Y(
        n17122) );
  CLKINVX1 U47528 ( .A(n17124), .Y(n49735) );
  OAI222XL U47529 ( .A0(net266276), .A1(n42146), .B0(n40181), .B1(n42147),
        .C0(n40293), .C1(n42148), .Y(n17124) );
  OA22X1 U47530 ( .A0(net261905), .A1(n42152), .B0(n42151), .B1(n40149), .Y(
        n17098) );
  CLKINVX1 U47531 ( .A(n17100), .Y(n49737) );
  OAI222XL U47532 ( .A0(net266255), .A1(n42147), .B0(n40181), .B1(n42148),
        .C0(n40293), .C1(n42149), .Y(n17100) );
  OA22X1 U47533 ( .A0(net261905), .A1(n42153), .B0(n42152), .B1(n40148), .Y(
        n17074) );
  CLKINVX1 U47534 ( .A(n17076), .Y(n49739) );
  OAI222XL U47535 ( .A0(net266255), .A1(n42148), .B0(n40181), .B1(n42149),
        .C0(n40293), .C1(n42150), .Y(n17076) );
  OA22X1 U47536 ( .A0(net261924), .A1(n42154), .B0(n42153), .B1(n40148), .Y(
        n17050) );
  CLKINVX1 U47537 ( .A(n17052), .Y(n49741) );
  OAI222XL U47538 ( .A0(net266255), .A1(n42149), .B0(n40181), .B1(n42150),
        .C0(n40293), .C1(n42151), .Y(n17052) );
  OA22X1 U47539 ( .A0(net261924), .A1(n42155), .B0(n42154), .B1(n40147), .Y(
        n17026) );
  CLKINVX1 U47540 ( .A(n17028), .Y(n49743) );
  OAI222XL U47541 ( .A0(net266255), .A1(n42150), .B0(n40182), .B1(n42151),
        .C0(n40293), .C1(n42152), .Y(n17028) );
  OAI211X1 U47542 ( .A0(n42154), .A1(n42756), .B0(n17002), .C0(n49745), .Y(
        n35840) );
  OA22X1 U47543 ( .A0(net261943), .A1(n42156), .B0(n42155), .B1(n40147), .Y(
        n17002) );
  CLKINVX1 U47544 ( .A(n17004), .Y(n49745) );
  OAI222XL U47545 ( .A0(net266255), .A1(n42151), .B0(n40182), .B1(n42152),
        .C0(n40293), .C1(n42153), .Y(n17004) );
  OA22X1 U47546 ( .A0(net261943), .A1(n42157), .B0(n42156), .B1(n40146), .Y(
        n16978) );
  CLKINVX1 U47547 ( .A(n16980), .Y(n49747) );
  OAI222XL U47548 ( .A0(net266255), .A1(n42152), .B0(n40182), .B1(n42153),
        .C0(n40293), .C1(n42154), .Y(n16980) );
  OA22X1 U47549 ( .A0(net261943), .A1(n42158), .B0(n42157), .B1(n40146), .Y(
        n16954) );
  CLKINVX1 U47550 ( .A(n16956), .Y(n49749) );
  OAI222XL U47551 ( .A0(net266255), .A1(n42153), .B0(n40182), .B1(n42154),
        .C0(n40293), .C1(n42155), .Y(n16956) );
  OA22X1 U47552 ( .A0(net218438), .A1(n42159), .B0(n42158), .B1(n40145), .Y(
        n16930) );
  CLKINVX1 U47553 ( .A(n16932), .Y(n49751) );
  OAI222XL U47554 ( .A0(net266255), .A1(n42154), .B0(n40182), .B1(n42155),
        .C0(n40293), .C1(n42156), .Y(n16932) );
  OA22X1 U47555 ( .A0(net218440), .A1(n42160), .B0(n42159), .B1(n40145), .Y(
        n16906) );
  CLKINVX1 U47556 ( .A(n16908), .Y(n49753) );
  OAI222XL U47557 ( .A0(net266276), .A1(n42155), .B0(n40182), .B1(n42156),
        .C0(net217168), .C1(n42157), .Y(n16908) );
  OA22X1 U47558 ( .A0(net261981), .A1(n42161), .B0(n42160), .B1(n40144), .Y(
        n16882) );
  CLKINVX1 U47559 ( .A(n16884), .Y(n49755) );
  OAI222XL U47560 ( .A0(net266318), .A1(n42156), .B0(n40178), .B1(n42157),
        .C0(net217126), .C1(n42158), .Y(n16884) );
  OA22X1 U47561 ( .A0(net262247), .A1(n42162), .B0(n42161), .B1(n40130), .Y(
        n16858) );
  CLKINVX1 U47562 ( .A(n16860), .Y(n49757) );
  OAI222XL U47563 ( .A0(net266318), .A1(n42157), .B0(n40178), .B1(n42158),
        .C0(net217176), .C1(n42159), .Y(n16860) );
  OA22X1 U47564 ( .A0(net262266), .A1(n42163), .B0(n42162), .B1(n40129), .Y(
        n16834) );
  CLKINVX1 U47565 ( .A(n16836), .Y(n49759) );
  OAI222XL U47566 ( .A0(net266318), .A1(n42158), .B0(n40178), .B1(n42159),
        .C0(net217258), .C1(n42160), .Y(n16836) );
  OA22X1 U47567 ( .A0(net262266), .A1(n42164), .B0(n42163), .B1(n40129), .Y(
        n16810) );
  CLKINVX1 U47568 ( .A(n16812), .Y(n49761) );
  OAI222XL U47569 ( .A0(net266318), .A1(n42159), .B0(n40178), .B1(n42160),
        .C0(net217276), .C1(n42161), .Y(n16812) );
  OA22X1 U47570 ( .A0(net262285), .A1(n42166), .B0(n42165), .B1(n40078), .Y(
        n16762) );
  CLKINVX1 U47571 ( .A(n16764), .Y(n49765) );
  OAI222XL U47572 ( .A0(net266318), .A1(n42161), .B0(n40178), .B1(n42162),
        .C0(net217212), .C1(n42163), .Y(n16764) );
  OA22X1 U47573 ( .A0(net262304), .A1(n42167), .B0(n42166), .B1(n40128), .Y(
        n16738) );
  CLKINVX1 U47574 ( .A(n16740), .Y(n49767) );
  OAI222XL U47575 ( .A0(net266339), .A1(n42162), .B0(n40178), .B1(n42163),
        .C0(net217150), .C1(n42164), .Y(n16740) );
  OA22X1 U47576 ( .A0(net262304), .A1(n42168), .B0(n42167), .B1(n40128), .Y(
        n16714) );
  CLKINVX1 U47577 ( .A(n16716), .Y(n49769) );
  OAI222XL U47578 ( .A0(net266339), .A1(n42163), .B0(n40177), .B1(n42164),
        .C0(net217158), .C1(n42165), .Y(n16716) );
  OA22X1 U47579 ( .A0(net262323), .A1(n42169), .B0(n42168), .B1(n40127), .Y(
        n16690) );
  CLKINVX1 U47580 ( .A(n16692), .Y(n49771) );
  OAI222XL U47581 ( .A0(net266339), .A1(n42164), .B0(n40177), .B1(n42165),
        .C0(n40309), .C1(n42166), .Y(n16692) );
  OAI211X1 U47582 ( .A0(n42168), .A1(n42740), .B0(n16666), .C0(n49773), .Y(
        n35728) );
  OA22X1 U47583 ( .A0(net262323), .A1(n42170), .B0(n42169), .B1(n40127), .Y(
        n16666) );
  CLKINVX1 U47584 ( .A(n16668), .Y(n49773) );
  OAI222XL U47585 ( .A0(net266339), .A1(n42165), .B0(n40177), .B1(n42166),
        .C0(n40309), .C1(n42167), .Y(n16668) );
  OA22X1 U47586 ( .A0(net262323), .A1(n42171), .B0(n42170), .B1(n40126), .Y(
        n16642) );
  CLKINVX1 U47587 ( .A(n16644), .Y(n49775) );
  OAI222XL U47588 ( .A0(net266339), .A1(n42166), .B0(n40177), .B1(n42167),
        .C0(n40309), .C1(n42168), .Y(n16644) );
  OA22X1 U47589 ( .A0(net262342), .A1(n42172), .B0(n42171), .B1(n40126), .Y(
        n16618) );
  CLKINVX1 U47590 ( .A(n16620), .Y(n49777) );
  OAI222XL U47591 ( .A0(net266339), .A1(n42167), .B0(n40177), .B1(n42168),
        .C0(n40309), .C1(n42169), .Y(n16620) );
  OA22X1 U47592 ( .A0(net262342), .A1(n42173), .B0(n42172), .B1(n40125), .Y(
        n16594) );
  CLKINVX1 U47593 ( .A(n16596), .Y(n49779) );
  OAI222XL U47594 ( .A0(net266339), .A1(n42168), .B0(n40177), .B1(n42169),
        .C0(n40309), .C1(n42170), .Y(n16596) );
  OA22X1 U47595 ( .A0(net262361), .A1(n42174), .B0(n42173), .B1(n40125), .Y(
        n16570) );
  CLKINVX1 U47596 ( .A(n16572), .Y(n49781) );
  OAI222XL U47597 ( .A0(net266339), .A1(n42169), .B0(n40177), .B1(n42170),
        .C0(n40309), .C1(n42171), .Y(n16572) );
  OA22X1 U47598 ( .A0(net262361), .A1(n42175), .B0(n42174), .B1(n40124), .Y(
        n16546) );
  CLKINVX1 U47599 ( .A(n16548), .Y(n49783) );
  OAI222XL U47600 ( .A0(net266339), .A1(n42170), .B0(n40177), .B1(n42171),
        .C0(n40309), .C1(n42172), .Y(n16548) );
  OA22X1 U47601 ( .A0(net262380), .A1(n42176), .B0(n42175), .B1(n40124), .Y(
        n16522) );
  CLKINVX1 U47602 ( .A(n16524), .Y(n49785) );
  OAI222XL U47603 ( .A0(net266339), .A1(n42171), .B0(n40177), .B1(n42172),
        .C0(n40309), .C1(n42173), .Y(n16524) );
  OA22X1 U47604 ( .A0(net262380), .A1(n42177), .B0(n42176), .B1(n40123), .Y(
        n16498) );
  CLKINVX1 U47605 ( .A(n16500), .Y(n49787) );
  OAI222XL U47606 ( .A0(net266360), .A1(n42172), .B0(n40176), .B1(n42173),
        .C0(n40309), .C1(n42174), .Y(n16500) );
  OA22X1 U47607 ( .A0(net262114), .A1(n42178), .B0(n42177), .B1(n40138), .Y(
        n16474) );
  CLKINVX1 U47608 ( .A(n16476), .Y(n49789) );
  OAI222XL U47609 ( .A0(net266360), .A1(n42173), .B0(n40176), .B1(n42174),
        .C0(n40310), .C1(n42175), .Y(n16476) );
  OA22X1 U47610 ( .A0(net262133), .A1(n42179), .B0(n42178), .B1(n40137), .Y(
        n16450) );
  CLKINVX1 U47611 ( .A(n16452), .Y(n49791) );
  OAI222XL U47612 ( .A0(net266360), .A1(n42174), .B0(n40176), .B1(n42175),
        .C0(n40310), .C1(n42176), .Y(n16452) );
  OA22X1 U47613 ( .A0(net262133), .A1(n42180), .B0(n42179), .B1(n40137), .Y(
        n16426) );
  CLKINVX1 U47614 ( .A(n16428), .Y(n49793) );
  OAI222XL U47615 ( .A0(net266360), .A1(n42175), .B0(n40176), .B1(n42176),
        .C0(n40310), .C1(n42177), .Y(n16428) );
  OA22X1 U47616 ( .A0(net262152), .A1(n42181), .B0(n42180), .B1(n40136), .Y(
        n16402) );
  CLKINVX1 U47617 ( .A(n16404), .Y(n49795) );
  OAI222XL U47618 ( .A0(net266360), .A1(n42176), .B0(n40176), .B1(n42177),
        .C0(n40310), .C1(n42178), .Y(n16404) );
  OAI211X1 U47619 ( .A0(n42180), .A1(n42786), .B0(n16378), .C0(n49797), .Y(
        n35632) );
  OA22X1 U47620 ( .A0(net262152), .A1(n42182), .B0(n42181), .B1(n40136), .Y(
        n16378) );
  CLKINVX1 U47621 ( .A(n16380), .Y(n49797) );
  OAI222XL U47622 ( .A0(net266360), .A1(n42177), .B0(n40176), .B1(n42178),
        .C0(n40310), .C1(n42179), .Y(n16380) );
  OA22X1 U47623 ( .A0(net262171), .A1(n42183), .B0(n42182), .B1(n40135), .Y(
        n16354) );
  CLKINVX1 U47624 ( .A(n16356), .Y(n49799) );
  OAI222XL U47625 ( .A0(net266360), .A1(n42178), .B0(n40176), .B1(n42179),
        .C0(n40310), .C1(n42180), .Y(n16356) );
  OA22X1 U47626 ( .A0(net262171), .A1(n42184), .B0(n42183), .B1(n40135), .Y(
        n16330) );
  CLKINVX1 U47627 ( .A(n16332), .Y(n49801) );
  OAI222XL U47628 ( .A0(net266360), .A1(n42179), .B0(n40176), .B1(n42180),
        .C0(n40310), .C1(n42181), .Y(n16332) );
  OA22X1 U47629 ( .A0(net262171), .A1(n42185), .B0(n42184), .B1(n40134), .Y(
        n16306) );
  CLKINVX1 U47630 ( .A(n16308), .Y(n49803) );
  OAI222XL U47631 ( .A0(net266360), .A1(n42180), .B0(n40175), .B1(n42181),
        .C0(n40310), .C1(n42182), .Y(n16308) );
  OA22X1 U47632 ( .A0(net262190), .A1(n42186), .B0(n42185), .B1(n40134), .Y(
        n16282) );
  CLKINVX1 U47633 ( .A(n16284), .Y(n49805) );
  OAI222XL U47634 ( .A0(net266360), .A1(n42181), .B0(n40175), .B1(n42182),
        .C0(n40311), .C1(n42183), .Y(n16284) );
  OA22X1 U47635 ( .A0(net262190), .A1(n42187), .B0(n42186), .B1(n40133), .Y(
        n16258) );
  CLKINVX1 U47636 ( .A(n16260), .Y(n49807) );
  OAI222XL U47637 ( .A0(net266381), .A1(n42182), .B0(n40175), .B1(n42183),
        .C0(n40311), .C1(n42184), .Y(n16260) );
  OA22X1 U47638 ( .A0(net262209), .A1(n42188), .B0(n42187), .B1(n40133), .Y(
        n16234) );
  CLKINVX1 U47639 ( .A(n16236), .Y(n49809) );
  OAI222XL U47640 ( .A0(net266381), .A1(n42183), .B0(n40175), .B1(n42184),
        .C0(n40311), .C1(n42185), .Y(n16236) );
  OA22X1 U47641 ( .A0(net262209), .A1(n42189), .B0(n42188), .B1(n40132), .Y(
        n16210) );
  CLKINVX1 U47642 ( .A(n16212), .Y(n49811) );
  OAI222XL U47643 ( .A0(net266381), .A1(n42184), .B0(n40175), .B1(n42185),
        .C0(n40311), .C1(n42186), .Y(n16212) );
  OA22X1 U47644 ( .A0(net262228), .A1(n42190), .B0(n42189), .B1(n40132), .Y(
        n16186) );
  CLKINVX1 U47645 ( .A(n16188), .Y(n49813) );
  OAI222XL U47646 ( .A0(net266381), .A1(n42185), .B0(n40175), .B1(n42186),
        .C0(n40311), .C1(n42187), .Y(n16188) );
  OA22X1 U47647 ( .A0(net262228), .A1(n42191), .B0(n42190), .B1(n40131), .Y(
        n16162) );
  CLKINVX1 U47648 ( .A(n16164), .Y(n49815) );
  OAI222XL U47649 ( .A0(net266381), .A1(n42186), .B0(n40175), .B1(n42187),
        .C0(n40311), .C1(n42188), .Y(n16164) );
  OA22X1 U47650 ( .A0(net262247), .A1(n42192), .B0(n42191), .B1(n40131), .Y(
        n16138) );
  CLKINVX1 U47651 ( .A(n16140), .Y(n49817) );
  OAI222XL U47652 ( .A0(net266381), .A1(n42187), .B0(n40175), .B1(n42188),
        .C0(n40311), .C1(n42189), .Y(n16140) );
  OA22X1 U47653 ( .A0(net262247), .A1(n42193), .B0(n42192), .B1(n40130), .Y(
        n16114) );
  CLKINVX1 U47654 ( .A(n16116), .Y(n49819) );
  OAI222XL U47655 ( .A0(net266381), .A1(n42188), .B0(n40175), .B1(n42189),
        .C0(n40311), .C1(n42190), .Y(n16116) );
  OA22X1 U47656 ( .A0(net263596), .A1(n42194), .B0(n42193), .B1(n40061), .Y(
        n16090) );
  CLKINVX1 U47657 ( .A(n16092), .Y(n49821) );
  OAI222XL U47658 ( .A0(net266654), .A1(n42189), .B0(n40155), .B1(n42190),
        .C0(n40311), .C1(n42191), .Y(n16092) );
  OA22X1 U47659 ( .A0(net263615), .A1(n42195), .B0(n42194), .B1(n40061), .Y(
        n16066) );
  CLKINVX1 U47660 ( .A(n16068), .Y(n49823) );
  OAI222XL U47661 ( .A0(net266654), .A1(n42190), .B0(n40159), .B1(n42191),
        .C0(n40312), .C1(n42192), .Y(n16068) );
  OA22X1 U47662 ( .A0(net263615), .A1(n42196), .B0(n42195), .B1(n40060), .Y(
        n16042) );
  CLKINVX1 U47663 ( .A(n16044), .Y(n49825) );
  OAI222XL U47664 ( .A0(net266675), .A1(n42191), .B0(n40159), .B1(n42192),
        .C0(n40312), .C1(n42193), .Y(n16044) );
  OA22X1 U47665 ( .A0(net263634), .A1(n42197), .B0(n42196), .B1(n40060), .Y(
        n16018) );
  CLKINVX1 U47666 ( .A(n16020), .Y(n49827) );
  OAI222XL U47667 ( .A0(net266675), .A1(n42192), .B0(n40159), .B1(n42193),
        .C0(n40312), .C1(n42194), .Y(n16020) );
  OA22X1 U47668 ( .A0(net263634), .A1(n42198), .B0(n42197), .B1(n40059), .Y(
        n15994) );
  CLKINVX1 U47669 ( .A(n15996), .Y(n49829) );
  OAI222XL U47670 ( .A0(net266675), .A1(n42193), .B0(n40159), .B1(n42194),
        .C0(n40312), .C1(n42195), .Y(n15996) );
  OA22X1 U47671 ( .A0(net263653), .A1(n42199), .B0(n42198), .B1(n40059), .Y(
        n15970) );
  CLKINVX1 U47672 ( .A(n15972), .Y(n49831) );
  OAI222XL U47673 ( .A0(net266675), .A1(n42194), .B0(n40158), .B1(n42195),
        .C0(n40312), .C1(n42196), .Y(n15972) );
  OA22X1 U47674 ( .A0(net263653), .A1(n42200), .B0(n42199), .B1(n40058), .Y(
        n15946) );
  CLKINVX1 U47675 ( .A(n15948), .Y(n49833) );
  OAI222XL U47676 ( .A0(net266675), .A1(n42195), .B0(n40158), .B1(n42196),
        .C0(n40312), .C1(n42197), .Y(n15948) );
  OA22X1 U47677 ( .A0(net263672), .A1(n42201), .B0(n42200), .B1(n40058), .Y(
        n15922) );
  CLKINVX1 U47678 ( .A(n15924), .Y(n49835) );
  OAI222XL U47679 ( .A0(net266675), .A1(n42196), .B0(n40158), .B1(n42197),
        .C0(n40312), .C1(n42198), .Y(n15924) );
  OA22X1 U47680 ( .A0(net263672), .A1(n42202), .B0(n42201), .B1(net218636),
        .Y(n15898) );
  CLKINVX1 U47681 ( .A(n15900), .Y(n49837) );
  OAI222XL U47682 ( .A0(net266675), .A1(n42197), .B0(n40158), .B1(n42198),
        .C0(n40312), .C1(n42199), .Y(n15900) );
  OAI211X1 U47683 ( .A0(n42201), .A1(n42778), .B0(n15874), .C0(n49839), .Y(
        n35464) );
  OA22X1 U47684 ( .A0(net263691), .A1(n42203), .B0(n42202), .B1(n40057), .Y(
        n15874) );
  CLKINVX1 U47685 ( .A(n15876), .Y(n49839) );
  OAI222XL U47686 ( .A0(net266675), .A1(n42198), .B0(n40158), .B1(n42199),
        .C0(n40312), .C1(n42200), .Y(n15876) );
  OA22X1 U47687 ( .A0(net263691), .A1(n42204), .B0(n42203), .B1(n40057), .Y(
        n15850) );
  CLKINVX1 U47688 ( .A(n15852), .Y(n49841) );
  OAI222XL U47689 ( .A0(net266675), .A1(n42199), .B0(n40158), .B1(n42200),
        .C0(n40313), .C1(n42201), .Y(n15852) );
  OA22X1 U47690 ( .A0(net263691), .A1(n42205), .B0(n42204), .B1(n40056), .Y(
        n15826) );
  CLKINVX1 U47691 ( .A(n15828), .Y(n49843) );
  OAI222XL U47692 ( .A0(net266675), .A1(n42200), .B0(n40158), .B1(n42201),
        .C0(n40313), .C1(n42202), .Y(n15828) );
  OA22X1 U47693 ( .A0(net263710), .A1(n42206), .B0(n42205), .B1(n40056), .Y(
        n15802) );
  CLKINVX1 U47694 ( .A(n15804), .Y(n49845) );
  OAI222XL U47695 ( .A0(net266696), .A1(n42201), .B0(n40158), .B1(n42202),
        .C0(net217172), .C1(n42203), .Y(n15804) );
  OA22X1 U47696 ( .A0(net263710), .A1(n42207), .B0(n42206), .B1(n40055), .Y(
        n15778) );
  CLKINVX1 U47697 ( .A(n15780), .Y(n49847) );
  OAI222XL U47698 ( .A0(net266696), .A1(n42202), .B0(n40158), .B1(n42203),
        .C0(n40308), .C1(n42204), .Y(n15780) );
  OA22X1 U47699 ( .A0(net218480), .A1(n42208), .B0(n42207), .B1(n40055), .Y(
        n15754) );
  CLKINVX1 U47700 ( .A(n15756), .Y(n49849) );
  OAI222XL U47701 ( .A0(net266696), .A1(n42203), .B0(n40157), .B1(n42204),
        .C0(n40308), .C1(n42205), .Y(n15756) );
  OA22X1 U47702 ( .A0(net218340), .A1(n42209), .B0(n42208), .B1(n40054), .Y(
        n15730) );
  CLKINVX1 U47703 ( .A(n15732), .Y(n49851) );
  OAI222XL U47704 ( .A0(net266696), .A1(n42204), .B0(n40157), .B1(n42205),
        .C0(n40308), .C1(n42206), .Y(n15732) );
  OA22X1 U47705 ( .A0(net263463), .A1(n42210), .B0(n42209), .B1(n40069), .Y(
        n15706) );
  CLKINVX1 U47706 ( .A(n15708), .Y(n49853) );
  OAI222XL U47707 ( .A0(net266696), .A1(n42205), .B0(n40157), .B1(n42206),
        .C0(n40308), .C1(n42207), .Y(n15708) );
  OA22X1 U47708 ( .A0(net218428), .A1(n42211), .B0(n42210), .B1(n40068), .Y(
        n15682) );
  CLKINVX1 U47709 ( .A(n15684), .Y(n49855) );
  OAI222XL U47710 ( .A0(net266696), .A1(n42206), .B0(n40157), .B1(n42207),
        .C0(n40308), .C1(n42208), .Y(n15684) );
  OAI211X1 U47711 ( .A0(n42210), .A1(n42949), .B0(n15658), .C0(n49857), .Y(
        n35392) );
  OA22X1 U47712 ( .A0(net263178), .A1(n42212), .B0(n42211), .B1(n40068), .Y(
        n15658) );
  CLKINVX1 U47713 ( .A(n15660), .Y(n49857) );
  OAI222XL U47714 ( .A0(net266696), .A1(n42207), .B0(n40157), .B1(n42208),
        .C0(n40308), .C1(n42209), .Y(n15660) );
  OA22X1 U47715 ( .A0(net263501), .A1(n42213), .B0(n42212), .B1(n40067), .Y(
        n15634) );
  CLKINVX1 U47716 ( .A(n15636), .Y(n49859) );
  OAI222XL U47717 ( .A0(net266696), .A1(n42208), .B0(n40157), .B1(n42209),
        .C0(n40308), .C1(n42210), .Y(n15636) );
  OA22X1 U47718 ( .A0(net263501), .A1(n42214), .B0(n42213), .B1(n40067), .Y(
        n15610) );
  CLKINVX1 U47719 ( .A(n15612), .Y(n49861) );
  OAI222XL U47720 ( .A0(net266696), .A1(n42209), .B0(n40157), .B1(n42210),
        .C0(n40308), .C1(n42211), .Y(n15612) );
  OA22X1 U47721 ( .A0(net218572), .A1(n42215), .B0(n42214), .B1(n40066), .Y(
        n15586) );
  CLKINVX1 U47722 ( .A(n15588), .Y(n49863) );
  OAI222XL U47723 ( .A0(net266696), .A1(n42210), .B0(n40157), .B1(n42211),
        .C0(n40308), .C1(n42212), .Y(n15588) );
  OA22X1 U47724 ( .A0(net218526), .A1(n42216), .B0(n42215), .B1(n40066), .Y(
        n15562) );
  CLKINVX1 U47725 ( .A(n15564), .Y(n49865) );
  OAI222XL U47726 ( .A0(net266717), .A1(n42211), .B0(n40156), .B1(n42212),
        .C0(n40307), .C1(n42213), .Y(n15564) );
  OA22X1 U47727 ( .A0(net263539), .A1(n42217), .B0(n42216), .B1(n40065), .Y(
        n15538) );
  CLKINVX1 U47728 ( .A(n15540), .Y(n49867) );
  OAI222XL U47729 ( .A0(net266717), .A1(n42212), .B0(n40156), .B1(n42213),
        .C0(n40307), .C1(n42214), .Y(n15540) );
  OA22X1 U47730 ( .A0(net263539), .A1(n42218), .B0(n42217), .B1(n40065), .Y(
        n15514) );
  CLKINVX1 U47731 ( .A(n15516), .Y(n49869) );
  OAI222XL U47732 ( .A0(net266717), .A1(n42213), .B0(n40156), .B1(n42214),
        .C0(n40307), .C1(n42215), .Y(n15516) );
  OA22X1 U47733 ( .A0(net263539), .A1(n42219), .B0(n42218), .B1(n40064), .Y(
        n15490) );
  CLKINVX1 U47734 ( .A(n15492), .Y(n49871) );
  OAI222XL U47735 ( .A0(net266717), .A1(n42214), .B0(n40156), .B1(n42215),
        .C0(n40307), .C1(n42216), .Y(n15492) );
  OAI211X1 U47736 ( .A0(n42218), .A1(n42958), .B0(n15466), .C0(n49873), .Y(
        n35328) );
  OA22X1 U47737 ( .A0(net263558), .A1(n42220), .B0(n42219), .B1(n40064), .Y(
        n15466) );
  OAI222XL U47738 ( .A0(net266717), .A1(n42215), .B0(n40156), .B1(n42216),
        .C0(n40307), .C1(n42217), .Y(n15468) );
  OAI211X1 U47739 ( .A0(n42219), .A1(n42959), .B0(n15442), .C0(n49875), .Y(
        n35320) );
  OA22X1 U47740 ( .A0(net263558), .A1(n42221), .B0(n42220), .B1(n40063), .Y(
        n15442) );
  OAI222XL U47741 ( .A0(net266717), .A1(n42216), .B0(n40156), .B1(n42217),
        .C0(n40307), .C1(n42218), .Y(n15444) );
  OAI211X1 U47742 ( .A0(n42220), .A1(n42928), .B0(n15418), .C0(n49877), .Y(
        n35312) );
  OA22X1 U47743 ( .A0(net263577), .A1(n42222), .B0(n42221), .B1(n40063), .Y(
        n15418) );
  OAI222XL U47744 ( .A0(net266717), .A1(n42217), .B0(n40156), .B1(n42218),
        .C0(n40307), .C1(n42219), .Y(n15420) );
  OAI211X1 U47745 ( .A0(n42221), .A1(n42929), .B0(n15394), .C0(n49879), .Y(
        n35304) );
  OA22X1 U47746 ( .A0(net263577), .A1(n42223), .B0(n42222), .B1(n40062), .Y(
        n15394) );
  OAI222XL U47747 ( .A0(net266717), .A1(n42218), .B0(n40156), .B1(n42219),
        .C0(n40307), .C1(n42220), .Y(n15396) );
  OAI211X1 U47748 ( .A0(n42222), .A1(n42931), .B0(n15370), .C0(n49881), .Y(
        n35296) );
  OA22X1 U47749 ( .A0(net263596), .A1(n42224), .B0(n42223), .B1(n40062), .Y(
        n15370) );
  OAI222XL U47750 ( .A0(net266717), .A1(n42219), .B0(n40156), .B1(n42220),
        .C0(n40307), .C1(n42221), .Y(n15372) );
  OAI211X1 U47751 ( .A0(n42223), .A1(n42932), .B0(n15346), .C0(n49883), .Y(
        n35288) );
  OA22X1 U47752 ( .A0(net263596), .A1(n42225), .B0(n42224), .B1(n40061), .Y(
        n15346) );
  OAI222XL U47753 ( .A0(net266717), .A1(n42220), .B0(n40155), .B1(n42221),
        .C0(n40306), .C1(n42222), .Y(n15348) );
  OAI211X1 U47754 ( .A0(n42224), .A1(n42933), .B0(n15322), .C0(n49885), .Y(
        n35280) );
  OA22X1 U47755 ( .A0(net263881), .A1(n42226), .B0(n42225), .B1(n40046), .Y(
        n15322) );
  OAI222XL U47756 ( .A0(net266738), .A1(n42221), .B0(n40155), .B1(n42222),
        .C0(n40306), .C1(n42223), .Y(n15324) );
  OAI211X1 U47757 ( .A0(n42225), .A1(n42934), .B0(n15298), .C0(n49887), .Y(
        n35272) );
  OA22X1 U47758 ( .A0(net263881), .A1(n42227), .B0(n42226), .B1(n40045), .Y(
        n15298) );
  OAI222XL U47759 ( .A0(net266738), .A1(n42222), .B0(n40155), .B1(n42223),
        .C0(n40306), .C1(n42224), .Y(n15300) );
  OAI211X1 U47760 ( .A0(n42226), .A1(n42935), .B0(n15274), .C0(n49889), .Y(
        n35264) );
  OA22X1 U47761 ( .A0(net263900), .A1(n42228), .B0(n42227), .B1(n40045), .Y(
        n15274) );
  OAI222XL U47762 ( .A0(net266738), .A1(n42223), .B0(n40155), .B1(n42224),
        .C0(n40306), .C1(n42225), .Y(n15276) );
  OAI211X1 U47763 ( .A0(n42227), .A1(n42936), .B0(n15250), .C0(n49891), .Y(
        n35256) );
  OA22X1 U47764 ( .A0(net263900), .A1(n42229), .B0(n42228), .B1(n40044), .Y(
        n15250) );
  OAI222XL U47765 ( .A0(net266738), .A1(n42224), .B0(n40155), .B1(n42225),
        .C0(n40306), .C1(n42226), .Y(n15252) );
  OAI211X1 U47766 ( .A0(n42228), .A1(n42938), .B0(n15226), .C0(n49893), .Y(
        n35248) );
  OA22X1 U47767 ( .A0(net263919), .A1(n42230), .B0(n42229), .B1(n40044), .Y(
        n15226) );
  OAI222XL U47768 ( .A0(net266738), .A1(n42225), .B0(n40155), .B1(n42226),
        .C0(n40306), .C1(n42227), .Y(n15228) );
  OAI211X1 U47769 ( .A0(n42229), .A1(n42939), .B0(n15202), .C0(n49895), .Y(
        n35240) );
  OA22X1 U47770 ( .A0(net263919), .A1(n42231), .B0(n42230), .B1(n40043), .Y(
        n15202) );
  OAI222XL U47771 ( .A0(net266738), .A1(n42226), .B0(n40155), .B1(n42227),
        .C0(n40306), .C1(n42228), .Y(n15204) );
  OAI211X1 U47772 ( .A0(n42230), .A1(n42940), .B0(n15178), .C0(n49897), .Y(
        n35232) );
  OA22X1 U47773 ( .A0(net263919), .A1(n42232), .B0(n42231), .B1(n40043), .Y(
        n15178) );
  OAI222XL U47774 ( .A0(net266738), .A1(n42227), .B0(n40154), .B1(n42228),
        .C0(n40306), .C1(n42229), .Y(n15180) );
  OAI211X1 U47775 ( .A0(n42231), .A1(n42941), .B0(n15154), .C0(n49899), .Y(
        n35224) );
  OA22X1 U47776 ( .A0(net262931), .A1(n42233), .B0(n42232), .B1(n40069), .Y(
        n15154) );
  OAI222XL U47777 ( .A0(net266738), .A1(n42228), .B0(n40154), .B1(n42229),
        .C0(n40306), .C1(n42230), .Y(n15156) );
  OAI211X1 U47778 ( .A0(n42232), .A1(n42942), .B0(n15130), .C0(n49901), .Y(
        n35216) );
  OA22X1 U47779 ( .A0(net262931), .A1(n42234), .B0(n42233), .B1(n40069), .Y(
        n15130) );
  OAI222XL U47780 ( .A0(net266738), .A1(n42229), .B0(n40154), .B1(n42230),
        .C0(n40305), .C1(n42231), .Y(n15132) );
  OAI211X1 U47781 ( .A0(n42233), .A1(n42943), .B0(n15106), .C0(n49903), .Y(
        n35208) );
  OA22X1 U47782 ( .A0(net263957), .A1(n42235), .B0(n42234), .B1(n40042), .Y(
        n15106) );
  OAI222XL U47783 ( .A0(net266759), .A1(n42230), .B0(n40154), .B1(n42231),
        .C0(n40305), .C1(n42232), .Y(n15108) );
  OAI211X1 U47784 ( .A0(n42234), .A1(n42977), .B0(n15082), .C0(n49905), .Y(
        n35200) );
  OA22X1 U47785 ( .A0(net263957), .A1(n42236), .B0(n42235), .B1(n40042), .Y(
        n15082) );
  OAI222XL U47786 ( .A0(net266759), .A1(n42231), .B0(n40154), .B1(n42232),
        .C0(n40305), .C1(n42233), .Y(n15084) );
  OAI211X1 U47787 ( .A0(n42235), .A1(n42978), .B0(n15058), .C0(n49907), .Y(
        n35192) );
  OA22X1 U47788 ( .A0(net263976), .A1(n42237), .B0(n42236), .B1(n40041), .Y(
        n15058) );
  OAI222XL U47789 ( .A0(net266759), .A1(n42232), .B0(n40154), .B1(n42233),
        .C0(n40305), .C1(n42234), .Y(n15060) );
  OAI211X1 U47790 ( .A0(n42236), .A1(n42979), .B0(n15034), .C0(n49909), .Y(
        n35184) );
  OA22X1 U47791 ( .A0(net263976), .A1(n42238), .B0(n42237), .B1(n40041), .Y(
        n15034) );
  OAI222XL U47792 ( .A0(net266759), .A1(n42233), .B0(n40154), .B1(n42234),
        .C0(n40305), .C1(n42235), .Y(n15036) );
  OAI211X1 U47793 ( .A0(n42237), .A1(n42980), .B0(n15010), .C0(n49911), .Y(
        n35176) );
  OA22X1 U47794 ( .A0(net263995), .A1(n42239), .B0(n42238), .B1(n40040), .Y(
        n15010) );
  OAI222XL U47795 ( .A0(net266738), .A1(n42234), .B0(n40154), .B1(n42235),
        .C0(n40305), .C1(n42236), .Y(n15012) );
  OAI211X1 U47796 ( .A0(n42238), .A1(n42981), .B0(n14986), .C0(n49913), .Y(
        n35168) );
  OA22X1 U47797 ( .A0(net263995), .A1(n42240), .B0(n42239), .B1(n40040), .Y(
        n14986) );
  OAI222XL U47798 ( .A0(net266759), .A1(n42235), .B0(n40154), .B1(n42236),
        .C0(n40305), .C1(n42237), .Y(n14988) );
  OAI211X1 U47799 ( .A0(n42239), .A1(n42982), .B0(n14962), .C0(n49915), .Y(
        n35160) );
  OA22X1 U47800 ( .A0(net263995), .A1(n42241), .B0(n42240), .B1(net218866),
        .Y(n14962) );
  OAI222XL U47801 ( .A0(net266759), .A1(n42236), .B0(n40153), .B1(n42237),
        .C0(n40305), .C1(n42238), .Y(n14964) );
  OAI211X1 U47802 ( .A0(n42240), .A1(n42983), .B0(n14938), .C0(n49917), .Y(
        n35152) );
  OA22X1 U47803 ( .A0(net263748), .A1(n42242), .B0(n42241), .B1(n40054), .Y(
        n14938) );
  OAI222XL U47804 ( .A0(net266759), .A1(n42237), .B0(n40153), .B1(n42238),
        .C0(n40305), .C1(n42239), .Y(n14940) );
  OAI211X1 U47805 ( .A0(n42241), .A1(n42985), .B0(n14914), .C0(n49919), .Y(
        n35144) );
  OA22X1 U47806 ( .A0(net263748), .A1(n42243), .B0(n42242), .B1(n40053), .Y(
        n14914) );
  OAI222XL U47807 ( .A0(net266759), .A1(n42238), .B0(n40153), .B1(n42239),
        .C0(n40304), .C1(n42240), .Y(n14916) );
  OAI211X1 U47808 ( .A0(n42242), .A1(n42986), .B0(n14890), .C0(n49921), .Y(
        n35136) );
  OA22X1 U47809 ( .A0(net263767), .A1(n42244), .B0(n42243), .B1(n40053), .Y(
        n14890) );
  OAI222XL U47810 ( .A0(net266759), .A1(n42239), .B0(n40153), .B1(n42240),
        .C0(n40304), .C1(n42241), .Y(n14892) );
  OAI211X1 U47811 ( .A0(n42243), .A1(n42987), .B0(n14866), .C0(n49923), .Y(
        n35128) );
  OA22X1 U47812 ( .A0(net263767), .A1(n42245), .B0(n42244), .B1(n40052), .Y(
        n14866) );
  OAI222XL U47813 ( .A0(net266780), .A1(n42240), .B0(n40153), .B1(n42241),
        .C0(n40304), .C1(n42242), .Y(n14868) );
  OAI211X1 U47814 ( .A0(n42244), .A1(n42988), .B0(n14842), .C0(n49925), .Y(
        n35120) );
  OA22X1 U47815 ( .A0(net263767), .A1(n42246), .B0(n42245), .B1(n40052), .Y(
        n14842) );
  OAI222XL U47816 ( .A0(net266780), .A1(n42241), .B0(n40153), .B1(n42242),
        .C0(n40304), .C1(n42243), .Y(n14844) );
  OAI211X1 U47817 ( .A0(n42245), .A1(n42989), .B0(n14818), .C0(n49927), .Y(
        n35112) );
  OA22X1 U47818 ( .A0(net218478), .A1(n42247), .B0(n42246), .B1(n40051), .Y(
        n14818) );
  OAI222XL U47819 ( .A0(net266780), .A1(n42242), .B0(n40153), .B1(n42243),
        .C0(n40304), .C1(n42244), .Y(n14820) );
  OAI211X1 U47820 ( .A0(n42246), .A1(n42990), .B0(n14794), .C0(n49929), .Y(
        n35104) );
  OA22X1 U47821 ( .A0(net218376), .A1(n42248), .B0(n42247), .B1(n40051), .Y(
        n14794) );
  OAI222XL U47822 ( .A0(net266780), .A1(n42243), .B0(n40153), .B1(n42244),
        .C0(n40304), .C1(n42245), .Y(n14796) );
  OAI211X1 U47823 ( .A0(n42247), .A1(n42965), .B0(n14770), .C0(n49931), .Y(
        n35096) );
  OA22X1 U47824 ( .A0(net263805), .A1(n42249), .B0(n42248), .B1(n40050), .Y(
        n14770) );
  OAI222XL U47825 ( .A0(net266780), .A1(n42244), .B0(n40152), .B1(n42245),
        .C0(n40304), .C1(n42246), .Y(n14772) );
  OAI211X1 U47826 ( .A0(n42248), .A1(n42960), .B0(n14746), .C0(n49933), .Y(
        n35088) );
  OA22X1 U47827 ( .A0(net263805), .A1(n42250), .B0(n42249), .B1(n40050), .Y(
        n14746) );
  OAI222XL U47828 ( .A0(net266780), .A1(n42245), .B0(n40152), .B1(n42246),
        .C0(n40304), .C1(n42247), .Y(n14748) );
  OAI211X1 U47829 ( .A0(n42249), .A1(n42962), .B0(n14722), .C0(n49935), .Y(
        n35080) );
  OA22X1 U47830 ( .A0(net263824), .A1(n42251), .B0(n42250), .B1(n40049), .Y(
        n14722) );
  OAI222XL U47831 ( .A0(net266780), .A1(n42246), .B0(n40152), .B1(n42247),
        .C0(n40304), .C1(n42248), .Y(n14724) );
  OAI211X1 U47832 ( .A0(n42250), .A1(n42963), .B0(n14698), .C0(n49937), .Y(
        n35072) );
  OA22X1 U47833 ( .A0(net263824), .A1(n42252), .B0(n42251), .B1(n40049), .Y(
        n14698) );
  OAI222XL U47834 ( .A0(net266780), .A1(n42247), .B0(n40152), .B1(n42248),
        .C0(n40303), .C1(n42249), .Y(n14700) );
  OAI211X1 U47835 ( .A0(n42251), .A1(n42964), .B0(n14674), .C0(n49939), .Y(
        n35064) );
  OA22X1 U47836 ( .A0(net263843), .A1(n42253), .B0(n42252), .B1(n40048), .Y(
        n14674) );
  OAI222XL U47837 ( .A0(net266780), .A1(n42248), .B0(n40152), .B1(n42249),
        .C0(n40303), .C1(n42250), .Y(n14676) );
  OAI211X1 U47838 ( .A0(n42252), .A1(n42965), .B0(n14650), .C0(n49941), .Y(
        n35056) );
  OA22X1 U47839 ( .A0(net263843), .A1(n42254), .B0(n42253), .B1(n40048), .Y(
        n14650) );
  OAI222XL U47840 ( .A0(net266780), .A1(n42249), .B0(n40152), .B1(n42250),
        .C0(n40303), .C1(n42251), .Y(n14652) );
  OAI211X1 U47841 ( .A0(n42253), .A1(n42966), .B0(n14626), .C0(n49943), .Y(
        n35048) );
  OA22X1 U47842 ( .A0(net263862), .A1(n42255), .B0(n42254), .B1(n40047), .Y(
        n14626) );
  OAI222XL U47843 ( .A0(net266780), .A1(n42250), .B0(n40152), .B1(n42251),
        .C0(n40288), .C1(n42252), .Y(n14628) );
  OAI211X1 U47844 ( .A0(n42254), .A1(n42967), .B0(n14602), .C0(n49945), .Y(
        n35040) );
  OA22X1 U47845 ( .A0(net263862), .A1(n42256), .B0(n42255), .B1(n40047), .Y(
        n14602) );
  OAI222XL U47846 ( .A0(net266780), .A1(n42251), .B0(n40152), .B1(n42252),
        .C0(n40288), .C1(n42253), .Y(n14604) );
  OAI211X1 U47847 ( .A0(n42255), .A1(n42969), .B0(n14578), .C0(n49947), .Y(
        n35032) );
  OA22X1 U47848 ( .A0(net263862), .A1(n42257), .B0(n42256), .B1(n40046), .Y(
        n14578) );
  OAI222XL U47849 ( .A0(net266780), .A1(n42252), .B0(n40152), .B1(n42253),
        .C0(n40288), .C1(n42254), .Y(n14580) );
  OAI211X1 U47850 ( .A0(n42256), .A1(n42970), .B0(n14554), .C0(n49949), .Y(
        n35024) );
  OA22X1 U47851 ( .A0(net263064), .A1(n42258), .B0(n42257), .B1(n40092), .Y(
        n14554) );
  CLKINVX1 U47852 ( .A(n14556), .Y(n49949) );
  OAI222XL U47853 ( .A0(net221954), .A1(n42253), .B0(net218220), .B1(n42254),
        .C0(n40288), .C1(n42255), .Y(n14556) );
  OAI211X1 U47854 ( .A0(n42257), .A1(n42971), .B0(n14530), .C0(n49951), .Y(
        n35016) );
  OA22X1 U47855 ( .A0(net263083), .A1(n42259), .B0(n42258), .B1(n40091), .Y(
        n14530) );
  OAI222XL U47856 ( .A0(net266591), .A1(n42254), .B0(n40163), .B1(n42255),
        .C0(n40288), .C1(n42256), .Y(n14532) );
  OAI211X1 U47857 ( .A0(n42258), .A1(n42972), .B0(n14506), .C0(n49953), .Y(
        n35008) );
  OA22X1 U47858 ( .A0(net263083), .A1(n42260), .B0(n42259), .B1(n40091), .Y(
        n14506) );
  OAI222XL U47859 ( .A0(net266528), .A1(n42255), .B0(n40167), .B1(n42256),
        .C0(n40288), .C1(n42257), .Y(n14508) );
  OAI211X1 U47860 ( .A0(n42259), .A1(n42973), .B0(n14482), .C0(n49955), .Y(
        n35000) );
  OA22X1 U47861 ( .A0(net263083), .A1(n42261), .B0(n42260), .B1(n40090), .Y(
        n14482) );
  OAI222XL U47862 ( .A0(net266528), .A1(n42256), .B0(n40167), .B1(n42257),
        .C0(n40288), .C1(n42258), .Y(n14484) );
  OAI211X1 U47863 ( .A0(n42260), .A1(n42974), .B0(n14458), .C0(n49957), .Y(
        n34992) );
  OA22X1 U47864 ( .A0(net263102), .A1(n42262), .B0(n42261), .B1(n40090), .Y(
        n14458) );
  OAI222XL U47865 ( .A0(net266528), .A1(n42257), .B0(n40166), .B1(n42258),
        .C0(n40288), .C1(n42259), .Y(n14460) );
  OAI211X1 U47866 ( .A0(n42261), .A1(n42975), .B0(n14434), .C0(n49959), .Y(
        n34984) );
  OA22X1 U47867 ( .A0(net263102), .A1(n42263), .B0(n42262), .B1(n40089), .Y(
        n14434) );
  OAI222XL U47868 ( .A0(net266528), .A1(n42258), .B0(n40166), .B1(n42259),
        .C0(n40288), .C1(n42260), .Y(n14436) );
  OAI211X1 U47869 ( .A0(n42262), .A1(n42879), .B0(n14410), .C0(n49961), .Y(
        n34976) );
  OA22X1 U47870 ( .A0(net263121), .A1(n42264), .B0(n42263), .B1(n40089), .Y(
        n14410) );
  OAI222XL U47871 ( .A0(net266528), .A1(n42259), .B0(n40166), .B1(n42260),
        .C0(n40287), .C1(n42261), .Y(n14412) );
  OAI211X1 U47872 ( .A0(n42263), .A1(n42881), .B0(n14386), .C0(n49963), .Y(
        n34968) );
  OA22X1 U47873 ( .A0(net263121), .A1(n42265), .B0(n42264), .B1(n40088), .Y(
        n14386) );
  OAI222XL U47874 ( .A0(net266528), .A1(n42260), .B0(n40166), .B1(n42261),
        .C0(n40287), .C1(n42262), .Y(n14388) );
  OAI211X1 U47875 ( .A0(n42264), .A1(n42882), .B0(n14362), .C0(n49965), .Y(
        n34960) );
  OA22X1 U47876 ( .A0(net263140), .A1(n42266), .B0(n42265), .B1(n40088), .Y(
        n14362) );
  OAI222XL U47877 ( .A0(net266528), .A1(n42261), .B0(n40166), .B1(n42262),
        .C0(n40287), .C1(n42263), .Y(n14364) );
  OAI211X1 U47878 ( .A0(n42265), .A1(n42883), .B0(n14338), .C0(n49967), .Y(
        n34952) );
  OA22X1 U47879 ( .A0(net263140), .A1(n42267), .B0(n42266), .B1(n40087), .Y(
        n14338) );
  OAI222XL U47880 ( .A0(net266549), .A1(n42262), .B0(n40166), .B1(n42263),
        .C0(n40287), .C1(n42264), .Y(n14340) );
  OAI211X1 U47881 ( .A0(n42266), .A1(n42884), .B0(n14314), .C0(n49969), .Y(
        n34944) );
  OA22X1 U47882 ( .A0(net263159), .A1(n42268), .B0(n42267), .B1(n40087), .Y(
        n14314) );
  OAI222XL U47883 ( .A0(net266549), .A1(n42263), .B0(n40166), .B1(n42264),
        .C0(n40287), .C1(n42265), .Y(n14316) );
  OAI211X1 U47884 ( .A0(n42267), .A1(n42885), .B0(n14290), .C0(n49971), .Y(
        n34936) );
  OA22X1 U47885 ( .A0(net263159), .A1(n42269), .B0(n42268), .B1(n40086), .Y(
        n14290) );
  OAI222XL U47886 ( .A0(net266549), .A1(n42264), .B0(n40166), .B1(n42265),
        .C0(n40287), .C1(n42266), .Y(n14292) );
  OAI211X1 U47887 ( .A0(n42268), .A1(n42886), .B0(n14266), .C0(n49973), .Y(
        n34928) );
  OA22X1 U47888 ( .A0(net263159), .A1(n42270), .B0(n42269), .B1(n40086), .Y(
        n14266) );
  OAI222XL U47889 ( .A0(net266549), .A1(n42265), .B0(n40165), .B1(n42266),
        .C0(n40287), .C1(n42267), .Y(n14268) );
  OAI211X1 U47890 ( .A0(n42269), .A1(n42888), .B0(n14242), .C0(n49975), .Y(
        n34920) );
  OA22X1 U47891 ( .A0(net263178), .A1(n42271), .B0(n42270), .B1(n40085), .Y(
        n14242) );
  OAI222XL U47892 ( .A0(net266549), .A1(n42266), .B0(n40165), .B1(n42267),
        .C0(n40287), .C1(n42268), .Y(n14244) );
  OAI211X1 U47893 ( .A0(n42270), .A1(n42889), .B0(n14218), .C0(n49977), .Y(
        n34912) );
  OA22X1 U47894 ( .A0(net263178), .A1(n42272), .B0(n42271), .B1(n40085), .Y(
        n14218) );
  OAI222XL U47895 ( .A0(net266549), .A1(n42267), .B0(n40165), .B1(n42268),
        .C0(n40287), .C1(n42269), .Y(n14220) );
  OAI211X1 U47896 ( .A0(n42271), .A1(n42890), .B0(n14194), .C0(n49979), .Y(
        n34904) );
  OA22X1 U47897 ( .A0(net218394), .A1(n42273), .B0(n42272), .B1(n40084), .Y(
        n14194) );
  OAI222XL U47898 ( .A0(net266549), .A1(n42268), .B0(n40165), .B1(n42269),
        .C0(n40286), .C1(n42270), .Y(n14196) );
  OAI211X1 U47899 ( .A0(n42272), .A1(n42891), .B0(n14170), .C0(n49981), .Y(
        n34896) );
  OA22X1 U47900 ( .A0(net262931), .A1(n42274), .B0(n42273), .B1(n40100), .Y(
        n14170) );
  OAI222XL U47901 ( .A0(net266549), .A1(n42269), .B0(n40165), .B1(n42270),
        .C0(n40286), .C1(n42271), .Y(n14172) );
  OAI211X1 U47902 ( .A0(n42273), .A1(n42892), .B0(n14146), .C0(n49983), .Y(
        n34888) );
  OA22X1 U47903 ( .A0(net262931), .A1(n42275), .B0(n42274), .B1(n40099), .Y(
        n14146) );
  OAI222XL U47904 ( .A0(net266549), .A1(n42270), .B0(n40165), .B1(n42271),
        .C0(n40286), .C1(n42272), .Y(n14148) );
  OAI211X1 U47905 ( .A0(n42274), .A1(n42893), .B0(n14122), .C0(n49985), .Y(
        n34880) );
  OA22X1 U47906 ( .A0(net262950), .A1(n42276), .B0(n42275), .B1(n40099), .Y(
        n14122) );
  OAI222XL U47907 ( .A0(net266549), .A1(n42271), .B0(n40165), .B1(n42272),
        .C0(n40286), .C1(n42273), .Y(n14124) );
  OAI211X1 U47908 ( .A0(n42275), .A1(n42894), .B0(n14098), .C0(n49987), .Y(
        n34872) );
  OA22X1 U47909 ( .A0(net262950), .A1(n42277), .B0(n42276), .B1(n40098), .Y(
        n14098) );
  OAI222XL U47910 ( .A0(net266570), .A1(n42272), .B0(n40165), .B1(n42273),
        .C0(n40286), .C1(n42274), .Y(n14100) );
  OAI211X1 U47911 ( .A0(n42276), .A1(n42863), .B0(n14074), .C0(n49989), .Y(
        n34864) );
  OA22X1 U47912 ( .A0(net262969), .A1(n42278), .B0(n42277), .B1(n40098), .Y(
        n14074) );
  OAI222XL U47913 ( .A0(net266570), .A1(n42273), .B0(n40165), .B1(n42274),
        .C0(n40286), .C1(n42275), .Y(n14076) );
  OAI211X1 U47914 ( .A0(n42277), .A1(n42865), .B0(n14050), .C0(n49991), .Y(
        n34856) );
  OA22X1 U47915 ( .A0(net262969), .A1(n42279), .B0(n42278), .B1(n40097), .Y(
        n14050) );
  OAI222XL U47916 ( .A0(net266570), .A1(n42274), .B0(n40164), .B1(n42275),
        .C0(n40286), .C1(n42276), .Y(n14052) );
  OAI211X1 U47917 ( .A0(n42278), .A1(n42866), .B0(n14026), .C0(n49993), .Y(
        n34848) );
  OA22X1 U47918 ( .A0(net262988), .A1(n42280), .B0(n42279), .B1(n40097), .Y(
        n14026) );
  OAI222XL U47919 ( .A0(net266570), .A1(n42275), .B0(n40164), .B1(n42276),
        .C0(n40286), .C1(n42277), .Y(n14028) );
  OAI211X1 U47920 ( .A0(n42279), .A1(n42867), .B0(n14002), .C0(n49995), .Y(
        n34840) );
  OA22X1 U47921 ( .A0(net262988), .A1(n42281), .B0(n42280), .B1(n40096), .Y(
        n14002) );
  OAI222XL U47922 ( .A0(net266570), .A1(n42276), .B0(n40164), .B1(n42277),
        .C0(n40286), .C1(n42278), .Y(n14004) );
  OAI211X1 U47923 ( .A0(n42280), .A1(n42868), .B0(n13978), .C0(n49997), .Y(
        n34832) );
  OA22X1 U47924 ( .A0(net263007), .A1(n42282), .B0(n42281), .B1(n40096), .Y(
        n13978) );
  OAI222XL U47925 ( .A0(net266570), .A1(n42277), .B0(n40164), .B1(n42278),
        .C0(net217178), .C1(n42279), .Y(n13980) );
  OAI211X1 U47926 ( .A0(n42281), .A1(n42869), .B0(n13954), .C0(n49999), .Y(
        n34824) );
  OA22X1 U47927 ( .A0(net263007), .A1(n42283), .B0(n42282), .B1(n40095), .Y(
        n13954) );
  OAI222XL U47928 ( .A0(net266570), .A1(n42278), .B0(n40164), .B1(n42279),
        .C0(net217178), .C1(n42280), .Y(n13956) );
  OAI211X1 U47929 ( .A0(n42282), .A1(n42870), .B0(n13930), .C0(n50001), .Y(
        n34816) );
  OA22X1 U47930 ( .A0(net263026), .A1(n42284), .B0(n42283), .B1(n40095), .Y(
        n13930) );
  OAI222XL U47931 ( .A0(net266570), .A1(n42279), .B0(n40164), .B1(n42280),
        .C0(net217178), .C1(n42281), .Y(n13932) );
  OAI211X1 U47932 ( .A0(n42283), .A1(n42872), .B0(n13906), .C0(n50003), .Y(
        n34808) );
  OA22X1 U47933 ( .A0(net263026), .A1(n42285), .B0(n42284), .B1(n40094), .Y(
        n13906) );
  OAI222XL U47934 ( .A0(net266570), .A1(n42280), .B0(n40164), .B1(n42281),
        .C0(net217178), .C1(n42282), .Y(n13908) );
  OAI211X1 U47935 ( .A0(n42284), .A1(n42873), .B0(n13882), .C0(n50005), .Y(
        n34800) );
  OA22X1 U47936 ( .A0(net263026), .A1(n42286), .B0(n42285), .B1(n40094), .Y(
        n13882) );
  OAI222XL U47937 ( .A0(net266570), .A1(n42281), .B0(n40164), .B1(n42282),
        .C0(net217178), .C1(n42283), .Y(n13884) );
  OAI211X1 U47938 ( .A0(n42285), .A1(n42874), .B0(n13858), .C0(n50007), .Y(
        n34792) );
  OA22X1 U47939 ( .A0(net263045), .A1(n42287), .B0(n42286), .B1(n40093), .Y(
        n13858) );
  OAI222XL U47940 ( .A0(net266591), .A1(n42282), .B0(n40163), .B1(n42283),
        .C0(net217178), .C1(n42284), .Y(n13860) );
  OAI211X1 U47941 ( .A0(n42286), .A1(n42875), .B0(n13834), .C0(n50009), .Y(
        n34784) );
  OA22X1 U47942 ( .A0(net263045), .A1(n42288), .B0(n42287), .B1(n40093), .Y(
        n13834) );
  OAI222XL U47943 ( .A0(net266591), .A1(n42283), .B0(n40163), .B1(n42284),
        .C0(net217178), .C1(n42285), .Y(n13836) );
  OAI211X1 U47944 ( .A0(n42287), .A1(n42876), .B0(n13810), .C0(n50011), .Y(
        n34776) );
  OA22X1 U47945 ( .A0(net263064), .A1(n42289), .B0(n42288), .B1(n40092), .Y(
        n13810) );
  OAI222XL U47946 ( .A0(net266591), .A1(n42284), .B0(n40163), .B1(n42285),
        .C0(net217178), .C1(n42286), .Y(n13812) );
  OAI211X1 U47947 ( .A0(n42288), .A1(n42877), .B0(n13786), .C0(n50013), .Y(
        n34768) );
  OA22X1 U47948 ( .A0(net263330), .A1(n42290), .B0(n42289), .B1(n40077), .Y(
        n13786) );
  OAI222XL U47949 ( .A0(net266591), .A1(n42285), .B0(n40163), .B1(n42286),
        .C0(n40289), .C1(n42287), .Y(n13788) );
  OAI211X1 U47950 ( .A0(n42289), .A1(n42878), .B0(n13762), .C0(n50015), .Y(
        n34760) );
  OA22X1 U47951 ( .A0(net263349), .A1(n42291), .B0(n42290), .B1(n40076), .Y(
        n13762) );
  OAI222XL U47952 ( .A0(net266591), .A1(n42286), .B0(n40163), .B1(n42287),
        .C0(n40289), .C1(n42288), .Y(n13764) );
  OAI211X1 U47953 ( .A0(n42290), .A1(n42912), .B0(n13738), .C0(n50017), .Y(
        n34752) );
  OA22X1 U47954 ( .A0(net263349), .A1(n42292), .B0(n42291), .B1(n40076), .Y(
        n13738) );
  OAI222XL U47955 ( .A0(net266591), .A1(n42287), .B0(n40163), .B1(n42288),
        .C0(n40289), .C1(n42289), .Y(n13740) );
  OAI211X1 U47956 ( .A0(n42291), .A1(n42913), .B0(n13714), .C0(n50019), .Y(
        n34744) );
  OA22X1 U47957 ( .A0(net263368), .A1(n42293), .B0(n42292), .B1(n40075), .Y(
        n13714) );
  OAI222XL U47958 ( .A0(net266591), .A1(n42288), .B0(n40163), .B1(n42289),
        .C0(n40289), .C1(n42290), .Y(n13716) );
  OAI211X1 U47959 ( .A0(n42292), .A1(n42914), .B0(n13690), .C0(n50021), .Y(
        n34736) );
  OA22X1 U47960 ( .A0(net263368), .A1(n42294), .B0(n42293), .B1(n40075), .Y(
        n13690) );
  OAI222XL U47961 ( .A0(net266591), .A1(n42289), .B0(n40163), .B1(n42290),
        .C0(n40289), .C1(n42291), .Y(n13692) );
  OAI211X1 U47962 ( .A0(n42293), .A1(n42915), .B0(n13666), .C0(n50023), .Y(
        n34728) );
  OA22X1 U47963 ( .A0(net263387), .A1(n42295), .B0(n42294), .B1(n40074), .Y(
        n13666) );
  OAI222XL U47964 ( .A0(net266591), .A1(n42290), .B0(n40163), .B1(n42291),
        .C0(n40289), .C1(n42292), .Y(n13668) );
  OAI211X1 U47965 ( .A0(n42294), .A1(n42916), .B0(n13642), .C0(n50025), .Y(
        n34720) );
  OA22X1 U47966 ( .A0(net263387), .A1(n42296), .B0(n42295), .B1(n40074), .Y(
        n13642) );
  OAI222XL U47967 ( .A0(net266591), .A1(n42291), .B0(n40162), .B1(n42292),
        .C0(n40289), .C1(n42293), .Y(n13644) );
  OAI211X1 U47968 ( .A0(n42295), .A1(n42917), .B0(n13618), .C0(n50027), .Y(
        n34712) );
  OA22X1 U47969 ( .A0(net263387), .A1(n42297), .B0(n42296), .B1(n40073), .Y(
        n13618) );
  OAI222XL U47970 ( .A0(net266612), .A1(n42292), .B0(n40162), .B1(n42293),
        .C0(n40289), .C1(n42294), .Y(n13620) );
  OAI211X1 U47971 ( .A0(n42296), .A1(n42918), .B0(n13594), .C0(n50029), .Y(
        n34704) );
  OA22X1 U47972 ( .A0(net263406), .A1(n42298), .B0(n42297), .B1(n40073), .Y(
        n13594) );
  OAI222XL U47973 ( .A0(net266612), .A1(n42293), .B0(n40162), .B1(n42294),
        .C0(n40290), .C1(n42295), .Y(n13596) );
  OAI211X1 U47974 ( .A0(n42297), .A1(n42920), .B0(n13570), .C0(n50031), .Y(
        n34696) );
  OA22X1 U47975 ( .A0(net263406), .A1(n42299), .B0(n42298), .B1(n40072), .Y(
        n13570) );
  OAI222XL U47976 ( .A0(net266612), .A1(n42294), .B0(n40162), .B1(n42295),
        .C0(n40290), .C1(n42296), .Y(n13572) );
  OAI211X1 U47977 ( .A0(n42298), .A1(n42921), .B0(n13546), .C0(n50033), .Y(
        n34688) );
  OA22X1 U47978 ( .A0(net218304), .A1(n42300), .B0(n42299), .B1(n40072), .Y(
        n13546) );
  OAI222XL U47979 ( .A0(net266612), .A1(n42295), .B0(n40162), .B1(n42296),
        .C0(n40290), .C1(n42297), .Y(n13548) );
  OAI211X1 U47980 ( .A0(n42299), .A1(n42922), .B0(n13522), .C0(n50035), .Y(
        n34680) );
  OA22X1 U47981 ( .A0(net218302), .A1(n42301), .B0(n42300), .B1(n40071), .Y(
        n13522) );
  OAI222XL U47982 ( .A0(net266612), .A1(n42296), .B0(n40162), .B1(n42297),
        .C0(n40290), .C1(n42298), .Y(n13524) );
  OAI211X1 U47983 ( .A0(n42300), .A1(n42923), .B0(n13498), .C0(n50037), .Y(
        n34672) );
  OA22X1 U47984 ( .A0(net263444), .A1(n42302), .B0(n42301), .B1(n40071), .Y(
        n13498) );
  OAI222XL U47985 ( .A0(net266612), .A1(n42297), .B0(n40162), .B1(n42298),
        .C0(n40290), .C1(n42299), .Y(n13500) );
  OAI211X1 U47986 ( .A0(n42301), .A1(n42924), .B0(n13474), .C0(n50039), .Y(
        n34664) );
  OA22X1 U47987 ( .A0(net263444), .A1(n42303), .B0(n42302), .B1(n40070), .Y(
        n13474) );
  OAI222XL U47988 ( .A0(net266612), .A1(n42298), .B0(n40162), .B1(n42299),
        .C0(n40290), .C1(n42300), .Y(n13476) );
  OAI211X1 U47989 ( .A0(n42302), .A1(n42925), .B0(n13450), .C0(n50041), .Y(
        n34656) );
  OA22X1 U47990 ( .A0(net263463), .A1(n42304), .B0(n42303), .B1(n40070), .Y(
        n13450) );
  OAI222XL U47991 ( .A0(net266612), .A1(n42299), .B0(n40161), .B1(n42300),
        .C0(n40290), .C1(n42301), .Y(n13452) );
  OAI211X1 U47992 ( .A0(n42303), .A1(n42927), .B0(n13426), .C0(n50043), .Y(
        n34648) );
  OA22X1 U47993 ( .A0(net263463), .A1(n42305), .B0(n42304), .B1(n40069), .Y(
        n13426) );
  OAI222XL U47994 ( .A0(net266612), .A1(n42300), .B0(n40161), .B1(n42301),
        .C0(n40290), .C1(n42302), .Y(n13428) );
  OAI211X1 U47995 ( .A0(n42304), .A1(n42895), .B0(n13402), .C0(n50045), .Y(
        n34640) );
  OA22X1 U47996 ( .A0(net218426), .A1(n42306), .B0(n42305), .B1(n40084), .Y(
        n13402) );
  OAI222XL U47997 ( .A0(net266612), .A1(n42301), .B0(n40161), .B1(n42302),
        .C0(n40290), .C1(n42303), .Y(n13404) );
  OAI211X1 U47998 ( .A0(n42305), .A1(n42897), .B0(n13378), .C0(n50047), .Y(
        n34632) );
  OA22X1 U47999 ( .A0(net263216), .A1(n42307), .B0(n42306), .B1(n40083), .Y(
        n13378) );
  OAI222XL U48000 ( .A0(net266633), .A1(n42302), .B0(n40161), .B1(n42303),
        .C0(n40291), .C1(n42304), .Y(n13380) );
  OAI211X1 U48001 ( .A0(n42306), .A1(n42898), .B0(n13354), .C0(n50049), .Y(
        n34624) );
  OA22X1 U48002 ( .A0(net263216), .A1(n42308), .B0(n42307), .B1(n40083), .Y(
        n13354) );
  OAI222XL U48003 ( .A0(net266633), .A1(n42303), .B0(n40161), .B1(n42304),
        .C0(n40291), .C1(n42305), .Y(n13356) );
  OAI211X1 U48004 ( .A0(n42307), .A1(n42899), .B0(n13330), .C0(n50051), .Y(
        n34616) );
  OA22X1 U48005 ( .A0(net263235), .A1(n42309), .B0(n42308), .B1(n40082), .Y(
        n13330) );
  OAI222XL U48006 ( .A0(net266633), .A1(n42304), .B0(n40161), .B1(n42305),
        .C0(n40291), .C1(n42306), .Y(n13332) );
  OAI211X1 U48007 ( .A0(n42308), .A1(n42900), .B0(n13306), .C0(n50053), .Y(
        n34608) );
  OA22X1 U48008 ( .A0(net263235), .A1(n42310), .B0(n42309), .B1(n40082), .Y(
        n13306) );
  OAI222XL U48009 ( .A0(net266633), .A1(n42305), .B0(n40161), .B1(n42306),
        .C0(n40291), .C1(n42307), .Y(n13308) );
  OAI211X1 U48010 ( .A0(n42309), .A1(n42901), .B0(n13282), .C0(n50055), .Y(
        n34600) );
  OA22X1 U48011 ( .A0(net263254), .A1(n42311), .B0(n42310), .B1(n40081), .Y(
        n13282) );
  OAI222XL U48012 ( .A0(net266633), .A1(n42306), .B0(n40161), .B1(n42307),
        .C0(n40291), .C1(n42308), .Y(n13284) );
  OAI211X1 U48013 ( .A0(n42310), .A1(n42902), .B0(n13258), .C0(n50057), .Y(
        n34592) );
  OA22X1 U48014 ( .A0(net263254), .A1(n42312), .B0(n42311), .B1(n40081), .Y(
        n13258) );
  OAI222XL U48015 ( .A0(net266633), .A1(n42307), .B0(n40161), .B1(n42308),
        .C0(n40291), .C1(n42309), .Y(n13260) );
  OAI211X1 U48016 ( .A0(n42311), .A1(n42904), .B0(n13234), .C0(n50059), .Y(
        n34584) );
  OA22X1 U48017 ( .A0(net263254), .A1(n42313), .B0(n42312), .B1(n40080), .Y(
        n13234) );
  OAI222XL U48018 ( .A0(net266633), .A1(n42308), .B0(n40160), .B1(n42309),
        .C0(n40291), .C1(n42310), .Y(n13236) );
  OAI211X1 U48019 ( .A0(n42312), .A1(n42905), .B0(n13210), .C0(n50061), .Y(
        n34576) );
  OA22X1 U48020 ( .A0(net218310), .A1(n42314), .B0(n42313), .B1(n40080), .Y(
        n13210) );
  OAI222XL U48021 ( .A0(net266633), .A1(n42309), .B0(n40160), .B1(n42310),
        .C0(n40291), .C1(n42311), .Y(n13212) );
  OAI211X1 U48022 ( .A0(n42313), .A1(n42906), .B0(n13186), .C0(n50063), .Y(
        n34568) );
  OA22X1 U48023 ( .A0(net218312), .A1(n42315), .B0(n42314), .B1(n40079), .Y(
        n13186) );
  OAI222XL U48024 ( .A0(net266633), .A1(n42310), .B0(n40160), .B1(n42311),
        .C0(n40291), .C1(n42312), .Y(n13188) );
  OAI211X1 U48025 ( .A0(n42314), .A1(n42907), .B0(n13162), .C0(n50065), .Y(
        n34560) );
  OA22X1 U48026 ( .A0(net263292), .A1(n36883), .B0(n42315), .B1(n40079), .Y(
        n13162) );
  OAI211X1 U48027 ( .A0(n42315), .A1(n42908), .B0(n13138), .C0(n50067), .Y(
        n34552) );
  OAI222XL U48028 ( .A0(net266654), .A1(n42312), .B0(n40160), .B1(n42313),
        .C0(n40292), .C1(n42314), .Y(n13140) );
  OAI222XL U48029 ( .A0(net266654), .A1(n42313), .B0(n40160), .B1(n42314),
        .C0(n40292), .C1(n42315), .Y(n13116) );
  OAI222XL U48030 ( .A0(net266654), .A1(n42314), .B0(n40160), .B1(n42315),
        .C0(n40292), .C1(n36880), .Y(n13092) );
  OAI222XL U48031 ( .A0(net266654), .A1(n42315), .B0(n40160), .B1(n36879),
        .C0(n40292), .C1(n42663), .Y(n13062) );
  NAND4BX1 U48032 ( .AN(n9991), .B(n9993), .C(n9992), .D(n20792), .Y(n9876) );
  AND3X2 U48033 ( .A(n10631), .B(n10630), .C(n10629), .Y(n20792) );
  OA22X1 U48034 ( .A0(net262285), .A1(n42165), .B0(n42164), .B1(n40078), .Y(
        n16786) );
  CLKINVX1 U48035 ( .A(n16788), .Y(n49763) );
  OAI222XL U48036 ( .A0(net266318), .A1(n42160), .B0(n40178), .B1(n42161),
        .C0(net217272), .C1(n42162), .Y(n16788) );
  NOR2X1 U48037 ( .A(n10819), .B(n10821), .Y(n22796) );
  XNOR2X1 U48038 ( .A(n50860), .B(n41290), .Y(n24412) );
  XNOR2X1 U48039 ( .A(n50867), .B(n42536), .Y(n30597) );
  XNOR2X1 U48040 ( .A(n50864), .B(n42537), .Y(n30477) );
  XNOR2X1 U48041 ( .A(n50861), .B(n42541), .Y(n30567) );
  XNOR2X1 U48042 ( .A(n50860), .B(n42535), .Y(n30295) );
  XNOR2X1 U48043 ( .A(n50862), .B(n42535), .Y(n30537) );
  XNOR2X1 U48044 ( .A(n50857), .B(n42542), .Y(n30235) );
  XNOR2X1 U48045 ( .A(n50858), .B(n42536), .Y(n30205) );
  XNOR2X1 U48046 ( .A(n50863), .B(n42539), .Y(n30447) );
  XNOR2X1 U48047 ( .A(n50866), .B(n42542), .Y(n30627) );
  XNOR2X1 U48048 ( .A(n50859), .B(n42535), .Y(n30265) );
  XNOR2X1 U48049 ( .A(n50856), .B(n42542), .Y(n30385) );
  XNOR2X1 U48050 ( .A(n50855), .B(n42543), .Y(n30415) );
  XNOR2X1 U48051 ( .A(n51298), .B(n42697), .Y(n30531) );
  XNOR2X1 U48052 ( .A(n51297), .B(n42697), .Y(n30621) );
  XNOR2X1 U48053 ( .A(n51288), .B(n42694), .Y(n30229) );
  XNOR2X1 U48054 ( .A(n51282), .B(n42694), .Y(n30138) );
  XNOR2X1 U48055 ( .A(n51279), .B(n42694), .Y(n30198) );
  XNOR2X1 U48056 ( .A(n51278), .B(n42694), .Y(n30078) );
  XNOR2X1 U48057 ( .A(n51277), .B(n42694), .Y(n30048) );
  XNOR2X1 U48058 ( .A(n51276), .B(n42694), .Y(n30018) );
  XNOR2X1 U48059 ( .A(n51281), .B(n42694), .Y(n30108) );
  XNOR2X1 U48060 ( .A(n51280), .B(n42694), .Y(n30168) );
  XNOR2X1 U48061 ( .A(n51267), .B(n42694), .Y(n29928) );
  XNOR2X1 U48062 ( .A(n51268), .B(n42694), .Y(n29868) );
  XNOR2X1 U48063 ( .A(n51275), .B(n42694), .Y(n29988) );
  XNOR2X1 U48064 ( .A(n51272), .B(n42694), .Y(n29838) );
  XNOR2X1 U48065 ( .A(n51269), .B(n42694), .Y(n29898) );
  XNOR2X1 U48066 ( .A(n51074), .B(n41328), .Y(n24413) );
  XNOR2X1 U48067 ( .A(n51297), .B(n42639), .Y(n30523) );
  XNOR2X1 U48068 ( .A(n50655), .B(n42587), .Y(n30519) );
  XNOR2X1 U48069 ( .A(n50654), .B(n42587), .Y(n30609) );
  XNOR2X1 U48070 ( .A(n51081), .B(n42552), .Y(n30598) );
  XNOR2X1 U48071 ( .A(n51078), .B(n42551), .Y(n30478) );
  XNOR2X1 U48072 ( .A(n51075), .B(n42552), .Y(n30568) );
  XNOR2X1 U48073 ( .A(n51074), .B(n36832), .Y(n30296) );
  XNOR2X1 U48074 ( .A(n51076), .B(n42549), .Y(n30538) );
  XNOR2X1 U48075 ( .A(n51071), .B(n36832), .Y(n30236) );
  XNOR2X1 U48076 ( .A(n51072), .B(n42552), .Y(n30206) );
  XNOR2X1 U48077 ( .A(n51278), .B(n36867), .Y(n30190) );
  XNOR2X1 U48078 ( .A(n51276), .B(n36867), .Y(n30040) );
  XNOR2X1 U48079 ( .A(n50634), .B(n42587), .Y(n30036) );
  XNOR2X1 U48080 ( .A(n51275), .B(n36867), .Y(n30010) );
  XNOR2X1 U48081 ( .A(n50633), .B(n42587), .Y(n30006) );
  XNOR2X1 U48082 ( .A(n51279), .B(n36867), .Y(n30160) );
  XNOR2X1 U48083 ( .A(n50637), .B(n42587), .Y(n30156) );
  XNOR2X1 U48084 ( .A(n51077), .B(n42552), .Y(n30448) );
  XNOR2X1 U48085 ( .A(n51073), .B(n42552), .Y(n30266) );
  XNOR2X1 U48086 ( .A(n51266), .B(n36867), .Y(n29920) );
  XNOR2X1 U48087 ( .A(n50624), .B(n42587), .Y(n29916) );
  XNOR2X1 U48088 ( .A(n51274), .B(n36867), .Y(n29980) );
  XNOR2X1 U48089 ( .A(n50632), .B(n42587), .Y(n29976) );
  XNOR2X1 U48090 ( .A(n51271), .B(n36867), .Y(n29830) );
  XNOR2X1 U48091 ( .A(n50629), .B(n42587), .Y(n29826) );
  XNOR2X1 U48092 ( .A(n50615), .B(net219434), .Y(n26133) );
  XNOR2X1 U48093 ( .A(n51070), .B(n36832), .Y(n30386) );
  XNOR2X1 U48094 ( .A(n51069), .B(n42552), .Y(n30416) );
  XNOR2X1 U48095 ( .A(n50614), .B(net219434), .Y(n26103) );
  XNOR2X1 U48096 ( .A(n50606), .B(net258207), .Y(n25923) );
  XNOR2X1 U48097 ( .A(n50434), .B(n42717), .Y(n30197) );
  XNOR2X1 U48098 ( .A(n50432), .B(n42724), .Y(n30047) );
  XNOR2X1 U48099 ( .A(n50431), .B(n42719), .Y(n30017) );
  XNOR2X1 U48100 ( .A(n50436), .B(n36875), .Y(n30107) );
  XNOR2X1 U48101 ( .A(n50435), .B(n42719), .Y(n30167) );
  XNOR2X1 U48102 ( .A(n50422), .B(n36875), .Y(n29927) );
  XNOR2X1 U48103 ( .A(n50430), .B(n36875), .Y(n29987) );
  XNOR2X1 U48104 ( .A(n50427), .B(n42724), .Y(n29837) );
  XNOR2X1 U48105 ( .A(n50646), .B(n36854), .Y(n24414) );
  XNOR2X1 U48106 ( .A(n50238), .B(n42706), .Y(n30529) );
  XNOR2X1 U48107 ( .A(n50237), .B(n42671), .Y(n30521) );
  XNOR2X1 U48108 ( .A(n50869), .B(n42616), .Y(n30517) );
  XNOR2X1 U48109 ( .A(n50236), .B(n42671), .Y(n30611) );
  XNOR2X1 U48110 ( .A(n50868), .B(n42616), .Y(n30607) );
  XNOR2X1 U48111 ( .A(n50219), .B(n42704), .Y(n30196) );
  XNOR2X1 U48112 ( .A(n50217), .B(n42712), .Y(n30046) );
  XNOR2X1 U48113 ( .A(n50216), .B(n42675), .Y(n30038) );
  XNOR2X1 U48114 ( .A(n50848), .B(n42615), .Y(n30034) );
  XNOR2X1 U48115 ( .A(n50216), .B(n42707), .Y(n30016) );
  XNOR2X1 U48116 ( .A(n50215), .B(n42675), .Y(n30008) );
  XNOR2X1 U48117 ( .A(n50847), .B(n42619), .Y(n30004) );
  XNOR2X1 U48118 ( .A(n50220), .B(n41642), .Y(n30166) );
  XNOR2X1 U48119 ( .A(n50219), .B(n42675), .Y(n30158) );
  XNOR2X1 U48120 ( .A(n50207), .B(n42711), .Y(n29926) );
  XNOR2X1 U48121 ( .A(n50206), .B(n42675), .Y(n29918) );
  XNOR2X1 U48122 ( .A(n50838), .B(n42616), .Y(n29914) );
  XNOR2X1 U48123 ( .A(n50215), .B(n41641), .Y(n29986) );
  XNOR2X1 U48124 ( .A(n50214), .B(n42675), .Y(n29978) );
  XNOR2X1 U48125 ( .A(n50846), .B(n42615), .Y(n29974) );
  XNOR2X1 U48126 ( .A(n50212), .B(n42711), .Y(n29836) );
  XNOR2X1 U48127 ( .A(n50211), .B(n42675), .Y(n29828) );
  XNOR2X1 U48128 ( .A(n50843), .B(n42615), .Y(n29824) );
  XNOR2X1 U48129 ( .A(n50452), .B(n36834), .Y(n30522) );
  XNOR2X1 U48130 ( .A(n51083), .B(n42625), .Y(n30518) );
  XNOR2X1 U48131 ( .A(n50451), .B(n41379), .Y(n30612) );
  XNOR2X1 U48132 ( .A(n51082), .B(n42624), .Y(n30608) );
  XNOR2X1 U48133 ( .A(n50646), .B(n42503), .Y(n30297) );
  XNOR2X1 U48134 ( .A(n50643), .B(n36731), .Y(n30237) );
  XNOR2X1 U48135 ( .A(n50644), .B(n42504), .Y(n30207) );
  XNOR2X1 U48136 ( .A(n50431), .B(n36903), .Y(n30039) );
  XNOR2X1 U48137 ( .A(n51062), .B(n42633), .Y(n30035) );
  XNOR2X1 U48138 ( .A(n50430), .B(n36903), .Y(n30009) );
  XNOR2X1 U48139 ( .A(n51061), .B(n42628), .Y(n30005) );
  XNOR2X1 U48140 ( .A(n50434), .B(n36834), .Y(n30159) );
  XNOR2X1 U48141 ( .A(n51065), .B(n42627), .Y(n30155) );
  XNOR2X1 U48142 ( .A(n50645), .B(n42503), .Y(n30267) );
  XNOR2X1 U48143 ( .A(n50421), .B(n36903), .Y(n29919) );
  XNOR2X1 U48144 ( .A(n51052), .B(n42625), .Y(n29915) );
  XNOR2X1 U48145 ( .A(n50429), .B(n36903), .Y(n29979) );
  XNOR2X1 U48146 ( .A(n51060), .B(n42626), .Y(n29975) );
  XNOR2X1 U48147 ( .A(n50426), .B(n36903), .Y(n29829) );
  XNOR2X1 U48148 ( .A(n51057), .B(n34447), .Y(n29825) );
  XOR2X1 U48149 ( .A(n41994), .B(n36892), .Y(n30256) );
  XOR2X1 U48150 ( .A(n42253), .B(n36879), .Y(n30260) );
  XOR2X1 U48151 ( .A(n42254), .B(n42654), .Y(n30252) );
  XOR2X1 U48152 ( .A(n41995), .B(n36711), .Y(n30248) );
  XOR2X1 U48153 ( .A(n41993), .B(n36901), .Y(n30226) );
  XOR2X1 U48154 ( .A(n42252), .B(n36886), .Y(n30230) );
  XOR2X1 U48155 ( .A(n42253), .B(n42654), .Y(n30222) );
  XOR2X1 U48156 ( .A(n41994), .B(n36711), .Y(n30218) );
  XOR2X1 U48157 ( .A(n41999), .B(n36901), .Y(n30135) );
  XOR2X1 U48158 ( .A(n42258), .B(n36879), .Y(n30139) );
  XOR2X1 U48159 ( .A(n42259), .B(n42654), .Y(n30131) );
  XOR2X1 U48160 ( .A(n42000), .B(n36711), .Y(n30127) );
  XOR2X1 U48161 ( .A(n42002), .B(n36898), .Y(n30195) );
  XOR2X1 U48162 ( .A(n42261), .B(n36885), .Y(n30199) );
  XOR2X1 U48163 ( .A(n42262), .B(n42654), .Y(n30191) );
  XOR2X1 U48164 ( .A(n42003), .B(n36711), .Y(n30187) );
  XOR2X1 U48165 ( .A(n42003), .B(n36894), .Y(n30075) );
  XOR2X1 U48166 ( .A(n42262), .B(n36883), .Y(n30079) );
  XOR2X1 U48167 ( .A(n42004), .B(n36894), .Y(n30045) );
  XOR2X1 U48168 ( .A(n42263), .B(n36885), .Y(n30049) );
  XOR2X1 U48169 ( .A(n42264), .B(n42654), .Y(n30041) );
  XOR2X1 U48170 ( .A(n42005), .B(n36711), .Y(n30037) );
  XOR2X1 U48171 ( .A(n42005), .B(n36897), .Y(n30015) );
  XOR2X1 U48172 ( .A(n42264), .B(n36889), .Y(n30019) );
  XOR2X1 U48173 ( .A(n42265), .B(n42654), .Y(n30011) );
  XOR2X1 U48174 ( .A(n42006), .B(n36711), .Y(n30007) );
  XOR2X1 U48175 ( .A(n42000), .B(n36901), .Y(n30105) );
  XOR2X1 U48176 ( .A(n42259), .B(n36886), .Y(n30109) );
  XOR2X1 U48177 ( .A(n42260), .B(n42654), .Y(n30101) );
  XOR2X1 U48178 ( .A(n42001), .B(n36711), .Y(n30097) );
  XOR2X1 U48179 ( .A(n42010), .B(n36894), .Y(n29805) );
  XOR2X1 U48180 ( .A(n42269), .B(n36881), .Y(n29809) );
  XOR2X1 U48181 ( .A(n42001), .B(n36900), .Y(n30165) );
  XOR2X1 U48182 ( .A(n42260), .B(n36879), .Y(n30169) );
  XOR2X1 U48183 ( .A(n42261), .B(n42654), .Y(n30161) );
  XOR2X1 U48184 ( .A(n42002), .B(n36711), .Y(n30157) );
  XOR2X1 U48185 ( .A(n42011), .B(n36899), .Y(n29955) );
  XOR2X1 U48186 ( .A(n42270), .B(n36885), .Y(n29959) );
  XOR2X1 U48187 ( .A(n42019), .B(n36893), .Y(n29624) );
  XOR2X1 U48188 ( .A(n42278), .B(n36882), .Y(n29628) );
  XOR2X1 U48189 ( .A(n42014), .B(n36898), .Y(n29925) );
  XOR2X1 U48190 ( .A(n42273), .B(n36889), .Y(n29929) );
  XOR2X1 U48191 ( .A(n42274), .B(n42661), .Y(n29921) );
  XOR2X1 U48192 ( .A(n42015), .B(n42602), .Y(n29917) );
  XOR2X1 U48193 ( .A(n41997), .B(n36894), .Y(n30346) );
  XOR2X1 U48194 ( .A(n42256), .B(n36888), .Y(n30350) );
  XOR2X1 U48195 ( .A(n42257), .B(n42654), .Y(n30342) );
  XOR2X1 U48196 ( .A(n41998), .B(n36711), .Y(n30338) );
  XOR2X1 U48197 ( .A(n42013), .B(n36895), .Y(n29865) );
  XOR2X1 U48198 ( .A(n42272), .B(n36889), .Y(n29869) );
  XOR2X1 U48199 ( .A(n42273), .B(n42648), .Y(n29861) );
  XOR2X1 U48200 ( .A(n42282), .B(n36888), .Y(n26168) );
  XOR2X1 U48201 ( .A(n42258), .B(n42654), .Y(n30372) );
  XOR2X1 U48202 ( .A(n41999), .B(n36711), .Y(n30368) );
  XOR2X1 U48203 ( .A(n42285), .B(n36887), .Y(n26078) );
  XOR2X1 U48204 ( .A(n42288), .B(n36888), .Y(n26018) );
  XOR2X1 U48205 ( .A(n42007), .B(n36898), .Y(n29775) );
  XOR2X1 U48206 ( .A(n42266), .B(n36889), .Y(n29779) );
  XOR2X1 U48207 ( .A(n42267), .B(n42665), .Y(n29771) );
  XOR2X1 U48208 ( .A(n42008), .B(n42602), .Y(n29767) );
  XOR2X1 U48209 ( .A(n42006), .B(n36891), .Y(n29985) );
  XOR2X1 U48210 ( .A(n42265), .B(n36888), .Y(n29989) );
  XOR2X1 U48211 ( .A(n42266), .B(n42665), .Y(n29981) );
  XOR2X1 U48212 ( .A(n42007), .B(n42602), .Y(n29977) );
  XOR2X1 U48213 ( .A(n42008), .B(n36895), .Y(n29745) );
  XOR2X1 U48214 ( .A(n42267), .B(n36889), .Y(n29749) );
  XOR2X1 U48215 ( .A(n42268), .B(n42664), .Y(n29741) );
  XOR2X1 U48216 ( .A(n42009), .B(n42602), .Y(n29737) );
  XOR2X1 U48217 ( .A(n42009), .B(n36894), .Y(n29835) );
  XOR2X1 U48218 ( .A(n42268), .B(n36881), .Y(n29839) );
  XOR2X1 U48219 ( .A(n42269), .B(n42652), .Y(n29831) );
  XOR2X1 U48220 ( .A(n42010), .B(n42602), .Y(n29827) );
  XOR2X1 U48221 ( .A(n42012), .B(n36899), .Y(n29895) );
  XOR2X1 U48222 ( .A(n42271), .B(n36880), .Y(n29899) );
  XOR2X1 U48223 ( .A(n42287), .B(n36883), .Y(n25988) );
  XOR2X1 U48224 ( .A(n42289), .B(n36887), .Y(n26048) );
  XOR2X1 U48225 ( .A(n42015), .B(n36894), .Y(n29594) );
  XOR2X1 U48226 ( .A(n42274), .B(n36885), .Y(n29598) );
  XOR2X1 U48227 ( .A(n42283), .B(n36885), .Y(n26138) );
  XOR2X1 U48228 ( .A(n42024), .B(n36893), .Y(n26134) );
  XOR2X1 U48229 ( .A(n42284), .B(n42654), .Y(n26130) );
  XOR2X1 U48230 ( .A(n42025), .B(n42606), .Y(n26126) );
  XOR2X1 U48231 ( .A(n42020), .B(n36900), .Y(n29654) );
  XOR2X1 U48232 ( .A(n42279), .B(n36882), .Y(n29658) );
  XOR2X1 U48233 ( .A(n42280), .B(n42655), .Y(n29650) );
  XOR2X1 U48234 ( .A(n42021), .B(n42602), .Y(n29646) );
  XOR2X1 U48235 ( .A(n42021), .B(n36891), .Y(n29684) );
  XOR2X1 U48236 ( .A(n42280), .B(n36880), .Y(n29688) );
  XOR2X1 U48237 ( .A(n42284), .B(n36879), .Y(n26108) );
  XOR2X1 U48238 ( .A(n42025), .B(n36892), .Y(n26104) );
  XOR2X1 U48239 ( .A(n42285), .B(n42653), .Y(n26100) );
  XOR2X1 U48240 ( .A(n42026), .B(n42606), .Y(n26096) );
  XOR2X1 U48241 ( .A(n42022), .B(n36893), .Y(n29714) );
  XOR2X1 U48242 ( .A(n42281), .B(n36887), .Y(n29718) );
  XOR2X1 U48243 ( .A(n42282), .B(n42652), .Y(n29710) );
  XOR2X1 U48244 ( .A(n42023), .B(n42602), .Y(n29706) );
  XOR2X1 U48245 ( .A(n41991), .B(n36893), .Y(n30316) );
  XOR2X1 U48246 ( .A(n42250), .B(n36881), .Y(n30320) );
  XOR2X1 U48247 ( .A(n42251), .B(n42654), .Y(n30312) );
  XOR2X1 U48248 ( .A(n41992), .B(n36711), .Y(n30308) );
  XOR2X1 U48249 ( .A(n42301), .B(n36889), .Y(n26198) );
  XOR2X1 U48250 ( .A(n42298), .B(n36881), .Y(n26288) );
  XOR2X1 U48251 ( .A(n42292), .B(n36887), .Y(n25928) );
  XOR2X1 U48252 ( .A(n42033), .B(n36891), .Y(n25924) );
  XOR2X1 U48253 ( .A(n42293), .B(n42654), .Y(n25920) );
  XOR2X1 U48254 ( .A(n42034), .B(n42606), .Y(n25916) );
  XOR2X1 U48255 ( .A(n42300), .B(n36879), .Y(n26228) );
  XOR2X1 U48256 ( .A(n42299), .B(n36888), .Y(n26258) );
  XOR2X1 U48257 ( .A(n41992), .B(n36901), .Y(n30286) );
  XOR2X1 U48258 ( .A(n42251), .B(n36883), .Y(n30290) );
  XOR2X1 U48259 ( .A(n42252), .B(n42654), .Y(n30282) );
  XOR2X1 U48260 ( .A(n41993), .B(n36711), .Y(n30278) );
  XOR2X1 U48261 ( .A(n41993), .B(n41318), .Y(n24415) );
  XOR2X1 U48262 ( .A(n41996), .B(n42515), .Y(n30238) );
  XOR2X1 U48263 ( .A(n41995), .B(n42515), .Y(n30208) );
  XOR2X1 U48264 ( .A(n42008), .B(n42515), .Y(n29967) );
  XOR2X1 U48265 ( .A(n42006), .B(n42515), .Y(n30027) );
  XOR2X1 U48266 ( .A(n42009), .B(n42518), .Y(n29757) );
  AND4X1 U48267 ( .A(n10007), .B(n36926), .C(net151440), .D(n10010), .Y(n10006) );
  AOI31X1 U48268 ( .A0(n50088), .A1(n10015), .A2(n10016), .B0(n9884), .Y(
        n10011) );
  CLKINVX1 U48269 ( .A(n10017), .Y(n50088) );
  NAND4X1 U48270 ( .A(n10968), .B(n10969), .C(n10965), .D(n10966), .Y(n10218)
         );
  XNOR2X1 U48271 ( .A(n50451), .B(n42576), .Y(n30512) );
  XNOR2X1 U48272 ( .A(n50450), .B(n42582), .Y(n30602) );
  XNOR2X1 U48273 ( .A(n50447), .B(n42581), .Y(n30482) );
  XNOR2X1 U48274 ( .A(n50444), .B(n42582), .Y(n30572) );
  XNOR2X1 U48275 ( .A(n50445), .B(n42582), .Y(n30542) );
  XNOR2X1 U48276 ( .A(n50440), .B(n42577), .Y(n30240) );
  XNOR2X1 U48277 ( .A(n50446), .B(n42582), .Y(n30452) );
  XNOR2X1 U48278 ( .A(n50449), .B(n42584), .Y(n30632) );
  XNOR2X1 U48279 ( .A(n50442), .B(n42576), .Y(n30270) );
  XNOR2X1 U48280 ( .A(n50439), .B(n42584), .Y(n30390) );
  XOR2X1 U48281 ( .A(n42252), .B(n36807), .Y(n24416) );
  XOR2X1 U48282 ( .A(n42255), .B(n41321), .Y(n30239) );
  XOR2X1 U48283 ( .A(n42254), .B(n36801), .Y(n30209) );
  XOR2X1 U48284 ( .A(n42267), .B(n41321), .Y(n29968) );
  NOR4X1 U48285 ( .A(n10222), .B(n10223), .C(net171476), .D(n10225), .Y(n10220) );
  AOI211X1 U48286 ( .A0(n9863), .A1(n10226), .B0(n10227), .C0(n10228), .Y(
        n10225) );
  OAI31XL U48287 ( .A0(n10229), .A1(n10230), .A2(n10231), .B0(n50112), .Y(
        n10226) );
  NOR4X1 U48288 ( .A(n21343), .B(n21342), .C(n21341), .D(n21340), .Y(n46835)
         );
  NOR4X1 U48289 ( .A(n21363), .B(n21362), .C(n21361), .D(n21360), .Y(n46825)
         );
  NOR4X1 U48290 ( .A(n26075), .B(n26076), .C(n26077), .D(n26078), .Y(n44378)
         );
  XNOR2X1 U48291 ( .A(n50195), .B(n42711), .Y(n26075) );
  XNOR2X1 U48292 ( .A(n50410), .B(n42717), .Y(n26076) );
  XNOR2X1 U48293 ( .A(n51255), .B(n42700), .Y(n26077) );
  NOR4X1 U48294 ( .A(n26015), .B(n26016), .C(n26017), .D(n26018), .Y(net215050) );
  XNOR2X1 U48295 ( .A(n50192), .B(n42711), .Y(n26015) );
  XNOR2X1 U48296 ( .A(n50407), .B(n42717), .Y(n26016) );
  NOR4X1 U48297 ( .A(n25985), .B(n25986), .C(n25987), .D(n25988), .Y(net215041) );
  XNOR2X1 U48298 ( .A(n50193), .B(n42705), .Y(n25985) );
  XNOR2X1 U48299 ( .A(n50408), .B(n42723), .Y(n25986) );
  NOR4X1 U48300 ( .A(n26045), .B(n26046), .C(n26047), .D(n26048), .Y(net215059) );
  XNOR2X1 U48301 ( .A(n50191), .B(n42705), .Y(n26045) );
  XNOR2X1 U48302 ( .A(n50406), .B(n42725), .Y(n26046) );
  XNOR2X1 U48303 ( .A(n51251), .B(n41385), .Y(n26047) );
  NOR4X1 U48304 ( .A(n26195), .B(n26196), .C(n26197), .D(n26198), .Y(net214750) );
  XNOR2X1 U48305 ( .A(n50179), .B(n42706), .Y(n26195) );
  XNOR2X1 U48306 ( .A(n50394), .B(n41287), .Y(n26196) );
  XNOR2X1 U48307 ( .A(n51239), .B(n41385), .Y(n26197) );
  NOR4X1 U48308 ( .A(n25925), .B(n25926), .C(n25927), .D(n25928), .Y(net215005) );
  XNOR2X1 U48309 ( .A(n50188), .B(n41642), .Y(n25925) );
  XNOR2X1 U48310 ( .A(n50403), .B(n34435), .Y(n25926) );
  NOR4X1 U48311 ( .A(n25865), .B(n25866), .C(n25867), .D(n25868), .Y(net215023) );
  XNOR2X1 U48312 ( .A(n50189), .B(n42705), .Y(n25865) );
  XNOR2X1 U48313 ( .A(n50404), .B(n42719), .Y(n25866) );
  NOR4X1 U48314 ( .A(n26345), .B(n26346), .C(n26347), .D(n26348), .Y(net215131) );
  XNOR2X1 U48315 ( .A(n50178), .B(n42706), .Y(n26345) );
  XNOR2X1 U48316 ( .A(n50393), .B(n41287), .Y(n26346) );
  XNOR2X1 U48317 ( .A(n51238), .B(n42697), .Y(n26347) );
  NOR4X1 U48318 ( .A(n26315), .B(n26316), .C(n26317), .D(n26318), .Y(net215122) );
  XNOR2X1 U48319 ( .A(n50177), .B(n42711), .Y(n26315) );
  XNOR2X1 U48320 ( .A(n50392), .B(n41287), .Y(n26316) );
  XNOR2X1 U48321 ( .A(n51237), .B(n42697), .Y(n26317) );
  NOR4X1 U48322 ( .A(n26375), .B(n26376), .C(n26377), .D(n26378), .Y(n44346)
         );
  XNOR2X1 U48323 ( .A(n50175), .B(n42706), .Y(n26375) );
  XNOR2X1 U48324 ( .A(n50390), .B(n42717), .Y(n26376) );
  XNOR2X1 U48325 ( .A(n51235), .B(n42697), .Y(n26377) );
  NOR4X1 U48326 ( .A(n26165), .B(n26166), .C(n26167), .D(n26168), .Y(net215095) );
  XNOR2X1 U48327 ( .A(n50198), .B(n42705), .Y(n26165) );
  XNOR2X1 U48328 ( .A(n50413), .B(n42717), .Y(n26166) );
  XNOR2X1 U48329 ( .A(n51258), .B(n42697), .Y(n26167) );
  NOR4X1 U48330 ( .A(n26135), .B(n26136), .C(n26137), .D(n26138), .Y(n44368)
         );
  XNOR2X1 U48331 ( .A(n50197), .B(n42712), .Y(n26135) );
  XNOR2X1 U48332 ( .A(n50412), .B(n42717), .Y(n26136) );
  XNOR2X1 U48333 ( .A(n51257), .B(n42696), .Y(n26137) );
  NOR4X1 U48334 ( .A(n26105), .B(n26106), .C(n26107), .D(n26108), .Y(n44373)
         );
  XNOR2X1 U48335 ( .A(n50196), .B(n42705), .Y(n26105) );
  XNOR2X1 U48336 ( .A(n50411), .B(n42724), .Y(n26106) );
  XNOR2X1 U48337 ( .A(n51256), .B(n42690), .Y(n26107) );
  NOR4X1 U48338 ( .A(n26285), .B(n26286), .C(n26287), .D(n26288), .Y(n44353)
         );
  XNOR2X1 U48339 ( .A(n50182), .B(n42711), .Y(n26285) );
  XNOR2X1 U48340 ( .A(n50397), .B(n42720), .Y(n26286) );
  XNOR2X1 U48341 ( .A(n51242), .B(n42697), .Y(n26287) );
  NOR4X1 U48342 ( .A(n26225), .B(n26226), .C(n26227), .D(n26228), .Y(net214754) );
  XNOR2X1 U48343 ( .A(n50180), .B(n42706), .Y(n26225) );
  XNOR2X1 U48344 ( .A(n50395), .B(n42717), .Y(n26226) );
  XNOR2X1 U48345 ( .A(n51240), .B(n41385), .Y(n26227) );
  NOR4X1 U48346 ( .A(n26255), .B(n26256), .C(n26257), .D(n26258), .Y(net215104) );
  XNOR2X1 U48347 ( .A(n50181), .B(n41642), .Y(n26255) );
  XNOR2X1 U48348 ( .A(n50396), .B(n42720), .Y(n26256) );
  XNOR2X1 U48349 ( .A(n51241), .B(n42697), .Y(n26257) );
  XNOR2X1 U48350 ( .A(n50173), .B(n42706), .Y(n26526) );
  XNOR2X1 U48351 ( .A(n50388), .B(n42717), .Y(n26527) );
  NOR4X1 U48352 ( .A(n26496), .B(n26497), .C(n26498), .D(n26499), .Y(n44326)
         );
  XNOR2X1 U48353 ( .A(n50174), .B(n42706), .Y(n26496) );
  XNOR2X1 U48354 ( .A(n50389), .B(n34435), .Y(n26497) );
  XNOR2X1 U48355 ( .A(n50172), .B(n42706), .Y(n26466) );
  XNOR2X1 U48356 ( .A(n50387), .B(n34435), .Y(n26467) );
  OAI21XL U48357 ( .A0(n9988), .A1(n9989), .B0(n49518), .Y(n9986) );
  OAI211X1 U48358 ( .A0(n9990), .A1(n9991), .B0(n9992), .C0(n9993), .Y(n9989)
         );
  NOR3X1 U48359 ( .A(n9994), .B(net171528), .C(n9996), .Y(n9990) );
  NOR4X1 U48360 ( .A(net171530), .B(n9998), .C(n9999), .D(n9900), .Y(n9996) );
  NOR4X1 U48361 ( .A(n30916), .B(n30917), .C(n30918), .D(n30919), .Y(n43415)
         );
  NOR4X1 U48362 ( .A(n30525), .B(n30526), .C(n30527), .D(n30528), .Y(n43454)
         );
  XNOR2X1 U48363 ( .A(n50656), .B(net219434), .Y(n30527) );
  NOR4X1 U48364 ( .A(n30615), .B(n30616), .C(n30617), .D(n30618), .Y(n43465)
         );
  NOR4X1 U48365 ( .A(n30223), .B(n30224), .C(n30225), .D(n30226), .Y(n43489)
         );
  NOR4X1 U48366 ( .A(n30132), .B(n30133), .C(n30134), .D(n30135), .Y(net216299) );
  XNOR2X1 U48367 ( .A(n51068), .B(n41281), .Y(n30133) );
  XNOR2X1 U48368 ( .A(n50640), .B(net219442), .Y(n30134) );
  NOR4X1 U48369 ( .A(n30192), .B(n30193), .C(n30194), .D(n30195), .Y(n43497)
         );
  XNOR2X1 U48370 ( .A(n50851), .B(net219310), .Y(n30192) );
  NOR4X1 U48371 ( .A(n30072), .B(n30073), .C(n30074), .D(n30075), .Y(n43509)
         );
  XNOR2X1 U48372 ( .A(n50850), .B(n40039), .Y(n30072) );
  XNOR2X1 U48373 ( .A(n51064), .B(n41281), .Y(n30073) );
  XNOR2X1 U48374 ( .A(n50636), .B(net219442), .Y(n30074) );
  NOR4X1 U48375 ( .A(n30042), .B(n30043), .C(n30044), .D(n30045), .Y(net216272) );
  XNOR2X1 U48376 ( .A(n50849), .B(net258262), .Y(n30042) );
  XNOR2X1 U48377 ( .A(n51063), .B(n41282), .Y(n30043) );
  XNOR2X1 U48378 ( .A(n50635), .B(net219442), .Y(n30044) );
  NOR4X1 U48379 ( .A(n30012), .B(n30013), .C(n30014), .D(n30015), .Y(net216263) );
  XNOR2X1 U48380 ( .A(n50848), .B(net219330), .Y(n30012) );
  XNOR2X1 U48381 ( .A(n51062), .B(n41283), .Y(n30013) );
  XNOR2X1 U48382 ( .A(n50634), .B(net219442), .Y(n30014) );
  NOR4X1 U48383 ( .A(n30102), .B(n30103), .C(n30104), .D(n30105), .Y(net216290) );
  XNOR2X1 U48384 ( .A(n50853), .B(net219310), .Y(n30102) );
  XNOR2X1 U48385 ( .A(n51067), .B(n41282), .Y(n30103) );
  XNOR2X1 U48386 ( .A(n50639), .B(net219442), .Y(n30104) );
  NOR4X1 U48387 ( .A(n29802), .B(n29803), .C(n29804), .D(n29805), .Y(n43518)
         );
  XNOR2X1 U48388 ( .A(n51057), .B(n41282), .Y(n29803) );
  XNOR2X1 U48389 ( .A(n50629), .B(net219442), .Y(n29804) );
  NOR4X1 U48390 ( .A(n30162), .B(n30163), .C(n30164), .D(n30165), .Y(net216308) );
  XNOR2X1 U48391 ( .A(n50852), .B(net219308), .Y(n30162) );
  XNOR2X1 U48392 ( .A(n51066), .B(n41281), .Y(n30163) );
  XNOR2X1 U48393 ( .A(n50638), .B(net219442), .Y(n30164) );
  NOR4X1 U48394 ( .A(n30826), .B(n30827), .C(n30828), .D(n30829), .Y(net216488) );
  NOR4X1 U48395 ( .A(n30675), .B(n30676), .C(n30677), .D(n30678), .Y(net216407) );
  NOR4X1 U48396 ( .A(n30495), .B(n30496), .C(n30497), .D(n30498), .Y(net216434) );
  NOR4X1 U48397 ( .A(n30465), .B(n30466), .C(n30467), .D(n30468), .Y(net216425) );
  NOR4X1 U48398 ( .A(n29501), .B(n29502), .C(n29503), .D(n29504), .Y(n43537)
         );
  NOR4X1 U48399 ( .A(n29952), .B(n29953), .C(n29954), .D(n29955), .Y(n44579)
         );
  XNOR2X1 U48400 ( .A(n50842), .B(net219310), .Y(n29952) );
  XNOR2X1 U48401 ( .A(n51056), .B(n41282), .Y(n29953) );
  XNOR2X1 U48402 ( .A(n50628), .B(net219442), .Y(n29954) );
  NOR4X1 U48403 ( .A(n29621), .B(n29622), .C(n29623), .D(n29624), .Y(n43542)
         );
  XNOR2X1 U48404 ( .A(n50839), .B(net219314), .Y(n29922) );
  XNOR2X1 U48405 ( .A(n51053), .B(n41281), .Y(n29923) );
  XNOR2X1 U48406 ( .A(n50625), .B(net219442), .Y(n29924) );
  NOR4X1 U48407 ( .A(n30433), .B(n30434), .C(n30435), .D(n30436), .Y(net216344) );
  NOR4X1 U48408 ( .A(n30343), .B(n30344), .C(n30345), .D(n30346), .Y(net214786) );
  XNOR2X1 U48409 ( .A(n50840), .B(n36870), .Y(n29862) );
  XNOR2X1 U48410 ( .A(n51054), .B(n41283), .Y(n29863) );
  XNOR2X1 U48411 ( .A(n50626), .B(net219442), .Y(n29864) );
  NOR4X1 U48412 ( .A(n30373), .B(n30374), .C(n30375), .D(n30376), .Y(net216326) );
  XNOR2X1 U48413 ( .A(n51058), .B(n41283), .Y(n29833) );
  XNOR2X1 U48414 ( .A(n50630), .B(net219442), .Y(n29834) );
  XNOR2X1 U48415 ( .A(n50841), .B(net219310), .Y(n29892) );
  XNOR2X1 U48416 ( .A(n51055), .B(n41281), .Y(n29893) );
  XNOR2X1 U48417 ( .A(n50627), .B(net219442), .Y(n29894) );
  NOR4X1 U48418 ( .A(n29561), .B(n29562), .C(n29563), .D(n29564), .Y(net216191) );
  NOR4X1 U48419 ( .A(n30555), .B(n30556), .C(n30557), .D(n30558), .Y(net216443) );
  XNOR2X1 U48420 ( .A(n50864), .B(net219336), .Y(n30555) );
  XNOR2X1 U48421 ( .A(n51078), .B(n41283), .Y(n30556) );
  NOR4X1 U48422 ( .A(n30585), .B(n30586), .C(n30587), .D(n30588), .Y(n43434)
         );
  NOR4X1 U48423 ( .A(n30313), .B(n30314), .C(n30315), .D(n30316), .Y(n43474)
         );
  NOR4X1 U48424 ( .A(n30283), .B(n30284), .C(n30285), .D(n30286), .Y(n43483)
         );
  XNOR2X1 U48425 ( .A(n50861), .B(net219310), .Y(n30283) );
  XNOR2X1 U48426 ( .A(n51075), .B(n41282), .Y(n30284) );
  NOR4X1 U48427 ( .A(n26405), .B(n26406), .C(n26407), .D(n26408), .Y(net215147) );
  XNOR2X1 U48428 ( .A(n50176), .B(n42706), .Y(n26405) );
  XNOR2X1 U48429 ( .A(n50391), .B(n42720), .Y(n26406) );
  XNOR2X1 U48430 ( .A(n51236), .B(n42697), .Y(n26407) );
  NOR4X1 U48431 ( .A(n30645), .B(n30646), .C(n30647), .D(n30648), .Y(net216396) );
  XNOR2X1 U48432 ( .A(n50847), .B(n40039), .Y(n29982) );
  XNOR2X1 U48433 ( .A(n51061), .B(n41282), .Y(n29983) );
  XNOR2X1 U48434 ( .A(n50633), .B(net219442), .Y(n29984) );
  NAND4BX1 U48435 ( .AN(n10641), .B(net271515), .C(n39342), .D(n21862), .Y(
        n9994) );
  AND3X2 U48436 ( .A(n10761), .B(n10760), .C(n10759), .Y(n21862) );
  NAND4X1 U48437 ( .A(n10763), .B(net210556), .C(net210555), .D(n23606), .Y(
        n10198) );
  AND2X2 U48438 ( .A(n10762), .B(n37348), .Y(n23606) );
  NAND4BBXL U48439 ( .AN(net210531), .BN(n48468), .C(net212664), .D(n10257),
        .Y(n47805) );
  OAI21XL U48440 ( .A0(n42316), .A1(n9750), .B0(n9751), .Y(nxt_data_num[0]) );
  OAI31XL U48441 ( .A0(n9748), .A1(n9743), .A2(n41790), .B0(n42316), .Y(n9751)
         );
  NOR2X1 U48442 ( .A(n41789), .B(n9744), .Y(n9750) );
  AND2X2 U48443 ( .A(n10848), .B(n10852), .Y(n24010) );
  CLKINVX1 U48444 ( .A(n10484), .Y(net171152) );
  NAND4X1 U48445 ( .A(n10847), .B(n10845), .C(n10846), .D(n24091), .Y(n47807)
         );
  NAND2X1 U48446 ( .A(n12855), .B(n12858), .Y(n11521) );
  NAND4BBXL U48447 ( .AN(net210522), .BN(net210525), .C(net210524), .D(n47663),
        .Y(n47823) );
  NAND4X1 U48448 ( .A(n10638), .B(n10635), .C(n39341), .D(n20877), .Y(n9991)
         );
  AND2X2 U48449 ( .A(n10639), .B(n10632), .Y(n20877) );
  OAI21XL U48450 ( .A0(n47811), .A1(n47835), .B0(n47810), .Y(n47813) );
  OAI21XL U48451 ( .A0(n47825), .A1(n47824), .B0(n41744), .Y(n47827) );
  AOI211X1 U48452 ( .A0(n10000), .A1(n10001), .B0(n10002), .C0(n39923), .Y(
        n9998) );
  NAND2X1 U48453 ( .A(n10004), .B(n10005), .Y(n10002) );
  OAI21XL U48454 ( .A0(n10006), .A1(n9880), .B0(n50108), .Y(n10001) );
  NOR3X1 U48455 ( .A(n43038), .B(n50134), .C(n9726), .Y(n9724) );
  NAND2X1 U48456 ( .A(n23687), .B(n23688), .Y(n9979) );
  OAI21XL U48457 ( .A0(n10255), .A1(n9978), .B0(n50096), .Y(n10252) );
  NOR2X1 U48458 ( .A(n47806), .B(n47805), .Y(n10255) );
  NOR2X1 U48459 ( .A(n47804), .B(n47803), .Y(n47806) );
  OAI21XL U48460 ( .A0(n10152), .A1(n10153), .B0(n49498), .Y(n10149) );
  CLKINVX1 U48461 ( .A(n9840), .Y(n49498) );
  OAI211X1 U48462 ( .A0(n10155), .A1(n10156), .B0(n10157), .C0(n10158), .Y(
        n10153) );
  OAI31XL U48463 ( .A0(n50100), .A1(net171214), .A2(n10161), .B0(n10162), .Y(
        n10156) );
  AND4X1 U48464 ( .A(net151587), .B(n10959), .C(n24174), .D(n24175), .Y(n9969)
         );
  NOR4X1 U48465 ( .A(net151586), .B(net171412), .C(net151584), .D(net171414),
        .Y(n24175) );
  NOR2X1 U48466 ( .A(n39537), .B(n10215), .Y(n24174) );
  AND4X1 U48467 ( .A(n10983), .B(n_cell_303546_net275959), .C(n24376), .D(
        n24377), .Y(n10216) );
  AND2X2 U48468 ( .A(n_cell_303546_net275923), .B(net271956), .Y(n24376) );
  NOR4X1 U48469 ( .A(net171398), .B(net171401), .C(net151536), .D(net151541),
        .Y(n24377) );
  NAND3X1 U48470 ( .A(n20424), .B(n10614), .C(n37342), .Y(n47822) );
  AND2X2 U48471 ( .A(n37016), .B(n10619), .Y(n20424) );
  NAND4BX1 U48472 ( .AN(n48715), .B(n48714), .C(n48713), .D(n48712), .Y(n34529) );
  NAND2X1 U48473 ( .A(n51225), .B(net265207), .Y(n48712) );
  NAND2X1 U48474 ( .A(n40273), .B(n49513), .Y(n49174) );
  NAND4X1 U48475 ( .A(n13096), .B(n48870), .C(n48869), .D(n48868), .Y(n34538)
         );
  NAND4X1 U48476 ( .A(n13099), .B(n49022), .C(n49021), .D(n49020), .Y(n34539)
         );
  NAND4X1 U48477 ( .A(n13105), .B(n49177), .C(n49176), .D(n49175), .Y(n34541)
         );
  NAND4X1 U48478 ( .A(n13084), .B(n49332), .C(n49331), .D(n49330), .Y(n34534)
         );
  NAND4X1 U48479 ( .A(n13079), .B(n49180), .C(n49179), .D(n49178), .Y(n34533)
         );
  NAND4X1 U48480 ( .A(n13052), .B(n49335), .C(n49334), .D(n49333), .Y(n34526)
         );
  NAND4X1 U48481 ( .A(n13056), .B(n49490), .C(n49489), .D(n49488), .Y(n34527)
         );
  NAND4X1 U48482 ( .A(n13093), .B(n48711), .C(n48710), .D(n48709), .Y(n34537)
         );
  NAND4X1 U48483 ( .A(n13087), .B(n49487), .C(n49486), .D(n49485), .Y(n34535)
         );
  OAI211X1 U48484 ( .A0(n10235), .A1(n10236), .B0(n10237), .C0(net151652), .Y(
        n10234) );
  CLKINVX1 U48485 ( .A(n10239), .Y(net151652) );
  OAI31XL U48486 ( .A0(n10240), .A1(n10241), .A2(n10242), .B0(n10243), .Y(
        n10236) );
  AND4X1 U48487 ( .A(n10000), .B(n10004), .C(n10005), .D(n10646), .Y(n9898) );
  NAND2X1 U48488 ( .A(n51438), .B(n40243), .Y(n48708) );
  NAND2X1 U48489 ( .A(n51011), .B(n40256), .Y(n48870) );
  NAND2X1 U48490 ( .A(n50797), .B(n40225), .Y(n49022) );
  NAND2X1 U48491 ( .A(n50583), .B(n40222), .Y(n49177) );
  CLKINVX1 U48492 ( .A(n12639), .Y(net209733) );
  NAND4X1 U48493 ( .A(n10626), .B(n10625), .C(n10624), .D(n20015), .Y(n9877)
         );
  NOR2X1 U48494 ( .A(net151785), .B(n10621), .Y(n20015) );
  CLKINVX1 U48495 ( .A(n10622), .Y(net151785) );
  NAND2X1 U48496 ( .A(n40195), .B(n49515), .Y(n49019) );
  NAND2X1 U48497 ( .A(net217942), .B(n49512), .Y(n49329) );
  NAND2X1 U48498 ( .A(n40220), .B(n49510), .Y(n49484) );
  NAND2X1 U48499 ( .A(n40276), .B(n49164), .Y(n49163) );
  NAND2X1 U48500 ( .A(n40271), .B(n48598), .Y(n48597) );
  NAND2X1 U48501 ( .A(n40271), .B(n48602), .Y(n48601) );
  NAND2X1 U48502 ( .A(n40271), .B(n48606), .Y(n48605) );
  NAND2X1 U48503 ( .A(n40271), .B(n48610), .Y(n48609) );
  NAND2X1 U48504 ( .A(n40271), .B(n48614), .Y(n48613) );
  NAND2X1 U48505 ( .A(n40271), .B(n48618), .Y(n48617) );
  NAND2X1 U48506 ( .A(n40271), .B(n48622), .Y(n48621) );
  NAND2X1 U48507 ( .A(n40271), .B(n48626), .Y(n48625) );
  NAND2X1 U48508 ( .A(n40271), .B(n48630), .Y(n48629) );
  NAND2X1 U48509 ( .A(n40271), .B(n48634), .Y(n48633) );
  NAND2X1 U48510 ( .A(n40271), .B(n48638), .Y(n48637) );
  NAND2X1 U48511 ( .A(n40271), .B(n48642), .Y(n48641) );
  NAND2X1 U48512 ( .A(n40270), .B(n48646), .Y(n48645) );
  NAND2X1 U48513 ( .A(n40270), .B(n48650), .Y(n48649) );
  NAND2X1 U48514 ( .A(n40270), .B(n48654), .Y(n48653) );
  NAND2X1 U48515 ( .A(n40270), .B(n48658), .Y(n48657) );
  NAND2X1 U48516 ( .A(n40270), .B(n48662), .Y(n48661) );
  NAND2X1 U48517 ( .A(n40270), .B(n48666), .Y(n48665) );
  NAND2X1 U48518 ( .A(n40270), .B(n48670), .Y(n48669) );
  NAND2X1 U48519 ( .A(n40270), .B(n48674), .Y(n48673) );
  NAND2X1 U48520 ( .A(n40270), .B(n48682), .Y(n48681) );
  NAND2X1 U48521 ( .A(n40270), .B(n48686), .Y(n48685) );
  NAND2X1 U48522 ( .A(n40270), .B(n48690), .Y(n48689) );
  NAND2X1 U48523 ( .A(n40269), .B(n48694), .Y(n48693) );
  NAND2X1 U48524 ( .A(n40269), .B(n48698), .Y(n48697) );
  NAND2X1 U48525 ( .A(n40269), .B(n48705), .Y(n48704) );
  NAND2X1 U48526 ( .A(n40269), .B(n48726), .Y(n48725) );
  NAND2X1 U48527 ( .A(n40269), .B(n48730), .Y(n48729) );
  NAND2X1 U48528 ( .A(n40269), .B(n48746), .Y(n48745) );
  NAND2X1 U48529 ( .A(n40274), .B(n48790), .Y(n48789) );
  NAND2X1 U48530 ( .A(n40226), .B(n48794), .Y(n48793) );
  NAND2X1 U48531 ( .A(n40268), .B(n48798), .Y(n48797) );
  NAND2X1 U48532 ( .A(n40235), .B(n48802), .Y(n48801) );
  NAND2X1 U48533 ( .A(n40228), .B(n48806), .Y(n48805) );
  NAND2X1 U48534 ( .A(n40214), .B(n48810), .Y(n48809) );
  NAND2X1 U48535 ( .A(n40232), .B(n48814), .Y(n48813) );
  NAND2X1 U48536 ( .A(n40274), .B(n48818), .Y(n48817) );
  NAND2X1 U48537 ( .A(n40248), .B(n48822), .Y(n48821) );
  NAND2X1 U48538 ( .A(n40243), .B(n48826), .Y(n48825) );
  NAND2X1 U48539 ( .A(n40268), .B(n48830), .Y(n48829) );
  NAND2X1 U48540 ( .A(n40274), .B(n48834), .Y(n48833) );
  NAND2X1 U48541 ( .A(n40267), .B(n48842), .Y(n48841) );
  NAND2X1 U48542 ( .A(n40277), .B(n48846), .Y(n48845) );
  NAND2X1 U48543 ( .A(net217940), .B(n48850), .Y(n48849) );
  NAND2X1 U48544 ( .A(n40268), .B(n48854), .Y(n48853) );
  NAND2X1 U48545 ( .A(n40274), .B(n48864), .Y(n48863) );
  NAND2X1 U48546 ( .A(n40267), .B(n48884), .Y(n48883) );
  NAND2X1 U48547 ( .A(n40267), .B(n41367), .Y(n48887) );
  NAND2X1 U48548 ( .A(n40267), .B(n48902), .Y(n48901) );
  NAND2X1 U48549 ( .A(n40267), .B(n48906), .Y(n48905) );
  NAND2X1 U48550 ( .A(n40267), .B(n48910), .Y(n48909) );
  NAND2X1 U48551 ( .A(n40227), .B(n48914), .Y(n48913) );
  NAND2X1 U48552 ( .A(n40235), .B(n48918), .Y(n48917) );
  NAND2X1 U48553 ( .A(n40230), .B(n48922), .Y(n48921) );
  NAND2X1 U48554 ( .A(n40232), .B(n48926), .Y(n48925) );
  NAND2X1 U48555 ( .A(n40187), .B(n48930), .Y(n48929) );
  NAND2X1 U48556 ( .A(n40228), .B(n48934), .Y(n48933) );
  NAND2X1 U48557 ( .A(n40188), .B(n48938), .Y(n48937) );
  NAND2X1 U48558 ( .A(n40231), .B(n48942), .Y(n48941) );
  NAND2X1 U48559 ( .A(n40221), .B(n48946), .Y(n48945) );
  NAND2X1 U48560 ( .A(n40226), .B(n48950), .Y(n48949) );
  NAND2X1 U48561 ( .A(n40247), .B(n48954), .Y(n48953) );
  NAND2X1 U48562 ( .A(n40242), .B(n48958), .Y(n48957) );
  NAND2X1 U48563 ( .A(n40268), .B(n48962), .Y(n48961) );
  NAND2X1 U48564 ( .A(n40268), .B(n48966), .Y(n48965) );
  NAND2X1 U48565 ( .A(n40268), .B(n48970), .Y(n48969) );
  NAND2X1 U48566 ( .A(n40268), .B(n48974), .Y(n48973) );
  NAND2X1 U48567 ( .A(n40268), .B(n48978), .Y(n48977) );
  NAND2X1 U48568 ( .A(n40268), .B(n48982), .Y(n48981) );
  NAND2X1 U48569 ( .A(n40268), .B(n48986), .Y(n48985) );
  NAND2X1 U48570 ( .A(n40268), .B(n48990), .Y(n48989) );
  NAND2X1 U48571 ( .A(n40268), .B(n48998), .Y(n48997) );
  NAND2X1 U48572 ( .A(n40268), .B(n49002), .Y(n49001) );
  NAND2X1 U48573 ( .A(n40268), .B(n49006), .Y(n49005) );
  NAND2X1 U48574 ( .A(net217930), .B(n41234), .Y(n49035) );
  NAND2X1 U48575 ( .A(n40191), .B(n49039), .Y(n49038) );
  NAND2X1 U48576 ( .A(net217936), .B(n49192), .Y(n49191) );
  NAND2X1 U48577 ( .A(n40273), .B(n49196), .Y(n49195) );
  NAND2X1 U48578 ( .A(n40275), .B(n49216), .Y(n49215) );
  NAND2X1 U48579 ( .A(n40275), .B(n49220), .Y(n49219) );
  NAND2X1 U48580 ( .A(n40275), .B(n49224), .Y(n49223) );
  NAND2X1 U48581 ( .A(n40275), .B(n49228), .Y(n49227) );
  NAND2X1 U48582 ( .A(n40275), .B(n49232), .Y(n49231) );
  NAND2X1 U48583 ( .A(n40275), .B(n49236), .Y(n49235) );
  NAND2X1 U48584 ( .A(n40275), .B(n49240), .Y(n49239) );
  NAND2X1 U48585 ( .A(n40275), .B(n49244), .Y(n49243) );
  NAND2X1 U48586 ( .A(n40274), .B(n49248), .Y(n49247) );
  NAND2X1 U48587 ( .A(n40274), .B(n49252), .Y(n49251) );
  NAND2X1 U48588 ( .A(n40274), .B(n49256), .Y(n49255) );
  NAND2X1 U48589 ( .A(n40274), .B(n49260), .Y(n49259) );
  NAND2X1 U48590 ( .A(n40274), .B(n49264), .Y(n49263) );
  NAND2X1 U48591 ( .A(n40274), .B(n49268), .Y(n49267) );
  NAND2X1 U48592 ( .A(n40274), .B(n49272), .Y(n49271) );
  NAND2X1 U48593 ( .A(n40274), .B(n49276), .Y(n49275) );
  NAND2X1 U48594 ( .A(n40274), .B(n49280), .Y(n49279) );
  NAND2X1 U48595 ( .A(n40274), .B(n49284), .Y(n49283) );
  NAND2X1 U48596 ( .A(n40274), .B(n49288), .Y(n49287) );
  NAND2X1 U48597 ( .A(n40274), .B(n41227), .Y(n49291) );
  NAND2X1 U48598 ( .A(n40254), .B(n49295), .Y(n49294) );
  NAND2X1 U48599 ( .A(n40188), .B(n49299), .Y(n49298) );
  NAND2X1 U48600 ( .A(n40225), .B(n49307), .Y(n49306) );
  NAND2X1 U48601 ( .A(n40187), .B(n49311), .Y(n49310) );
  NAND2X1 U48602 ( .A(n40222), .B(n49315), .Y(n49314) );
  NAND2X1 U48603 ( .A(n40229), .B(n49319), .Y(n49318) );
  NAND2X1 U48604 ( .A(net217944), .B(n49347), .Y(n49346) );
  NAND2X1 U48605 ( .A(n40275), .B(n49351), .Y(n49350) );
  NAND2X1 U48606 ( .A(n40275), .B(n49367), .Y(n49366) );
  NAND2X1 U48607 ( .A(net217944), .B(n49371), .Y(n49370) );
  NAND2X1 U48608 ( .A(net217944), .B(n49375), .Y(n49374) );
  NAND2X1 U48609 ( .A(net217944), .B(n49379), .Y(n49378) );
  NAND2X1 U48610 ( .A(n40275), .B(n49383), .Y(n49382) );
  NAND2X1 U48611 ( .A(net217944), .B(n49387), .Y(n49386) );
  NAND2X1 U48612 ( .A(n40275), .B(n49391), .Y(n49390) );
  NAND2X1 U48613 ( .A(n40273), .B(n49395), .Y(n49394) );
  NAND2X1 U48614 ( .A(n40273), .B(n49399), .Y(n49398) );
  NAND2X1 U48615 ( .A(n40273), .B(n49403), .Y(n49402) );
  NAND2X1 U48616 ( .A(n40273), .B(n49407), .Y(n49406) );
  NAND2X1 U48617 ( .A(n40273), .B(n49411), .Y(n49410) );
  NAND2X1 U48618 ( .A(n40273), .B(n49415), .Y(n49414) );
  NAND2X1 U48619 ( .A(n40273), .B(n49419), .Y(n49418) );
  NAND2X1 U48620 ( .A(n40273), .B(n49423), .Y(n49422) );
  NAND2X1 U48621 ( .A(n40273), .B(n41221), .Y(n49426) );
  NAND2X1 U48622 ( .A(n40273), .B(n49430), .Y(n49429) );
  NAND2X1 U48623 ( .A(n40273), .B(n49434), .Y(n49433) );
  NAND2X1 U48624 ( .A(n40273), .B(n49438), .Y(n49437) );
  NAND2X1 U48625 ( .A(n40269), .B(n48742), .Y(n48741) );
  NAND2X1 U48626 ( .A(n40267), .B(n41655), .Y(n48898) );
  NAND2X1 U48627 ( .A(net217944), .B(n49363), .Y(n49362) );
  NAND2X1 U48628 ( .A(n40270), .B(n48678), .Y(n48677) );
  NAND2X1 U48629 ( .A(n40267), .B(n48838), .Y(n48837) );
  NAND2X1 U48630 ( .A(n40268), .B(n48994), .Y(n48993) );
  NAND2X1 U48631 ( .A(n40275), .B(n49212), .Y(n49211) );
  NAND2X1 U48632 ( .A(n40233), .B(n49303), .Y(n49302) );
  NAND2X1 U48633 ( .A(n40269), .B(n48734), .Y(n48733) );
  NAND2X1 U48634 ( .A(n40269), .B(n48738), .Y(n48737) );
  NAND2X1 U48635 ( .A(n40267), .B(n48891), .Y(n48890) );
  NAND2X1 U48636 ( .A(n40267), .B(n48895), .Y(n48894) );
  NAND2X1 U48637 ( .A(n40226), .B(n49043), .Y(n49042) );
  NAND2X1 U48638 ( .A(n40277), .B(n49066), .Y(n49065) );
  NAND2X1 U48639 ( .A(n40277), .B(n49082), .Y(n49081) );
  NAND2X1 U48640 ( .A(n40276), .B(n49152), .Y(n49151) );
  NAND2X1 U48641 ( .A(n40275), .B(n49208), .Y(n49207) );
  NAND2X1 U48642 ( .A(n40275), .B(n49359), .Y(n49358) );
  NAND2X1 U48643 ( .A(n40235), .B(n41349), .Y(n49054) );
  NAND2X1 U48644 ( .A(n40277), .B(n49078), .Y(n49077) );
  NAND2X1 U48645 ( .A(n40228), .B(n49047), .Y(n49046) );
  NAND2X1 U48646 ( .A(n40258), .B(n49051), .Y(n49050) );
  NAND2X1 U48647 ( .A(n40255), .B(n49058), .Y(n49057) );
  NAND2X1 U48648 ( .A(n40277), .B(n49062), .Y(n49061) );
  NAND2X1 U48649 ( .A(n40277), .B(n49070), .Y(n49069) );
  NAND2X1 U48650 ( .A(n40277), .B(n49074), .Y(n49073) );
  NAND2X1 U48651 ( .A(n40277), .B(n49086), .Y(n49085) );
  NAND2X1 U48652 ( .A(n40277), .B(n49090), .Y(n49089) );
  NAND2X1 U48653 ( .A(n40277), .B(n49094), .Y(n49093) );
  NAND2X1 U48654 ( .A(n40277), .B(n49098), .Y(n49097) );
  NAND2X1 U48655 ( .A(n40277), .B(n49102), .Y(n49101) );
  NAND2X1 U48656 ( .A(n40277), .B(n49106), .Y(n49105) );
  NAND2X1 U48657 ( .A(n40276), .B(n49110), .Y(n49109) );
  NAND2X1 U48658 ( .A(n40276), .B(n49114), .Y(n49113) );
  NAND2X1 U48659 ( .A(n40276), .B(n49118), .Y(n49117) );
  NAND2X1 U48660 ( .A(n40276), .B(n49122), .Y(n49121) );
  NAND2X1 U48661 ( .A(n40276), .B(n49126), .Y(n49125) );
  NAND2X1 U48662 ( .A(n40276), .B(n49130), .Y(n49129) );
  NAND2X1 U48663 ( .A(n40276), .B(n41231), .Y(n49133) );
  NAND2X1 U48664 ( .A(n40276), .B(n49137), .Y(n49136) );
  NAND2X1 U48665 ( .A(n40276), .B(n49141), .Y(n49140) );
  NAND2X1 U48666 ( .A(n40276), .B(n41259), .Y(n49144) );
  NAND2X1 U48667 ( .A(n40276), .B(n49148), .Y(n49147) );
  NAND2X1 U48668 ( .A(n40273), .B(n49156), .Y(n49155) );
  NAND2X1 U48669 ( .A(n40273), .B(n49160), .Y(n49159) );
  NAND2X1 U48670 ( .A(net217936), .B(n49171), .Y(n49170) );
  NAND2X1 U48671 ( .A(n40276), .B(n49200), .Y(n49199) );
  NAND2X1 U48672 ( .A(n40275), .B(n49204), .Y(n49203) );
  NAND2X1 U48673 ( .A(net217944), .B(n49355), .Y(n49354) );
  NAND2X1 U48674 ( .A(n40269), .B(n41643), .Y(n48719) );
  NAND2X1 U48675 ( .A(n40267), .B(n41345), .Y(n48877) );
  NAND2X1 U48676 ( .A(n40242), .B(n49029), .Y(n49028) );
  NAND2X1 U48677 ( .A(net217936), .B(n49185), .Y(n49184) );
  NAND2X1 U48678 ( .A(n40221), .B(n49340), .Y(n49339) );
  NAND2X1 U48679 ( .A(n51225), .B(n40214), .Y(n48711) );
  NAND2X1 U48680 ( .A(n50165), .B(n40248), .Y(n49487) );
  AOI31X1 U48681 ( .A0(n10199), .A1(n10200), .A2(n37346), .B0(n9870), .Y(n9982) );
  NAND3X1 U48682 ( .A(n37123), .B(n10203), .C(n10204), .Y(n10200) );
  NAND4X1 U48683 ( .A(n10205), .B(n10206), .C(net151587), .D(n10208), .Y(
        n10203) );
  OAI222XL U48684 ( .A0(n49553), .A1(n19493), .B0(n42544), .B1(n43040), .C0(
        n36796), .C1(n43044), .Y(n19498) );
  OAI222XL U48685 ( .A0(n49554), .A1(n19493), .B0(n42526), .B1(n43040), .C0(
        n36754), .C1(n43044), .Y(n19494) );
  OAI222XL U48686 ( .A0(n49555), .A1(n19493), .B0(n42508), .B1(n43040), .C0(
        n42473), .C1(n43044), .Y(n19488) );
  OAI222XL U48687 ( .A0(n49548), .A1(n19493), .B0(n42584), .B1(n43040), .C0(
        n36768), .C1(n43043), .Y(n19518) );
  OAI221XL U48688 ( .A0(n9708), .A1(n50087), .B0(n50147), .B1(n49522), .C0(
        n9712), .Y(n9706) );
  CLKINVX1 U48689 ( .A(n9689), .Y(n49522) );
  AOI211X1 U48690 ( .A0(net171349), .A1(n9714), .B0(n50147), .C0(n9715), .Y(
        n9708) );
  OAI21XL U48691 ( .A0(n42316), .A1(n9716), .B0(n50135), .Y(n9714) );
  NOR4X1 U48692 ( .A(n10532), .B(n39815), .C(net171205), .D(net171210), .Y(
        n10196) );
  NAND4X1 U48693 ( .A(net260449), .B(net260394), .C(n10438), .D(n26409), .Y(
        n9922) );
  NOR4X1 U48694 ( .A(net171259), .B(net171262), .C(net151773), .D(net151775),
        .Y(n26409) );
  NAND4X1 U48695 ( .A(n11883), .B(n11884), .C(n11885), .D(n11886), .Y(n10130)
         );
  NOR2X1 U48696 ( .A(net171145), .B(n10492), .Y(n30683) );
  NAND4X1 U48697 ( .A(n10520), .B(n10519), .C(n11994), .D(n31645), .Y(n9840)
         );
  NOR3X1 U48698 ( .A(n10522), .B(net171117), .C(n10518), .Y(n31645) );
  XNOR2X1 U48699 ( .A(n50826), .B(n36797), .Y(n20923) );
  XNOR2X1 U48700 ( .A(n50823), .B(n36793), .Y(n20892) );
  XNOR2X1 U48701 ( .A(n50820), .B(n36795), .Y(n20850) );
  XNOR2X1 U48702 ( .A(n50819), .B(n36791), .Y(n20839) );
  XNOR2X1 U48703 ( .A(n50824), .B(n36792), .Y(n20882) );
  XNOR2X1 U48704 ( .A(n50818), .B(n36789), .Y(n20870) );
  XNOR2X1 U48705 ( .A(n50817), .B(n36790), .Y(n20860) );
  XNOR2X1 U48706 ( .A(n50815), .B(n36795), .Y(n20807) );
  XNOR2X1 U48707 ( .A(n50814), .B(n36789), .Y(n20828) );
  XNOR2X1 U48708 ( .A(n50813), .B(n36793), .Y(n20818) );
  XNOR2X1 U48709 ( .A(n50859), .B(n41290), .Y(n24452) );
  XNOR2X1 U48710 ( .A(n50859), .B(n36796), .Y(n22058) );
  XNOR2X1 U48711 ( .A(n50858), .B(n41294), .Y(n24442) );
  XNOR2X1 U48712 ( .A(n50860), .B(n36798), .Y(n22068) );
  XNOR2X1 U48713 ( .A(n50858), .B(n36792), .Y(n22048) );
  XNOR2X1 U48714 ( .A(n50855), .B(n41293), .Y(n24402) );
  XNOR2X1 U48715 ( .A(n50857), .B(n36789), .Y(n22038) );
  XNOR2X1 U48716 ( .A(n50854), .B(n41292), .Y(n24392) );
  XNOR2X1 U48717 ( .A(n50851), .B(n41296), .Y(n24472) );
  XNOR2X1 U48718 ( .A(n50850), .B(n41293), .Y(n24462) );
  XNOR2X1 U48719 ( .A(n50850), .B(n36798), .Y(n21988) );
  XNOR2X1 U48720 ( .A(n50849), .B(n36795), .Y(n21978) );
  XNOR2X1 U48721 ( .A(n50847), .B(n36790), .Y(n21948) );
  XNOR2X1 U48722 ( .A(n50844), .B(n41294), .Y(n24270) );
  XNOR2X1 U48723 ( .A(n50856), .B(n41297), .Y(n24422) );
  XNOR2X1 U48724 ( .A(n50846), .B(n36797), .Y(n21968) );
  XNOR2X1 U48725 ( .A(n50843), .B(n41292), .Y(n24260) );
  XNOR2X1 U48726 ( .A(n50857), .B(n41292), .Y(n24432) );
  XNOR2X1 U48727 ( .A(n50845), .B(n36796), .Y(n21958) );
  XNOR2X1 U48728 ( .A(n50842), .B(n41296), .Y(n24250) );
  XNOR2X1 U48729 ( .A(n50840), .B(n41291), .Y(n24290) );
  XNOR2X1 U48730 ( .A(n50852), .B(n41295), .Y(n24482) );
  XNOR2X1 U48731 ( .A(n50846), .B(n41296), .Y(n24350) );
  XNOR2X1 U48732 ( .A(n50845), .B(n41291), .Y(n24340) );
  XNOR2X1 U48733 ( .A(n50838), .B(n41291), .Y(n24240) );
  XNOR2X1 U48734 ( .A(n50839), .B(n36797), .Y(n21856) );
  XNOR2X1 U48735 ( .A(n50848), .B(n41293), .Y(n24370) );
  XNOR2X1 U48736 ( .A(n50847), .B(n41297), .Y(n24360) );
  XNOR2X1 U48737 ( .A(n50856), .B(n36796), .Y(n22018) );
  XNOR2X1 U48738 ( .A(n50855), .B(n36799), .Y(n22028) );
  XNOR2X1 U48739 ( .A(n50851), .B(n36792), .Y(n21998) );
  XNOR2X1 U48740 ( .A(n50852), .B(n36798), .Y(n22008) );
  XNOR2X1 U48741 ( .A(n50841), .B(n41296), .Y(n24280) );
  XNOR2X1 U48742 ( .A(n50835), .B(n36793), .Y(n21907) );
  XNOR2X1 U48743 ( .A(n50832), .B(n41292), .Y(n24330) );
  XNOR2X1 U48744 ( .A(n50836), .B(n36798), .Y(n21826) );
  XNOR2X1 U48745 ( .A(n50834), .B(n36799), .Y(n21928) );
  XNOR2X1 U48746 ( .A(n50831), .B(n41294), .Y(n24320) );
  XNOR2X1 U48747 ( .A(n50833), .B(n36795), .Y(n21918) );
  XNOR2X1 U48748 ( .A(n50831), .B(n36795), .Y(n21887) );
  XNOR2X1 U48749 ( .A(n50830), .B(n41291), .Y(n24300) );
  XNOR2X1 U48750 ( .A(n50829), .B(n41296), .Y(n24310) );
  XNOR2X1 U48751 ( .A(n50840), .B(n36789), .Y(n21816) );
  XNOR2X1 U48752 ( .A(n50837), .B(n36793), .Y(n21836) );
  XNOR2X1 U48753 ( .A(n50838), .B(n36798), .Y(n21846) );
  XNOR2X1 U48754 ( .A(n50828), .B(n41291), .Y(n24604) );
  XNOR2X1 U48755 ( .A(n50827), .B(n41293), .Y(n24614) );
  XNOR2X1 U48756 ( .A(n50832), .B(n36791), .Y(n21897) );
  XNOR2X1 U48757 ( .A(n50830), .B(n36795), .Y(n21867) );
  XNOR2X1 U48758 ( .A(n50825), .B(n41295), .Y(n24584) );
  XNOR2X1 U48759 ( .A(n50826), .B(n41294), .Y(n24594) );
  XNOR2X1 U48760 ( .A(n50829), .B(n36796), .Y(n21877) );
  XNOR2X1 U48761 ( .A(n50824), .B(n41290), .Y(n24564) );
  XNOR2X1 U48762 ( .A(n50821), .B(n41297), .Y(n24574) );
  XNOR2X1 U48763 ( .A(n50817), .B(n41296), .Y(n24624) );
  XNOR2X1 U48764 ( .A(n50823), .B(n41296), .Y(n24542) );
  XNOR2X1 U48765 ( .A(n50822), .B(n41293), .Y(n24553) );
  XNOR2X1 U48766 ( .A(n50816), .B(n41297), .Y(n24522) );
  XNOR2X1 U48767 ( .A(n50815), .B(n41293), .Y(n24532) );
  XNOR2X1 U48768 ( .A(n50853), .B(n41294), .Y(n24382) );
  XNOR2X1 U48769 ( .A(n50849), .B(n41292), .Y(n24492) );
  XNOR2X1 U48770 ( .A(n50813), .B(n41293), .Y(n24502) );
  XNOR2X1 U48771 ( .A(n50814), .B(n41292), .Y(n24512) );
  XNOR2X1 U48772 ( .A(n50848), .B(n36789), .Y(n21938) );
  XNOR2X1 U48773 ( .A(n50852), .B(n42539), .Y(n30114) );
  XNOR2X1 U48774 ( .A(n50849), .B(n42540), .Y(n30174) );
  XNOR2X1 U48775 ( .A(n50848), .B(n42539), .Y(n30054) );
  XNOR2X1 U48776 ( .A(n50845), .B(n42542), .Y(n29964) );
  XNOR2X1 U48777 ( .A(n50847), .B(n42540), .Y(n30024) );
  XNOR2X1 U48778 ( .A(n50844), .B(n42539), .Y(n29754) );
  XNOR2X1 U48779 ( .A(n50846), .B(n42533), .Y(n29994) );
  XNOR2X1 U48780 ( .A(n50841), .B(n42537), .Y(n29784) );
  XNOR2X1 U48781 ( .A(n50842), .B(n42540), .Y(n29814) );
  XNOR2X1 U48782 ( .A(n50834), .B(n42544), .Y(n29513) );
  XNOR2X1 U48783 ( .A(n50833), .B(n42539), .Y(n29483) );
  XNOR2X1 U48784 ( .A(n50832), .B(n42541), .Y(n29603) );
  XNOR2X1 U48785 ( .A(n50851), .B(n42540), .Y(n30084) );
  XNOR2X1 U48786 ( .A(n50850), .B(n42542), .Y(n30144) );
  XNOR2X1 U48787 ( .A(n50828), .B(n42542), .Y(n26143) );
  XNOR2X1 U48788 ( .A(n50826), .B(n42537), .Y(n26083) );
  XNOR2X1 U48789 ( .A(n50843), .B(n42543), .Y(n29724) );
  XNOR2X1 U48790 ( .A(n50825), .B(n42534), .Y(n26053) );
  XNOR2X1 U48791 ( .A(n50820), .B(n42537), .Y(n25813) );
  XNOR2X1 U48792 ( .A(n50822), .B(n42534), .Y(n25993) );
  XNOR2X1 U48793 ( .A(n50824), .B(n42537), .Y(n25933) );
  XNOR2X1 U48794 ( .A(n50838), .B(n42539), .Y(n29844) );
  XNOR2X1 U48795 ( .A(n50854), .B(n42540), .Y(n30325) );
  XNOR2X1 U48796 ( .A(n50853), .B(n42541), .Y(n30355) );
  XNOR2X1 U48797 ( .A(n50823), .B(n42538), .Y(n25963) );
  XNOR2X1 U48798 ( .A(n50821), .B(n42534), .Y(n26023) );
  XNOR2X1 U48799 ( .A(n50827), .B(n42535), .Y(n26113) );
  XNOR2X1 U48800 ( .A(n50837), .B(n42541), .Y(n29904) );
  XNOR2X1 U48801 ( .A(n50839), .B(n42533), .Y(n29874) );
  XNOR2X1 U48802 ( .A(n50840), .B(n42542), .Y(n29934) );
  XNOR2X1 U48803 ( .A(n50819), .B(n42534), .Y(n25843) );
  XNOR2X1 U48804 ( .A(n50835), .B(n42540), .Y(n29543) );
  XNOR2X1 U48805 ( .A(n50836), .B(n42537), .Y(n29573) );
  XNOR2X1 U48806 ( .A(n50808), .B(n42532), .Y(n26323) );
  XNOR2X1 U48807 ( .A(n50809), .B(n42532), .Y(n26173) );
  XNOR2X1 U48808 ( .A(n50830), .B(n42544), .Y(n29663) );
  XNOR2X1 U48809 ( .A(n50829), .B(n42536), .Y(n29693) );
  XNOR2X1 U48810 ( .A(n50831), .B(n42536), .Y(n29633) );
  XNOR2X1 U48811 ( .A(n50812), .B(n42532), .Y(n26263) );
  XNOR2X1 U48812 ( .A(n50818), .B(n42534), .Y(n25903) );
  XNOR2X1 U48813 ( .A(n50817), .B(n42534), .Y(n25873) );
  XNOR2X1 U48814 ( .A(n50811), .B(n42532), .Y(n26233) );
  XNOR2X1 U48815 ( .A(n50810), .B(n42532), .Y(n26203) );
  XNOR2X1 U48816 ( .A(n50814), .B(n42538), .Y(n25783) );
  XNOR2X1 U48817 ( .A(n50803), .B(n42532), .Y(n26504) );
  XNOR2X1 U48818 ( .A(n50804), .B(n42532), .Y(n26474) );
  XNOR2X1 U48819 ( .A(n50807), .B(n42532), .Y(n26293) );
  XNOR2X1 U48820 ( .A(n50805), .B(n42532), .Y(n26353) );
  XNOR2X1 U48821 ( .A(n50806), .B(n42532), .Y(n26383) );
  XNOR2X1 U48822 ( .A(n50798), .B(n42532), .Y(n26534) );
  XNOR2X1 U48823 ( .A(n50801), .B(n42532), .Y(n26414) );
  XNOR2X1 U48824 ( .A(n50802), .B(n42532), .Y(n26444) );
  XNOR2X1 U48825 ( .A(n51270), .B(n42694), .Y(n29958) );
  XNOR2X1 U48826 ( .A(n51040), .B(n36715), .Y(n20924) );
  XNOR2X1 U48827 ( .A(n51034), .B(n36722), .Y(n20851) );
  XNOR2X1 U48828 ( .A(n51038), .B(n36716), .Y(n20883) );
  XNOR2X1 U48829 ( .A(n51032), .B(n36717), .Y(n20871) );
  XNOR2X1 U48830 ( .A(n51031), .B(n36721), .Y(n20861) );
  XNOR2X1 U48831 ( .A(n51029), .B(n36722), .Y(n20808) );
  XNOR2X1 U48832 ( .A(n51028), .B(n36717), .Y(n20829) );
  XNOR2X1 U48833 ( .A(n51027), .B(n36721), .Y(n20819) );
  XNOR2X1 U48834 ( .A(n51073), .B(n41328), .Y(n24453) );
  XNOR2X1 U48835 ( .A(n51073), .B(n36718), .Y(n22059) );
  XNOR2X1 U48836 ( .A(n51072), .B(n41331), .Y(n24443) );
  XNOR2X1 U48837 ( .A(n51074), .B(n36721), .Y(n22069) );
  XNOR2X1 U48838 ( .A(n51072), .B(n36717), .Y(n22049) );
  XNOR2X1 U48839 ( .A(n51069), .B(n41331), .Y(n24403) );
  XNOR2X1 U48840 ( .A(n51071), .B(n36715), .Y(n22039) );
  XNOR2X1 U48841 ( .A(n51068), .B(n41333), .Y(n24393) );
  XNOR2X1 U48842 ( .A(n51065), .B(n41332), .Y(n24473) );
  XNOR2X1 U48843 ( .A(n51064), .B(n41329), .Y(n24463) );
  XNOR2X1 U48844 ( .A(n51064), .B(n36717), .Y(n21989) );
  XNOR2X1 U48845 ( .A(n51063), .B(n36722), .Y(n21979) );
  XNOR2X1 U48846 ( .A(n51061), .B(n36717), .Y(n21949) );
  XNOR2X1 U48847 ( .A(n51058), .B(n41330), .Y(n24271) );
  XNOR2X1 U48848 ( .A(n51070), .B(n41330), .Y(n24423) );
  XNOR2X1 U48849 ( .A(n51060), .B(n36720), .Y(n21969) );
  XNOR2X1 U48850 ( .A(n51057), .B(n41330), .Y(n24261) );
  XNOR2X1 U48851 ( .A(n51071), .B(n41330), .Y(n24433) );
  XNOR2X1 U48852 ( .A(n51059), .B(n36718), .Y(n21959) );
  XNOR2X1 U48853 ( .A(n51056), .B(n41328), .Y(n24251) );
  XNOR2X1 U48854 ( .A(n51054), .B(n41331), .Y(n24291) );
  XNOR2X1 U48855 ( .A(n51066), .B(n41332), .Y(n24483) );
  XNOR2X1 U48856 ( .A(n51060), .B(n41332), .Y(n24351) );
  XNOR2X1 U48857 ( .A(n51059), .B(n41331), .Y(n24341) );
  XNOR2X1 U48858 ( .A(n51052), .B(n41330), .Y(n24241) );
  XNOR2X1 U48859 ( .A(n51053), .B(n36715), .Y(n21857) );
  XNOR2X1 U48860 ( .A(n51062), .B(n41331), .Y(n24371) );
  XNOR2X1 U48861 ( .A(n51061), .B(n41333), .Y(n24361) );
  XNOR2X1 U48862 ( .A(n51070), .B(n36718), .Y(n22019) );
  XNOR2X1 U48863 ( .A(n51069), .B(n36715), .Y(n22029) );
  XNOR2X1 U48864 ( .A(n51065), .B(n36718), .Y(n21999) );
  XNOR2X1 U48865 ( .A(n51066), .B(n36722), .Y(n22009) );
  XNOR2X1 U48866 ( .A(n51055), .B(n41333), .Y(n24281) );
  XNOR2X1 U48867 ( .A(n51049), .B(n36718), .Y(n21908) );
  XNOR2X1 U48868 ( .A(n51046), .B(n41327), .Y(n24331) );
  XNOR2X1 U48869 ( .A(n51050), .B(n36718), .Y(n21827) );
  XNOR2X1 U48870 ( .A(n51048), .B(n36722), .Y(n21929) );
  XNOR2X1 U48871 ( .A(n51045), .B(n41331), .Y(n24321) );
  XNOR2X1 U48872 ( .A(n51047), .B(n36715), .Y(n21919) );
  XNOR2X1 U48873 ( .A(n51045), .B(n36721), .Y(n21888) );
  XNOR2X1 U48874 ( .A(n51044), .B(n41328), .Y(n24301) );
  XNOR2X1 U48875 ( .A(n51043), .B(n41332), .Y(n24311) );
  XNOR2X1 U48876 ( .A(n51054), .B(n36716), .Y(n21817) );
  XNOR2X1 U48877 ( .A(n51051), .B(n36721), .Y(n21837) );
  XNOR2X1 U48878 ( .A(n51052), .B(n36714), .Y(n21847) );
  XNOR2X1 U48879 ( .A(n51042), .B(n41327), .Y(n24605) );
  XNOR2X1 U48880 ( .A(n51041), .B(n41329), .Y(n24615) );
  XNOR2X1 U48881 ( .A(n51046), .B(n36716), .Y(n21898) );
  XNOR2X1 U48882 ( .A(n51044), .B(n36720), .Y(n21868) );
  XNOR2X1 U48883 ( .A(n51039), .B(n41332), .Y(n24585) );
  XNOR2X1 U48884 ( .A(n51040), .B(n41330), .Y(n24595) );
  XNOR2X1 U48885 ( .A(n51043), .B(n36714), .Y(n21878) );
  XNOR2X1 U48886 ( .A(n51038), .B(n41328), .Y(n24565) );
  XNOR2X1 U48887 ( .A(n51035), .B(n41327), .Y(n24575) );
  XNOR2X1 U48888 ( .A(n51031), .B(n41332), .Y(n24625) );
  XNOR2X1 U48889 ( .A(n51037), .B(n41333), .Y(n24543) );
  XNOR2X1 U48890 ( .A(n51036), .B(n41329), .Y(n24554) );
  XNOR2X1 U48891 ( .A(n51030), .B(n41333), .Y(n24523) );
  XNOR2X1 U48892 ( .A(n51029), .B(n41331), .Y(n24533) );
  XNOR2X1 U48893 ( .A(n51067), .B(n41330), .Y(n24383) );
  XNOR2X1 U48894 ( .A(n51063), .B(n41327), .Y(n24493) );
  XNOR2X1 U48895 ( .A(n51027), .B(n41331), .Y(n24503) );
  XNOR2X1 U48896 ( .A(n51028), .B(n41331), .Y(n24513) );
  XNOR2X1 U48897 ( .A(n51062), .B(n36717), .Y(n21939) );
  XNOR2X1 U48898 ( .A(n51281), .B(n36867), .Y(n30130) );
  XNOR2X1 U48899 ( .A(n50639), .B(n42587), .Y(n30126) );
  XNOR2X1 U48900 ( .A(n50636), .B(n42587), .Y(n30186) );
  XNOR2X1 U48901 ( .A(n51066), .B(n42552), .Y(n30115) );
  XNOR2X1 U48902 ( .A(n51277), .B(n36867), .Y(n30070) );
  XNOR2X1 U48903 ( .A(n50635), .B(n42587), .Y(n30066) );
  XNOR2X1 U48904 ( .A(n51063), .B(n42548), .Y(n30175) );
  XNOR2X1 U48905 ( .A(n51062), .B(n42552), .Y(n30055) );
  XNOR2X1 U48906 ( .A(n51280), .B(n36867), .Y(n30100) );
  XNOR2X1 U48907 ( .A(n50638), .B(n42587), .Y(n30096) );
  XNOR2X1 U48908 ( .A(n51059), .B(n42552), .Y(n29965) );
  XNOR2X1 U48909 ( .A(n51061), .B(n42553), .Y(n30025) );
  XNOR2X1 U48910 ( .A(n51060), .B(n42552), .Y(n29995) );
  XNOR2X1 U48911 ( .A(n51269), .B(n36867), .Y(n29950) );
  XNOR2X1 U48912 ( .A(n50627), .B(n42587), .Y(n29946) );
  XNOR2X1 U48913 ( .A(n51267), .B(n36867), .Y(n29860) );
  XNOR2X1 U48914 ( .A(n50625), .B(n42587), .Y(n29856) );
  XNOR2X1 U48915 ( .A(n50616), .B(net219460), .Y(n26163) );
  XNOR2X1 U48916 ( .A(n51257), .B(n42637), .Y(n26159) );
  XNOR2X1 U48917 ( .A(n50615), .B(n42589), .Y(n26155) );
  XNOR2X1 U48918 ( .A(n51065), .B(n42553), .Y(n30085) );
  XNOR2X1 U48919 ( .A(n50613), .B(net219434), .Y(n26073) );
  XNOR2X1 U48920 ( .A(n51254), .B(n42637), .Y(n26069) );
  XNOR2X1 U48921 ( .A(n50612), .B(n42588), .Y(n26065) );
  XNOR2X1 U48922 ( .A(n50610), .B(net219434), .Y(n26013) );
  XNOR2X1 U48923 ( .A(n51251), .B(n42637), .Y(n26009) );
  XNOR2X1 U48924 ( .A(n50609), .B(n42588), .Y(n26005) );
  XNOR2X1 U48925 ( .A(n51064), .B(n42553), .Y(n30145) );
  XNOR2X1 U48926 ( .A(n51042), .B(n42547), .Y(n26144) );
  XNOR2X1 U48927 ( .A(n51040), .B(n42552), .Y(n26084) );
  XNOR2X1 U48928 ( .A(n50612), .B(net258207), .Y(n25953) );
  XNOR2X1 U48929 ( .A(n51253), .B(n42637), .Y(n25949) );
  XNOR2X1 U48930 ( .A(n50611), .B(n42592), .Y(n25945) );
  XNOR2X1 U48931 ( .A(n51039), .B(n42548), .Y(n26054) );
  XNOR2X1 U48932 ( .A(n51034), .B(n42554), .Y(n25814) );
  XNOR2X1 U48933 ( .A(n51036), .B(n42550), .Y(n25994) );
  XNOR2X1 U48934 ( .A(n51268), .B(n36867), .Y(n29890) );
  XNOR2X1 U48935 ( .A(n50626), .B(n42587), .Y(n29886) );
  XNOR2X1 U48936 ( .A(n50611), .B(net219434), .Y(n25983) );
  XNOR2X1 U48937 ( .A(n51252), .B(n42638), .Y(n25979) );
  XNOR2X1 U48938 ( .A(n50610), .B(n42592), .Y(n25975) );
  XNOR2X1 U48939 ( .A(n50609), .B(net258207), .Y(n26043) );
  XNOR2X1 U48940 ( .A(n51250), .B(n42637), .Y(n26039) );
  XNOR2X1 U48941 ( .A(n50608), .B(n42588), .Y(n26035) );
  XNOR2X1 U48942 ( .A(n51038), .B(n42552), .Y(n25934) );
  XNOR2X1 U48943 ( .A(n51052), .B(n42553), .Y(n29845) );
  XNOR2X1 U48944 ( .A(n51256), .B(n42637), .Y(n26129) );
  XNOR2X1 U48945 ( .A(n50614), .B(n42592), .Y(n26125) );
  XNOR2X1 U48946 ( .A(n51068), .B(n42551), .Y(n30326) );
  XNOR2X1 U48947 ( .A(n51067), .B(n42551), .Y(n30356) );
  XNOR2X1 U48948 ( .A(n51037), .B(n42546), .Y(n25964) );
  XNOR2X1 U48949 ( .A(n51035), .B(n42552), .Y(n26024) );
  XNOR2X1 U48950 ( .A(n51255), .B(n42637), .Y(n26099) );
  XNOR2X1 U48951 ( .A(n50613), .B(n42586), .Y(n26095) );
  XNOR2X1 U48952 ( .A(n51041), .B(n42552), .Y(n26114) );
  XNOR2X1 U48953 ( .A(n50597), .B(net219460), .Y(n26193) );
  XNOR2X1 U48954 ( .A(n51238), .B(n36867), .Y(n26189) );
  XNOR2X1 U48955 ( .A(n50596), .B(n36863), .Y(n26185) );
  XNOR2X1 U48956 ( .A(n51051), .B(n42552), .Y(n29905) );
  XNOR2X1 U48957 ( .A(n51053), .B(n42552), .Y(n29875) );
  XNOR2X1 U48958 ( .A(n51054), .B(n42546), .Y(n29935) );
  XNOR2X1 U48959 ( .A(n51033), .B(n42554), .Y(n25844) );
  XNOR2X1 U48960 ( .A(n51249), .B(n42637), .Y(n25829) );
  XNOR2X1 U48961 ( .A(n50607), .B(n36863), .Y(n25825) );
  XNOR2X1 U48962 ( .A(n50600), .B(net219460), .Y(n26283) );
  XNOR2X1 U48963 ( .A(n51241), .B(n36867), .Y(n26279) );
  XNOR2X1 U48964 ( .A(n50599), .B(n42589), .Y(n26275) );
  XNOR2X1 U48965 ( .A(n50605), .B(net219460), .Y(n25893) );
  XNOR2X1 U48966 ( .A(n51022), .B(n42546), .Y(n26324) );
  XNOR2X1 U48967 ( .A(n51023), .B(n42546), .Y(n26174) );
  XNOR2X1 U48968 ( .A(n51247), .B(n42637), .Y(n25919) );
  XNOR2X1 U48969 ( .A(n50605), .B(n42588), .Y(n25915) );
  XNOR2X1 U48970 ( .A(n50607), .B(net219444), .Y(n25863) );
  XNOR2X1 U48971 ( .A(n51248), .B(n42637), .Y(n25859) );
  XNOR2X1 U48972 ( .A(n50606), .B(n42592), .Y(n25855) );
  XNOR2X1 U48973 ( .A(n50604), .B(net219460), .Y(n25743) );
  XNOR2X1 U48974 ( .A(n51026), .B(n42546), .Y(n26264) );
  XNOR2X1 U48975 ( .A(n51032), .B(n42546), .Y(n25904) );
  XNOR2X1 U48976 ( .A(n51031), .B(n42552), .Y(n25874) );
  XNOR2X1 U48977 ( .A(n50601), .B(net219444), .Y(n25773) );
  XNOR2X1 U48978 ( .A(n51242), .B(n42637), .Y(n25769) );
  XNOR2X1 U48979 ( .A(n50600), .B(n42592), .Y(n25765) );
  XNOR2X1 U48980 ( .A(n51025), .B(n42546), .Y(n26234) );
  XNOR2X1 U48981 ( .A(n51024), .B(n42546), .Y(n26204) );
  XNOR2X1 U48982 ( .A(n50598), .B(net219460), .Y(n26223) );
  XNOR2X1 U48983 ( .A(n51239), .B(n36867), .Y(n26219) );
  XNOR2X1 U48984 ( .A(n50597), .B(n42586), .Y(n26215) );
  XNOR2X1 U48985 ( .A(n50599), .B(net219460), .Y(n26253) );
  XNOR2X1 U48986 ( .A(n51240), .B(n36867), .Y(n26249) );
  XNOR2X1 U48987 ( .A(n50598), .B(n42589), .Y(n26245) );
  XNOR2X1 U48988 ( .A(n50591), .B(net219460), .Y(n26524) );
  XNOR2X1 U48989 ( .A(n51232), .B(n36867), .Y(n26520) );
  XNOR2X1 U48990 ( .A(n50590), .B(n42591), .Y(n26516) );
  XNOR2X1 U48991 ( .A(n50592), .B(net219460), .Y(n26494) );
  XNOR2X1 U48992 ( .A(n51233), .B(n36867), .Y(n26490) );
  XNOR2X1 U48993 ( .A(n50591), .B(n42586), .Y(n26486) );
  XNOR2X1 U48994 ( .A(n50602), .B(net258207), .Y(n25803) );
  XNOR2X1 U48995 ( .A(n51243), .B(n42637), .Y(n25799) );
  XNOR2X1 U48996 ( .A(n50601), .B(n42592), .Y(n25795) );
  XNOR2X1 U48997 ( .A(n51027), .B(n42546), .Y(n25754) );
  XNOR2X1 U48998 ( .A(n51028), .B(n42552), .Y(n25784) );
  XNOR2X1 U48999 ( .A(n50593), .B(net219460), .Y(n26373) );
  XNOR2X1 U49000 ( .A(n51234), .B(n36867), .Y(n26369) );
  XNOR2X1 U49001 ( .A(n50592), .B(n42586), .Y(n26365) );
  XNOR2X1 U49002 ( .A(n51235), .B(n42637), .Y(n26399) );
  XNOR2X1 U49003 ( .A(n50593), .B(n42586), .Y(n26395) );
  XNOR2X1 U49004 ( .A(n50594), .B(net219460), .Y(n26403) );
  XNOR2X1 U49005 ( .A(n51017), .B(n42546), .Y(n26505) );
  XNOR2X1 U49006 ( .A(n51018), .B(n42546), .Y(n26475) );
  XNOR2X1 U49007 ( .A(n51227), .B(n36867), .Y(n26550) );
  XNOR2X1 U49008 ( .A(n50585), .B(n42586), .Y(n26546) );
  XNOR2X1 U49009 ( .A(n51021), .B(n42546), .Y(n26294) );
  XNOR2X1 U49010 ( .A(n50596), .B(net219460), .Y(n26343) );
  XNOR2X1 U49011 ( .A(n51237), .B(n36867), .Y(n26339) );
  XNOR2X1 U49012 ( .A(n50595), .B(n36863), .Y(n26335) );
  XNOR2X1 U49013 ( .A(n50589), .B(net219460), .Y(n26434) );
  XNOR2X1 U49014 ( .A(n51230), .B(n42638), .Y(n26430) );
  XNOR2X1 U49015 ( .A(n50588), .B(n36863), .Y(n26426) );
  XNOR2X1 U49016 ( .A(n51019), .B(n42547), .Y(n26354) );
  XNOR2X1 U49017 ( .A(n51020), .B(n42546), .Y(n26384) );
  XNOR2X1 U49018 ( .A(n50595), .B(net219460), .Y(n26313) );
  XNOR2X1 U49019 ( .A(n51236), .B(n42638), .Y(n26309) );
  XNOR2X1 U49020 ( .A(n50594), .B(n42588), .Y(n26305) );
  XNOR2X1 U49021 ( .A(n51015), .B(n42546), .Y(n26415) );
  XNOR2X1 U49022 ( .A(n51016), .B(n42546), .Y(n26445) );
  XNOR2X1 U49023 ( .A(n50590), .B(net219460), .Y(n26464) );
  XNOR2X1 U49024 ( .A(n51231), .B(n42637), .Y(n26460) );
  XNOR2X1 U49025 ( .A(n50589), .B(n42589), .Y(n26456) );
  XNOR2X1 U49026 ( .A(n50437), .B(n42717), .Y(n30137) );
  XNOR2X1 U49027 ( .A(n50433), .B(n42717), .Y(n30077) );
  XNOR2X1 U49028 ( .A(n50425), .B(n42724), .Y(n29957) );
  XNOR2X1 U49029 ( .A(n50423), .B(n42719), .Y(n29867) );
  XNOR2X1 U49030 ( .A(n50424), .B(n42719), .Y(n29897) );
  XNOR2X1 U49031 ( .A(n50612), .B(n42463), .Y(n20925) );
  XNOR2X1 U49032 ( .A(n50606), .B(n42464), .Y(n20852) );
  XNOR2X1 U49033 ( .A(n50610), .B(n42464), .Y(n20884) );
  XNOR2X1 U49034 ( .A(n50604), .B(n42463), .Y(n20872) );
  XNOR2X1 U49035 ( .A(n50603), .B(n42463), .Y(n20862) );
  XNOR2X1 U49036 ( .A(n50601), .B(n42463), .Y(n20809) );
  XNOR2X1 U49037 ( .A(n50600), .B(n42464), .Y(n20830) );
  XNOR2X1 U49038 ( .A(n50599), .B(n42464), .Y(n20820) );
  XNOR2X1 U49039 ( .A(n50645), .B(n36850), .Y(n24454) );
  XNOR2X1 U49040 ( .A(n50645), .B(n42464), .Y(n22060) );
  XNOR2X1 U49041 ( .A(n50644), .B(n36856), .Y(n24444) );
  XNOR2X1 U49042 ( .A(n50646), .B(n42464), .Y(n22070) );
  XNOR2X1 U49043 ( .A(n50644), .B(n42464), .Y(n22050) );
  XNOR2X1 U49044 ( .A(n50641), .B(n36851), .Y(n24404) );
  XNOR2X1 U49045 ( .A(n50643), .B(n42464), .Y(n22040) );
  XNOR2X1 U49046 ( .A(n50640), .B(n36858), .Y(n24394) );
  XNOR2X1 U49047 ( .A(n50637), .B(n36851), .Y(n24474) );
  XNOR2X1 U49048 ( .A(n50636), .B(n36851), .Y(n24464) );
  XNOR2X1 U49049 ( .A(n50636), .B(n42464), .Y(n21990) );
  XNOR2X1 U49050 ( .A(n50635), .B(n42464), .Y(n21980) );
  XNOR2X1 U49051 ( .A(n50633), .B(n42464), .Y(n21950) );
  XNOR2X1 U49052 ( .A(n50630), .B(n36850), .Y(n24272) );
  XNOR2X1 U49053 ( .A(n50642), .B(n36854), .Y(n24424) );
  XNOR2X1 U49054 ( .A(n50632), .B(n42464), .Y(n21970) );
  XNOR2X1 U49055 ( .A(n50629), .B(n36857), .Y(n24262) );
  XNOR2X1 U49056 ( .A(n50643), .B(n36852), .Y(n24434) );
  XNOR2X1 U49057 ( .A(n50631), .B(n42464), .Y(n21960) );
  XNOR2X1 U49058 ( .A(n50628), .B(n36857), .Y(n24252) );
  XNOR2X1 U49059 ( .A(n50626), .B(n36857), .Y(n24292) );
  XNOR2X1 U49060 ( .A(n50638), .B(n36853), .Y(n24484) );
  XNOR2X1 U49061 ( .A(n50632), .B(n36858), .Y(n24352) );
  XNOR2X1 U49062 ( .A(n50631), .B(n36851), .Y(n24342) );
  XNOR2X1 U49063 ( .A(n50624), .B(n36856), .Y(n24242) );
  XNOR2X1 U49064 ( .A(n50625), .B(n42463), .Y(n21858) );
  XNOR2X1 U49065 ( .A(n50634), .B(n36859), .Y(n24372) );
  XNOR2X1 U49066 ( .A(n50633), .B(n36857), .Y(n24362) );
  XNOR2X1 U49067 ( .A(n50642), .B(n42464), .Y(n22020) );
  XNOR2X1 U49068 ( .A(n50641), .B(n42464), .Y(n22030) );
  XNOR2X1 U49069 ( .A(n50637), .B(n42464), .Y(n22000) );
  XNOR2X1 U49070 ( .A(n50638), .B(n42464), .Y(n22010) );
  XNOR2X1 U49071 ( .A(n50627), .B(n36860), .Y(n24282) );
  XNOR2X1 U49072 ( .A(n50621), .B(n42463), .Y(n21909) );
  XNOR2X1 U49073 ( .A(n50618), .B(n36858), .Y(n24332) );
  XNOR2X1 U49074 ( .A(n50622), .B(n42463), .Y(n21828) );
  XNOR2X1 U49075 ( .A(n50620), .B(n42463), .Y(n21930) );
  XNOR2X1 U49076 ( .A(n50617), .B(n36856), .Y(n24322) );
  XNOR2X1 U49077 ( .A(n50619), .B(n42463), .Y(n21920) );
  XNOR2X1 U49078 ( .A(n50617), .B(n42463), .Y(n21889) );
  XNOR2X1 U49079 ( .A(n50616), .B(n36859), .Y(n24302) );
  XNOR2X1 U49080 ( .A(n50615), .B(n36859), .Y(n24312) );
  XNOR2X1 U49081 ( .A(n50626), .B(n42463), .Y(n21818) );
  XNOR2X1 U49082 ( .A(n50623), .B(n42463), .Y(n21838) );
  XNOR2X1 U49083 ( .A(n50624), .B(n42463), .Y(n21848) );
  XNOR2X1 U49084 ( .A(n50614), .B(n36860), .Y(n24606) );
  XNOR2X1 U49085 ( .A(n50613), .B(n36853), .Y(n24616) );
  XNOR2X1 U49086 ( .A(n50618), .B(n42463), .Y(n21899) );
  XNOR2X1 U49087 ( .A(n50616), .B(n42463), .Y(n21869) );
  XNOR2X1 U49088 ( .A(n50611), .B(n36852), .Y(n24586) );
  XNOR2X1 U49089 ( .A(n50612), .B(n36852), .Y(n24596) );
  XNOR2X1 U49090 ( .A(n50615), .B(n42463), .Y(n21879) );
  XNOR2X1 U49091 ( .A(n50610), .B(n36856), .Y(n24566) );
  XNOR2X1 U49092 ( .A(n50607), .B(n36857), .Y(n24576) );
  XNOR2X1 U49093 ( .A(n50603), .B(n36850), .Y(n24626) );
  XNOR2X1 U49094 ( .A(n50609), .B(n36852), .Y(n24544) );
  XNOR2X1 U49095 ( .A(n50608), .B(n36853), .Y(n24555) );
  XNOR2X1 U49096 ( .A(n50602), .B(n36856), .Y(n24524) );
  XNOR2X1 U49097 ( .A(n50601), .B(n36854), .Y(n24534) );
  XNOR2X1 U49098 ( .A(n50639), .B(n36859), .Y(n24384) );
  XNOR2X1 U49099 ( .A(n50635), .B(n36854), .Y(n24494) );
  XNOR2X1 U49100 ( .A(n50599), .B(n36852), .Y(n24504) );
  XNOR2X1 U49101 ( .A(n50600), .B(n36853), .Y(n24514) );
  XNOR2X1 U49102 ( .A(n50634), .B(n42463), .Y(n21940) );
  XNOR2X1 U49103 ( .A(n50222), .B(n42704), .Y(n30136) );
  XNOR2X1 U49104 ( .A(n50221), .B(n42675), .Y(n30128) );
  XNOR2X1 U49105 ( .A(n50853), .B(n42618), .Y(n30124) );
  XNOR2X1 U49106 ( .A(n50218), .B(n42675), .Y(n30188) );
  XNOR2X1 U49107 ( .A(n50850), .B(n42619), .Y(n30184) );
  XNOR2X1 U49108 ( .A(n50218), .B(n42704), .Y(n30076) );
  XNOR2X1 U49109 ( .A(n50217), .B(n42674), .Y(n30068) );
  XNOR2X1 U49110 ( .A(n50849), .B(n42620), .Y(n30064) );
  XNOR2X1 U49111 ( .A(n50221), .B(n42708), .Y(n30106) );
  XNOR2X1 U49112 ( .A(n50220), .B(n42671), .Y(n30098) );
  XNOR2X1 U49113 ( .A(n50852), .B(n42620), .Y(n30094) );
  XNOR2X1 U49114 ( .A(n50851), .B(n42615), .Y(n30154) );
  XNOR2X1 U49115 ( .A(n50210), .B(n42710), .Y(n29956) );
  XNOR2X1 U49116 ( .A(n50209), .B(n42675), .Y(n29948) );
  XNOR2X1 U49117 ( .A(n50841), .B(n42615), .Y(n29944) );
  XNOR2X1 U49118 ( .A(n50208), .B(n42711), .Y(n29866) );
  XNOR2X1 U49119 ( .A(n50207), .B(n42675), .Y(n29858) );
  XNOR2X1 U49120 ( .A(n50839), .B(n42615), .Y(n29854) );
  XNOR2X1 U49121 ( .A(n50830), .B(net219310), .Y(n26161) );
  XNOR2X1 U49122 ( .A(n50197), .B(n42669), .Y(n26157) );
  XNOR2X1 U49123 ( .A(n50829), .B(n41284), .Y(n26153) );
  XNOR2X1 U49124 ( .A(n50827), .B(net219310), .Y(n26071) );
  XNOR2X1 U49125 ( .A(n50194), .B(n42676), .Y(n26067) );
  XNOR2X1 U49126 ( .A(n50826), .B(n42619), .Y(n26063) );
  XNOR2X1 U49127 ( .A(n50824), .B(n40039), .Y(n26011) );
  XNOR2X1 U49128 ( .A(n50191), .B(n42671), .Y(n26007) );
  XNOR2X1 U49129 ( .A(n50823), .B(n42615), .Y(n26003) );
  XNOR2X1 U49130 ( .A(n50826), .B(net219314), .Y(n25951) );
  XNOR2X1 U49131 ( .A(n50193), .B(n42669), .Y(n25947) );
  XNOR2X1 U49132 ( .A(n50825), .B(n42618), .Y(n25943) );
  XNOR2X1 U49133 ( .A(n50209), .B(n42711), .Y(n29896) );
  XNOR2X1 U49134 ( .A(n50208), .B(n42675), .Y(n29888) );
  XNOR2X1 U49135 ( .A(n50840), .B(n42615), .Y(n29884) );
  XNOR2X1 U49136 ( .A(n50825), .B(net219310), .Y(n25981) );
  XNOR2X1 U49137 ( .A(n50192), .B(n42676), .Y(n25977) );
  XNOR2X1 U49138 ( .A(n50824), .B(n42619), .Y(n25973) );
  XNOR2X1 U49139 ( .A(n50823), .B(net219330), .Y(n26041) );
  XNOR2X1 U49140 ( .A(n50190), .B(n42671), .Y(n26037) );
  XNOR2X1 U49141 ( .A(n50822), .B(n42615), .Y(n26033) );
  XNOR2X1 U49142 ( .A(n50829), .B(net219310), .Y(n26131) );
  XNOR2X1 U49143 ( .A(n50196), .B(n42676), .Y(n26127) );
  XNOR2X1 U49144 ( .A(n50828), .B(n42615), .Y(n26123) );
  XNOR2X1 U49145 ( .A(n50195), .B(n42672), .Y(n26097) );
  XNOR2X1 U49146 ( .A(n50827), .B(n42615), .Y(n26093) );
  XNOR2X1 U49147 ( .A(n50811), .B(net219336), .Y(n26191) );
  XNOR2X1 U49148 ( .A(n50178), .B(n42673), .Y(n26187) );
  XNOR2X1 U49149 ( .A(n50810), .B(n42618), .Y(n26183) );
  XNOR2X1 U49150 ( .A(n50189), .B(n34444), .Y(n25827) );
  XNOR2X1 U49151 ( .A(n50821), .B(n42614), .Y(n25823) );
  XNOR2X1 U49152 ( .A(n50181), .B(n42673), .Y(n26277) );
  XNOR2X1 U49153 ( .A(n50813), .B(n42619), .Y(n26273) );
  XNOR2X1 U49154 ( .A(n50819), .B(net219308), .Y(n25891) );
  XNOR2X1 U49155 ( .A(n50186), .B(n42671), .Y(n25887) );
  XNOR2X1 U49156 ( .A(n50818), .B(n42613), .Y(n25883) );
  XNOR2X1 U49157 ( .A(n50820), .B(n40039), .Y(n25921) );
  XNOR2X1 U49158 ( .A(n50187), .B(n42669), .Y(n25917) );
  XNOR2X1 U49159 ( .A(n50819), .B(n42613), .Y(n25913) );
  XNOR2X1 U49160 ( .A(n50821), .B(net258262), .Y(n25861) );
  XNOR2X1 U49161 ( .A(n50815), .B(net219330), .Y(n25771) );
  XNOR2X1 U49162 ( .A(n50182), .B(n42671), .Y(n25767) );
  XNOR2X1 U49163 ( .A(n50814), .B(n42618), .Y(n25763) );
  XNOR2X1 U49164 ( .A(n50812), .B(net219336), .Y(n26221) );
  XNOR2X1 U49165 ( .A(n50179), .B(n42673), .Y(n26217) );
  XNOR2X1 U49166 ( .A(n50811), .B(n42615), .Y(n26213) );
  XNOR2X1 U49167 ( .A(n50813), .B(n40039), .Y(n26251) );
  XNOR2X1 U49168 ( .A(n50180), .B(n42673), .Y(n26247) );
  XNOR2X1 U49169 ( .A(n50812), .B(n42618), .Y(n26243) );
  XNOR2X1 U49170 ( .A(n50805), .B(net219336), .Y(n26522) );
  XNOR2X1 U49171 ( .A(n50172), .B(n42673), .Y(n26518) );
  XNOR2X1 U49172 ( .A(n50804), .B(n42618), .Y(n26514) );
  XNOR2X1 U49173 ( .A(n50806), .B(n40039), .Y(n26492) );
  XNOR2X1 U49174 ( .A(n50173), .B(n42673), .Y(n26488) );
  XNOR2X1 U49175 ( .A(n50805), .B(n42615), .Y(n26484) );
  XNOR2X1 U49176 ( .A(n50816), .B(net219310), .Y(n25801) );
  XNOR2X1 U49177 ( .A(n50183), .B(n42669), .Y(n25797) );
  XNOR2X1 U49178 ( .A(n50815), .B(n36868), .Y(n25793) );
  XNOR2X1 U49179 ( .A(n50807), .B(net219308), .Y(n26371) );
  XNOR2X1 U49180 ( .A(n50174), .B(n42673), .Y(n26367) );
  XNOR2X1 U49181 ( .A(n50806), .B(n42618), .Y(n26363) );
  XNOR2X1 U49182 ( .A(n50175), .B(n42673), .Y(n26397) );
  XNOR2X1 U49183 ( .A(n50807), .B(n42618), .Y(n26393) );
  XNOR2X1 U49184 ( .A(n50808), .B(n36870), .Y(n26401) );
  XNOR2X1 U49185 ( .A(n50167), .B(n42673), .Y(n26548) );
  XNOR2X1 U49186 ( .A(n50799), .B(n42618), .Y(n26544) );
  XNOR2X1 U49187 ( .A(n50810), .B(net219310), .Y(n26341) );
  XNOR2X1 U49188 ( .A(n50177), .B(n42673), .Y(n26337) );
  XNOR2X1 U49189 ( .A(n50809), .B(n42615), .Y(n26333) );
  XNOR2X1 U49190 ( .A(n50803), .B(n36870), .Y(n26432) );
  XNOR2X1 U49191 ( .A(n50170), .B(n42673), .Y(n26428) );
  XNOR2X1 U49192 ( .A(n50802), .B(n42618), .Y(n26424) );
  XNOR2X1 U49193 ( .A(n50809), .B(net219330), .Y(n26311) );
  XNOR2X1 U49194 ( .A(n50176), .B(n42673), .Y(n26307) );
  XNOR2X1 U49195 ( .A(n50808), .B(n36868), .Y(n26303) );
  XNOR2X1 U49196 ( .A(n50804), .B(net219314), .Y(n26462) );
  XNOR2X1 U49197 ( .A(n50171), .B(n42673), .Y(n26458) );
  XNOR2X1 U49198 ( .A(n50803), .B(n42620), .Y(n26454) );
  XNOR2X1 U49199 ( .A(n50436), .B(n41379), .Y(n30129) );
  XNOR2X1 U49200 ( .A(n51067), .B(n42628), .Y(n30125) );
  XNOR2X1 U49201 ( .A(n50433), .B(n36903), .Y(n30189) );
  XNOR2X1 U49202 ( .A(n51064), .B(n42628), .Y(n30185) );
  XNOR2X1 U49203 ( .A(n50638), .B(n42504), .Y(n30116) );
  XNOR2X1 U49204 ( .A(n50432), .B(n36903), .Y(n30069) );
  XNOR2X1 U49205 ( .A(n51063), .B(n42629), .Y(n30065) );
  XNOR2X1 U49206 ( .A(n50635), .B(n42505), .Y(n30176) );
  XNOR2X1 U49207 ( .A(n50634), .B(n36731), .Y(n30056) );
  XNOR2X1 U49208 ( .A(n50435), .B(n36903), .Y(n30099) );
  XNOR2X1 U49209 ( .A(n51066), .B(n42624), .Y(n30095) );
  XNOR2X1 U49210 ( .A(n50631), .B(n36731), .Y(n29966) );
  XNOR2X1 U49211 ( .A(n50633), .B(n36730), .Y(n30026) );
  XNOR2X1 U49212 ( .A(n50630), .B(n42505), .Y(n29756) );
  XNOR2X1 U49213 ( .A(n50632), .B(n36730), .Y(n29996) );
  XNOR2X1 U49214 ( .A(n50627), .B(n42504), .Y(n29786) );
  XNOR2X1 U49215 ( .A(n50628), .B(n42505), .Y(n29816) );
  XNOR2X1 U49216 ( .A(n50424), .B(n36903), .Y(n29949) );
  XNOR2X1 U49217 ( .A(n51055), .B(n42632), .Y(n29945) );
  XNOR2X1 U49218 ( .A(n50422), .B(n36903), .Y(n29859) );
  XNOR2X1 U49219 ( .A(n51053), .B(n42625), .Y(n29855) );
  XNOR2X1 U49220 ( .A(n51044), .B(n41281), .Y(n26162) );
  XNOR2X1 U49221 ( .A(n50412), .B(n36903), .Y(n26158) );
  XNOR2X1 U49222 ( .A(n51043), .B(n42627), .Y(n26154) );
  XNOR2X1 U49223 ( .A(n50618), .B(n42505), .Y(n29605) );
  XNOR2X1 U49224 ( .A(n50637), .B(n42503), .Y(n30086) );
  XNOR2X1 U49225 ( .A(n51041), .B(n41282), .Y(n26072) );
  XNOR2X1 U49226 ( .A(n50409), .B(n41380), .Y(n26068) );
  XNOR2X1 U49227 ( .A(n51040), .B(n42628), .Y(n26064) );
  XNOR2X1 U49228 ( .A(n51038), .B(n41281), .Y(n26012) );
  XNOR2X1 U49229 ( .A(n50406), .B(n36903), .Y(n26008) );
  XNOR2X1 U49230 ( .A(n51037), .B(n42631), .Y(n26004) );
  XNOR2X1 U49231 ( .A(n50636), .B(n42502), .Y(n30146) );
  XNOR2X1 U49232 ( .A(n50614), .B(n42501), .Y(n26145) );
  XNOR2X1 U49233 ( .A(n50612), .B(n42501), .Y(n26085) );
  XNOR2X1 U49234 ( .A(n51040), .B(n41283), .Y(n25952) );
  XNOR2X1 U49235 ( .A(n50408), .B(n36903), .Y(n25948) );
  XNOR2X1 U49236 ( .A(n51039), .B(n34447), .Y(n25944) );
  XNOR2X1 U49237 ( .A(n50629), .B(n36737), .Y(n29726) );
  XNOR2X1 U49238 ( .A(n50611), .B(n42501), .Y(n26055) );
  XNOR2X1 U49239 ( .A(n50606), .B(n42501), .Y(n25815) );
  XNOR2X1 U49240 ( .A(n50608), .B(n42501), .Y(n25995) );
  XNOR2X1 U49241 ( .A(n50423), .B(n41379), .Y(n29889) );
  XNOR2X1 U49242 ( .A(n51054), .B(n42626), .Y(n29885) );
  XNOR2X1 U49243 ( .A(n51039), .B(n41281), .Y(n25982) );
  XNOR2X1 U49244 ( .A(n50407), .B(n36903), .Y(n25978) );
  XNOR2X1 U49245 ( .A(n51038), .B(n42633), .Y(n25974) );
  XNOR2X1 U49246 ( .A(n51037), .B(n41282), .Y(n26042) );
  XNOR2X1 U49247 ( .A(n50405), .B(n36903), .Y(n26038) );
  XNOR2X1 U49248 ( .A(n51036), .B(n42633), .Y(n26034) );
  XNOR2X1 U49249 ( .A(n50610), .B(n42501), .Y(n25935) );
  XNOR2X1 U49250 ( .A(n50624), .B(n42508), .Y(n29846) );
  XNOR2X1 U49251 ( .A(n51043), .B(n41283), .Y(n26132) );
  XNOR2X1 U49252 ( .A(n50411), .B(n36903), .Y(n26128) );
  XNOR2X1 U49253 ( .A(n51042), .B(n42629), .Y(n26124) );
  XNOR2X1 U49254 ( .A(n50609), .B(n42501), .Y(n25965) );
  XNOR2X1 U49255 ( .A(n50607), .B(n42501), .Y(n26025) );
  XNOR2X1 U49256 ( .A(n51042), .B(n41281), .Y(n26102) );
  XNOR2X1 U49257 ( .A(n50410), .B(n36903), .Y(n26098) );
  XNOR2X1 U49258 ( .A(n51041), .B(n42630), .Y(n26094) );
  XNOR2X1 U49259 ( .A(n50613), .B(n42501), .Y(n26115) );
  XNOR2X1 U49260 ( .A(n51025), .B(n41282), .Y(n26192) );
  XNOR2X1 U49261 ( .A(n50393), .B(n41319), .Y(n26188) );
  XNOR2X1 U49262 ( .A(n51024), .B(n42633), .Y(n26184) );
  XNOR2X1 U49263 ( .A(n50623), .B(n42505), .Y(n29906) );
  XNOR2X1 U49264 ( .A(n50625), .B(n42502), .Y(n29876) );
  XNOR2X1 U49265 ( .A(n50626), .B(n42501), .Y(n29936) );
  XNOR2X1 U49266 ( .A(n50605), .B(n42501), .Y(n25845) );
  XNOR2X1 U49267 ( .A(n50404), .B(n41380), .Y(n25828) );
  XNOR2X1 U49268 ( .A(n51035), .B(n42626), .Y(n25824) );
  XNOR2X1 U49269 ( .A(n51028), .B(n41281), .Y(n26282) );
  XNOR2X1 U49270 ( .A(n50396), .B(n36905), .Y(n26278) );
  XNOR2X1 U49271 ( .A(n51027), .B(n42631), .Y(n26274) );
  XNOR2X1 U49272 ( .A(n51033), .B(n41281), .Y(n25892) );
  XNOR2X1 U49273 ( .A(n50401), .B(n36903), .Y(n25888) );
  XNOR2X1 U49274 ( .A(n50621), .B(n42501), .Y(n29545) );
  XNOR2X1 U49275 ( .A(n50622), .B(n42503), .Y(n29575) );
  XNOR2X1 U49276 ( .A(n50594), .B(n42502), .Y(n26325) );
  XNOR2X1 U49277 ( .A(n50595), .B(n42501), .Y(n26175) );
  XNOR2X1 U49278 ( .A(n51034), .B(n41281), .Y(n25922) );
  XNOR2X1 U49279 ( .A(n50402), .B(n36903), .Y(n25918) );
  XNOR2X1 U49280 ( .A(n51033), .B(n42632), .Y(n25914) );
  XNOR2X1 U49281 ( .A(n51035), .B(n41281), .Y(n25862) );
  XNOR2X1 U49282 ( .A(n51034), .B(n42631), .Y(n25854) );
  XNOR2X1 U49283 ( .A(n51032), .B(n41283), .Y(n25742) );
  XNOR2X1 U49284 ( .A(n50616), .B(n42501), .Y(n29665) );
  XNOR2X1 U49285 ( .A(n50615), .B(n42506), .Y(n29695) );
  XNOR2X1 U49286 ( .A(n50617), .B(n42506), .Y(n29635) );
  XNOR2X1 U49287 ( .A(n50598), .B(n42503), .Y(n26265) );
  XNOR2X1 U49288 ( .A(n50604), .B(n42501), .Y(n25905) );
  XNOR2X1 U49289 ( .A(n50603), .B(n42501), .Y(n25875) );
  XNOR2X1 U49290 ( .A(n51029), .B(n41283), .Y(n25772) );
  XNOR2X1 U49291 ( .A(n50397), .B(n36903), .Y(n25768) );
  XNOR2X1 U49292 ( .A(n51028), .B(n42625), .Y(n25764) );
  XNOR2X1 U49293 ( .A(n50597), .B(n42502), .Y(n26235) );
  XNOR2X1 U49294 ( .A(n50596), .B(n42501), .Y(n26205) );
  XNOR2X1 U49295 ( .A(n51026), .B(n41283), .Y(n26222) );
  XNOR2X1 U49296 ( .A(n51025), .B(n42628), .Y(n26214) );
  XNOR2X1 U49297 ( .A(n51027), .B(n41283), .Y(n26252) );
  XNOR2X1 U49298 ( .A(n50395), .B(n34443), .Y(n26248) );
  XNOR2X1 U49299 ( .A(n51026), .B(n42625), .Y(n26244) );
  XNOR2X1 U49300 ( .A(n51019), .B(n41283), .Y(n26523) );
  XNOR2X1 U49301 ( .A(n50387), .B(n41319), .Y(n26519) );
  XNOR2X1 U49302 ( .A(n51018), .B(n42633), .Y(n26515) );
  XNOR2X1 U49303 ( .A(n51020), .B(n41283), .Y(n26493) );
  XNOR2X1 U49304 ( .A(n50388), .B(n41319), .Y(n26489) );
  XNOR2X1 U49305 ( .A(n51019), .B(n42632), .Y(n26485) );
  XNOR2X1 U49306 ( .A(n51030), .B(n41283), .Y(n25802) );
  XNOR2X1 U49307 ( .A(n50398), .B(n36903), .Y(n25798) );
  XNOR2X1 U49308 ( .A(n51029), .B(n42630), .Y(n25794) );
  XNOR2X1 U49309 ( .A(n51021), .B(n41282), .Y(n26372) );
  XNOR2X1 U49310 ( .A(n50389), .B(n36905), .Y(n26368) );
  XNOR2X1 U49311 ( .A(n51020), .B(n42631), .Y(n26364) );
  XNOR2X1 U49312 ( .A(n50390), .B(n36903), .Y(n26398) );
  XNOR2X1 U49313 ( .A(n51021), .B(n42624), .Y(n26394) );
  XNOR2X1 U49314 ( .A(n51022), .B(n41281), .Y(n26402) );
  XNOR2X1 U49315 ( .A(n50589), .B(n42508), .Y(n26506) );
  XNOR2X1 U49316 ( .A(n50590), .B(n42503), .Y(n26476) );
  XNOR2X1 U49317 ( .A(n50382), .B(n41319), .Y(n26549) );
  XNOR2X1 U49318 ( .A(n51013), .B(n42628), .Y(n26545) );
  XNOR2X1 U49319 ( .A(n50593), .B(n36731), .Y(n26295) );
  XNOR2X1 U49320 ( .A(n51024), .B(n41281), .Y(n26342) );
  XNOR2X1 U49321 ( .A(n50392), .B(n41319), .Y(n26338) );
  XNOR2X1 U49322 ( .A(n51023), .B(n42633), .Y(n26334) );
  XNOR2X1 U49323 ( .A(n51017), .B(n41282), .Y(n26433) );
  XNOR2X1 U49324 ( .A(n51016), .B(n42632), .Y(n26425) );
  XNOR2X1 U49325 ( .A(n50591), .B(n42503), .Y(n26355) );
  XNOR2X1 U49326 ( .A(n50592), .B(n42505), .Y(n26385) );
  XNOR2X1 U49327 ( .A(n51023), .B(n41283), .Y(n26312) );
  XNOR2X1 U49328 ( .A(n50391), .B(n41319), .Y(n26308) );
  XNOR2X1 U49329 ( .A(n51022), .B(n34447), .Y(n26304) );
  XNOR2X1 U49330 ( .A(n50584), .B(n36737), .Y(n26536) );
  XNOR2X1 U49331 ( .A(n50587), .B(n36730), .Y(n26416) );
  XNOR2X1 U49332 ( .A(n50588), .B(n42505), .Y(n26446) );
  XNOR2X1 U49333 ( .A(n51018), .B(n41283), .Y(n26463) );
  XNOR2X1 U49334 ( .A(n50386), .B(n41319), .Y(n26459) );
  XNOR2X1 U49335 ( .A(n51017), .B(n42629), .Y(n26455) );
  XOR2X1 U49336 ( .A(n42263), .B(n42654), .Y(n30071) );
  XOR2X1 U49337 ( .A(n42004), .B(n36711), .Y(n30067) );
  XOR2X1 U49338 ( .A(n42270), .B(n42647), .Y(n29801) );
  XOR2X1 U49339 ( .A(n42011), .B(n42602), .Y(n29797) );
  XOR2X1 U49340 ( .A(n42271), .B(n42667), .Y(n29951) );
  XOR2X1 U49341 ( .A(n42012), .B(n42602), .Y(n29947) );
  XOR2X1 U49342 ( .A(n42014), .B(n42602), .Y(n29857) );
  XOR2X1 U49343 ( .A(n42023), .B(n36891), .Y(n26164) );
  XOR2X1 U49344 ( .A(n42283), .B(n42654), .Y(n26160) );
  XOR2X1 U49345 ( .A(n42024), .B(n42606), .Y(n26156) );
  XOR2X1 U49346 ( .A(n42026), .B(n36899), .Y(n26074) );
  XOR2X1 U49347 ( .A(n42286), .B(n42654), .Y(n26070) );
  XOR2X1 U49348 ( .A(n42027), .B(n42606), .Y(n26066) );
  XOR2X1 U49349 ( .A(n42029), .B(n36892), .Y(n26014) );
  XOR2X1 U49350 ( .A(n42289), .B(n42654), .Y(n26010) );
  XOR2X1 U49351 ( .A(n42030), .B(n42606), .Y(n26006) );
  XOR2X1 U49352 ( .A(n42286), .B(n36885), .Y(n25958) );
  XOR2X1 U49353 ( .A(n42027), .B(n36893), .Y(n25954) );
  XOR2X1 U49354 ( .A(n42287), .B(n42648), .Y(n25950) );
  XOR2X1 U49355 ( .A(n42028), .B(n42606), .Y(n25946) );
  XOR2X1 U49356 ( .A(n42272), .B(n42665), .Y(n29891) );
  XOR2X1 U49357 ( .A(n42013), .B(n42602), .Y(n29887) );
  XOR2X1 U49358 ( .A(n42028), .B(n36894), .Y(n25984) );
  XOR2X1 U49359 ( .A(n42288), .B(n42654), .Y(n25980) );
  XOR2X1 U49360 ( .A(n42029), .B(n42606), .Y(n25976) );
  XOR2X1 U49361 ( .A(n42030), .B(n36895), .Y(n26044) );
  XOR2X1 U49362 ( .A(n42290), .B(n41286), .Y(n26040) );
  XOR2X1 U49363 ( .A(n42031), .B(n42606), .Y(n26036) );
  XOR2X1 U49364 ( .A(n42277), .B(n42657), .Y(n29530) );
  XOR2X1 U49365 ( .A(n42018), .B(n42602), .Y(n29526) );
  XOR2X1 U49366 ( .A(n42281), .B(n42651), .Y(n29680) );
  XOR2X1 U49367 ( .A(n42022), .B(n42602), .Y(n29676) );
  XOR2X1 U49368 ( .A(n42042), .B(n36901), .Y(n26194) );
  XOR2X1 U49369 ( .A(n42302), .B(n42663), .Y(n26190) );
  XOR2X1 U49370 ( .A(n42043), .B(n42606), .Y(n26186) );
  XOR2X1 U49371 ( .A(n42039), .B(n36899), .Y(n26284) );
  XOR2X1 U49372 ( .A(n42299), .B(n42665), .Y(n26280) );
  XOR2X1 U49373 ( .A(n42040), .B(n42606), .Y(n26276) );
  XOR2X1 U49374 ( .A(n42041), .B(n36901), .Y(n26224) );
  XOR2X1 U49375 ( .A(n42301), .B(n42664), .Y(n26220) );
  XOR2X1 U49376 ( .A(n42042), .B(n42606), .Y(n26216) );
  XOR2X1 U49377 ( .A(n42040), .B(n36897), .Y(n26254) );
  XOR2X1 U49378 ( .A(n42300), .B(n42648), .Y(n26250) );
  XOR2X1 U49379 ( .A(n42041), .B(n42606), .Y(n26246) );
  XOR2X1 U49380 ( .A(n42028), .B(n36754), .Y(n20916) );
  XOR2X1 U49381 ( .A(n42033), .B(n36761), .Y(n20853) );
  XOR2X1 U49382 ( .A(n42029), .B(n36759), .Y(n20885) );
  XOR2X1 U49383 ( .A(n42035), .B(n36753), .Y(n20873) );
  XOR2X1 U49384 ( .A(n42036), .B(n36753), .Y(n20863) );
  XOR2X1 U49385 ( .A(n42038), .B(n36757), .Y(n20810) );
  XOR2X1 U49386 ( .A(n42039), .B(n36755), .Y(n20831) );
  XOR2X1 U49387 ( .A(n42040), .B(n36756), .Y(n20821) );
  XOR2X1 U49388 ( .A(n41994), .B(n41317), .Y(n24455) );
  XOR2X1 U49389 ( .A(n41994), .B(n36754), .Y(n22061) );
  XOR2X1 U49390 ( .A(n41995), .B(n41310), .Y(n24445) );
  XOR2X1 U49391 ( .A(n41993), .B(n36760), .Y(n22071) );
  XOR2X1 U49392 ( .A(n41995), .B(n36753), .Y(n22051) );
  XOR2X1 U49393 ( .A(n41998), .B(n41318), .Y(n24405) );
  XOR2X1 U49394 ( .A(n41996), .B(n36761), .Y(n22041) );
  XOR2X1 U49395 ( .A(n41999), .B(n41314), .Y(n24395) );
  XOR2X1 U49396 ( .A(n42002), .B(n41311), .Y(n24475) );
  XOR2X1 U49397 ( .A(n42003), .B(n41309), .Y(n24465) );
  XOR2X1 U49398 ( .A(n42003), .B(n36755), .Y(n21991) );
  XOR2X1 U49399 ( .A(n42004), .B(n36753), .Y(n21981) );
  XOR2X1 U49400 ( .A(n42006), .B(n36755), .Y(n21951) );
  XOR2X1 U49401 ( .A(n42009), .B(n41314), .Y(n24273) );
  XOR2X1 U49402 ( .A(n41997), .B(n41318), .Y(n24425) );
  XOR2X1 U49403 ( .A(n42007), .B(n36760), .Y(n21971) );
  XOR2X1 U49404 ( .A(n42010), .B(n41309), .Y(n24263) );
  XOR2X1 U49405 ( .A(n41996), .B(n41318), .Y(n24435) );
  XOR2X1 U49406 ( .A(n42008), .B(n36761), .Y(n21961) );
  XOR2X1 U49407 ( .A(n42011), .B(n41317), .Y(n24253) );
  XOR2X1 U49408 ( .A(n42013), .B(n41316), .Y(n24293) );
  XOR2X1 U49409 ( .A(n42001), .B(n41313), .Y(n24485) );
  XOR2X1 U49410 ( .A(n42007), .B(n41311), .Y(n24353) );
  XOR2X1 U49411 ( .A(n42008), .B(n41310), .Y(n24343) );
  XOR2X1 U49412 ( .A(n42015), .B(n41311), .Y(n24243) );
  XOR2X1 U49413 ( .A(n42014), .B(n36754), .Y(n21859) );
  XOR2X1 U49414 ( .A(n42005), .B(n41313), .Y(n24373) );
  XOR2X1 U49415 ( .A(n42006), .B(n41316), .Y(n24363) );
  XOR2X1 U49416 ( .A(n41997), .B(n36757), .Y(n22021) );
  XOR2X1 U49417 ( .A(n41998), .B(n36760), .Y(n22031) );
  XOR2X1 U49418 ( .A(n42002), .B(n36754), .Y(n22001) );
  XOR2X1 U49419 ( .A(n42001), .B(n36756), .Y(n22011) );
  XOR2X1 U49420 ( .A(n42012), .B(n41317), .Y(n24283) );
  XOR2X1 U49421 ( .A(n42018), .B(n36761), .Y(n21910) );
  XOR2X1 U49422 ( .A(n42021), .B(n41310), .Y(n24333) );
  XOR2X1 U49423 ( .A(n42017), .B(n36757), .Y(n21829) );
  XOR2X1 U49424 ( .A(n42019), .B(n36754), .Y(n21931) );
  XOR2X1 U49425 ( .A(n42022), .B(n41316), .Y(n24323) );
  XOR2X1 U49426 ( .A(n42020), .B(n36756), .Y(n21921) );
  XOR2X1 U49427 ( .A(n42022), .B(n36754), .Y(n21890) );
  XOR2X1 U49428 ( .A(n42023), .B(n41309), .Y(n24303) );
  XOR2X1 U49429 ( .A(n42024), .B(n41317), .Y(n24313) );
  XOR2X1 U49430 ( .A(n42013), .B(n36760), .Y(n21819) );
  XOR2X1 U49431 ( .A(n42016), .B(n36754), .Y(n21839) );
  XOR2X1 U49432 ( .A(n42015), .B(n36755), .Y(n21849) );
  XOR2X1 U49433 ( .A(n42025), .B(n41311), .Y(n24607) );
  XOR2X1 U49434 ( .A(n42026), .B(n41312), .Y(n24617) );
  XOR2X1 U49435 ( .A(n42021), .B(n36756), .Y(n21900) );
  XOR2X1 U49436 ( .A(n42023), .B(n36756), .Y(n21870) );
  XOR2X1 U49437 ( .A(n42028), .B(n41318), .Y(n24587) );
  XOR2X1 U49438 ( .A(n42027), .B(n41317), .Y(n24597) );
  XOR2X1 U49439 ( .A(n42024), .B(n36755), .Y(n21880) );
  XOR2X1 U49440 ( .A(n42029), .B(n41309), .Y(n24567) );
  XOR2X1 U49441 ( .A(n42032), .B(n41316), .Y(n24577) );
  XOR2X1 U49442 ( .A(n42036), .B(n41312), .Y(n24627) );
  XOR2X1 U49443 ( .A(n42030), .B(n41311), .Y(n24545) );
  XOR2X1 U49444 ( .A(n42031), .B(n41313), .Y(n24556) );
  XOR2X1 U49445 ( .A(n42037), .B(n41313), .Y(n24525) );
  XOR2X1 U49446 ( .A(n42038), .B(n41310), .Y(n24535) );
  XOR2X1 U49447 ( .A(n42000), .B(n41318), .Y(n24385) );
  XOR2X1 U49448 ( .A(n42004), .B(n41318), .Y(n24495) );
  XOR2X1 U49449 ( .A(n42040), .B(n41316), .Y(n24505) );
  XOR2X1 U49450 ( .A(n42039), .B(n41309), .Y(n24515) );
  XOR2X1 U49451 ( .A(n42005), .B(n36756), .Y(n21941) );
  XOR2X1 U49452 ( .A(n42001), .B(n42515), .Y(n30117) );
  XOR2X1 U49453 ( .A(n42004), .B(n42515), .Y(n30177) );
  XOR2X1 U49454 ( .A(n42005), .B(n42522), .Y(n30057) );
  XOR2X1 U49455 ( .A(n42007), .B(n42515), .Y(n29997) );
  XOR2X1 U49456 ( .A(n42012), .B(n42518), .Y(n29787) );
  XOR2X1 U49457 ( .A(n42011), .B(n42518), .Y(n29817) );
  XOR2X1 U49458 ( .A(n42021), .B(n42518), .Y(n29606) );
  XOR2X1 U49459 ( .A(n42002), .B(n42515), .Y(n30087) );
  XOR2X1 U49460 ( .A(n42003), .B(n42529), .Y(n30147) );
  XOR2X1 U49461 ( .A(n42025), .B(n42522), .Y(n26146) );
  XOR2X1 U49462 ( .A(n42027), .B(n42512), .Y(n26086) );
  XOR2X1 U49463 ( .A(n42010), .B(n42518), .Y(n29727) );
  XOR2X1 U49464 ( .A(n42028), .B(n42522), .Y(n26056) );
  XOR2X1 U49465 ( .A(n42015), .B(n42518), .Y(n29847) );
  XOR2X1 U49466 ( .A(n42032), .B(n42521), .Y(n26026) );
  XOR2X1 U49467 ( .A(n42026), .B(n42528), .Y(n26116) );
  XOR2X1 U49468 ( .A(n42016), .B(n42515), .Y(n29907) );
  XOR2X1 U49469 ( .A(n42014), .B(n42518), .Y(n29877) );
  XOR2X1 U49470 ( .A(n42013), .B(n42515), .Y(n29937) );
  XOR2X1 U49471 ( .A(n42018), .B(n42518), .Y(n29546) );
  XOR2X1 U49472 ( .A(n42017), .B(n42518), .Y(n29576) );
  XOR2X1 U49473 ( .A(n42045), .B(n42521), .Y(n26326) );
  XOR2X1 U49474 ( .A(n42044), .B(n42528), .Y(n26176) );
  XOR2X1 U49475 ( .A(n42023), .B(n42518), .Y(n29666) );
  XOR2X1 U49476 ( .A(n42024), .B(n42518), .Y(n29696) );
  XOR2X1 U49477 ( .A(n42022), .B(n42518), .Y(n29636) );
  XOR2X1 U49478 ( .A(n42041), .B(n42529), .Y(n26266) );
  XOR2X1 U49479 ( .A(n42042), .B(n42519), .Y(n26236) );
  XOR2X1 U49480 ( .A(n42043), .B(n42528), .Y(n26206) );
  XOR2X1 U49481 ( .A(n42046), .B(n42518), .Y(n26296) );
  XOR2X1 U49482 ( .A(n42048), .B(n42512), .Y(n26356) );
  NAND4X1 U49483 ( .A(n10470), .B(n10469), .C(n10471), .D(n29719), .Y(n9950)
         );
  NOR2X1 U49484 ( .A(net171178), .B(n10611), .Y(n29719) );
  NAND4X1 U49485 ( .A(net260299), .B(n11915), .C(net260295), .D(n29478), .Y(
        n9951) );
  NOR2X1 U49486 ( .A(n_cell_301249_net269596), .B(n10463), .Y(n29478) );
  OR2X2 U49487 ( .A(n9689), .B(out_valid), .Y(n19180) );
  XNOR2X1 U49488 ( .A(n50429), .B(n36768), .Y(n21973) );
  XNOR2X1 U49489 ( .A(n50428), .B(n36773), .Y(n21963) );
  XNOR2X1 U49490 ( .A(n50422), .B(n36774), .Y(n21861) );
  XNOR2X1 U49491 ( .A(n50417), .B(n36772), .Y(n21933) );
  XNOR2X1 U49492 ( .A(n50416), .B(n36772), .Y(n21923) );
  XNOR2X1 U49493 ( .A(n50420), .B(n36771), .Y(n21841) );
  XNOR2X1 U49494 ( .A(n50415), .B(n36765), .Y(n21902) );
  XNOR2X1 U49495 ( .A(n51287), .B(n41305), .Y(n24457) );
  XNOR2X1 U49496 ( .A(n51287), .B(n36746), .Y(n22063) );
  XNOR2X1 U49497 ( .A(n51286), .B(n41301), .Y(n24447) );
  XNOR2X1 U49498 ( .A(n51286), .B(n36749), .Y(n22053) );
  XNOR2X1 U49499 ( .A(n51283), .B(n41300), .Y(n24407) );
  XNOR2X1 U49500 ( .A(n51285), .B(n36749), .Y(n22043) );
  XNOR2X1 U49501 ( .A(n51282), .B(n41305), .Y(n24397) );
  XNOR2X1 U49502 ( .A(n51279), .B(n41303), .Y(n24477) );
  XNOR2X1 U49503 ( .A(n51278), .B(n41300), .Y(n24467) );
  XNOR2X1 U49504 ( .A(n51278), .B(n36748), .Y(n21993) );
  XNOR2X1 U49505 ( .A(n51277), .B(n36750), .Y(n21983) );
  XNOR2X1 U49506 ( .A(n51275), .B(n36744), .Y(n21953) );
  XNOR2X1 U49507 ( .A(n51284), .B(n41304), .Y(n24427) );
  XNOR2X1 U49508 ( .A(n51271), .B(n41299), .Y(n24265) );
  XNOR2X1 U49509 ( .A(n51285), .B(n41302), .Y(n24437) );
  XNOR2X1 U49510 ( .A(n51271), .B(n36744), .Y(n21801) );
  XNOR2X1 U49511 ( .A(n51270), .B(n41304), .Y(n24255) );
  XNOR2X1 U49512 ( .A(n51268), .B(n41300), .Y(n24295) );
  XNOR2X1 U49513 ( .A(n51280), .B(n41302), .Y(n24487) );
  XNOR2X1 U49514 ( .A(n51266), .B(n41300), .Y(n24245) );
  XNOR2X1 U49515 ( .A(n51276), .B(n41303), .Y(n24375) );
  XNOR2X1 U49516 ( .A(n51275), .B(n41300), .Y(n24365) );
  XNOR2X1 U49517 ( .A(n51284), .B(n36741), .Y(n22023) );
  XNOR2X1 U49518 ( .A(n51283), .B(n36748), .Y(n22033) );
  XNOR2X1 U49519 ( .A(n51279), .B(n36748), .Y(n22003) );
  XNOR2X1 U49520 ( .A(n51280), .B(n36741), .Y(n22013) );
  XNOR2X1 U49521 ( .A(n51269), .B(n41299), .Y(n24285) );
  XNOR2X1 U49522 ( .A(n51268), .B(n36743), .Y(n21821) );
  XNOR2X1 U49523 ( .A(n51255), .B(n41304), .Y(n24619) );
  XNOR2X1 U49524 ( .A(n51253), .B(n41300), .Y(n24589) );
  XNOR2X1 U49525 ( .A(n51254), .B(n41304), .Y(n24599) );
  XNOR2X1 U49526 ( .A(n51252), .B(n41304), .Y(n24569) );
  XNOR2X1 U49527 ( .A(n51255), .B(n36746), .Y(n20908) );
  XNOR2X1 U49528 ( .A(n51249), .B(n41305), .Y(n24579) );
  XNOR2X1 U49529 ( .A(n51253), .B(n36746), .Y(n20918) );
  XNOR2X1 U49530 ( .A(n51251), .B(n41305), .Y(n24548) );
  XNOR2X1 U49531 ( .A(n51251), .B(n36744), .Y(n20897) );
  XNOR2X1 U49532 ( .A(n51250), .B(n41301), .Y(n24559) );
  XNOR2X1 U49533 ( .A(n51244), .B(n41305), .Y(n24527) );
  XNOR2X1 U49534 ( .A(n51248), .B(n36748), .Y(n20855) );
  XNOR2X1 U49535 ( .A(n51247), .B(n36743), .Y(n20845) );
  XNOR2X1 U49536 ( .A(n51252), .B(n36746), .Y(n20887) );
  XNOR2X1 U49537 ( .A(n51281), .B(n41303), .Y(n24387) );
  XNOR2X1 U49538 ( .A(n51277), .B(n41305), .Y(n24497) );
  XNOR2X1 U49539 ( .A(n51246), .B(n36744), .Y(n20876) );
  XNOR2X1 U49540 ( .A(n51245), .B(n36748), .Y(n20865) );
  XNOR2X1 U49541 ( .A(n51243), .B(n36742), .Y(n20813) );
  XNOR2X1 U49542 ( .A(n51231), .B(n36744), .Y(n20466) );
  XNOR2X1 U49543 ( .A(n51244), .B(n36749), .Y(n20802) );
  XNOR2X1 U49544 ( .A(n51276), .B(n36746), .Y(n21943) );
  XNOR2X1 U49545 ( .A(n51228), .B(n36741), .Y(n20496) );
  XNOR2X1 U49546 ( .A(n51227), .B(n36742), .Y(n20506) );
  NOR2X1 U49547 ( .A(net171108), .B(net171111), .Y(n31886) );
  XNOR2X1 U49548 ( .A(n50443), .B(n42581), .Y(n30300) );
  XNOR2X1 U49549 ( .A(n50441), .B(n42578), .Y(n30210) );
  XNOR2X1 U49550 ( .A(n50435), .B(n42577), .Y(n30119) );
  XNOR2X1 U49551 ( .A(n50432), .B(n42578), .Y(n30179) );
  XNOR2X1 U49552 ( .A(n50431), .B(n42578), .Y(n30059) );
  XNOR2X1 U49553 ( .A(n50428), .B(n42577), .Y(n29969) );
  XNOR2X1 U49554 ( .A(n50430), .B(n42581), .Y(n30029) );
  XNOR2X1 U49555 ( .A(n50427), .B(n42576), .Y(n29759) );
  XNOR2X1 U49556 ( .A(n50429), .B(n42577), .Y(n29999) );
  XNOR2X1 U49557 ( .A(n50424), .B(n34451), .Y(n29789) );
  XNOR2X1 U49558 ( .A(n50425), .B(n42579), .Y(n29819) );
  XNOR2X1 U49559 ( .A(n50417), .B(n42576), .Y(n29518) );
  XNOR2X1 U49560 ( .A(n50416), .B(n42579), .Y(n29488) );
  XNOR2X1 U49561 ( .A(n50415), .B(n42579), .Y(n29608) );
  XNOR2X1 U49562 ( .A(n50434), .B(n42579), .Y(n30089) );
  XNOR2X1 U49563 ( .A(n50433), .B(n42577), .Y(n30149) );
  XNOR2X1 U49564 ( .A(n50411), .B(n42575), .Y(n26148) );
  XNOR2X1 U49565 ( .A(n50409), .B(n42575), .Y(n26088) );
  XNOR2X1 U49566 ( .A(n50426), .B(n42576), .Y(n29729) );
  XNOR2X1 U49567 ( .A(n50408), .B(n42575), .Y(n26058) );
  XNOR2X1 U49568 ( .A(n50403), .B(n42576), .Y(n25818) );
  XNOR2X1 U49569 ( .A(n50405), .B(n42575), .Y(n25998) );
  XNOR2X1 U49570 ( .A(n50407), .B(n42576), .Y(n25938) );
  XNOR2X1 U49571 ( .A(n50421), .B(n42576), .Y(n29849) );
  XNOR2X1 U49572 ( .A(n50437), .B(n42583), .Y(n30330) );
  XNOR2X1 U49573 ( .A(n50438), .B(n42584), .Y(n30420) );
  XNOR2X1 U49574 ( .A(n50436), .B(n42580), .Y(n30360) );
  XNOR2X1 U49575 ( .A(n50406), .B(n42575), .Y(n25968) );
  XNOR2X1 U49576 ( .A(n50404), .B(n42576), .Y(n26028) );
  XNOR2X1 U49577 ( .A(n50410), .B(n42579), .Y(n26118) );
  XNOR2X1 U49578 ( .A(n50420), .B(n42579), .Y(n29909) );
  XNOR2X1 U49579 ( .A(n50422), .B(n42577), .Y(n29879) );
  XNOR2X1 U49580 ( .A(n50423), .B(n42577), .Y(n29939) );
  XNOR2X1 U49581 ( .A(n50402), .B(n42580), .Y(n25848) );
  XNOR2X1 U49582 ( .A(n50418), .B(n42576), .Y(n29548) );
  XNOR2X1 U49583 ( .A(n50419), .B(n42576), .Y(n29578) );
  XNOR2X1 U49584 ( .A(n50391), .B(n42577), .Y(n26328) );
  XNOR2X1 U49585 ( .A(n50392), .B(n34451), .Y(n26178) );
  XNOR2X1 U49586 ( .A(n50413), .B(n42576), .Y(n29668) );
  XNOR2X1 U49587 ( .A(n50412), .B(n42576), .Y(n29698) );
  XNOR2X1 U49588 ( .A(n50414), .B(n42576), .Y(n29638) );
  XNOR2X1 U49589 ( .A(n50395), .B(n42579), .Y(n26268) );
  XNOR2X1 U49590 ( .A(n50401), .B(n42580), .Y(n25908) );
  XNOR2X1 U49591 ( .A(n50400), .B(n42579), .Y(n25878) );
  XNOR2X1 U49592 ( .A(n50394), .B(n34451), .Y(n26238) );
  XNOR2X1 U49593 ( .A(n50393), .B(n34451), .Y(n26208) );
  XNOR2X1 U49594 ( .A(n50397), .B(n42580), .Y(n25788) );
  XNOR2X1 U49595 ( .A(n50386), .B(n42579), .Y(n26509) );
  XNOR2X1 U49596 ( .A(n50387), .B(n42576), .Y(n26479) );
  XNOR2X1 U49597 ( .A(n50390), .B(n42579), .Y(n26298) );
  XNOR2X1 U49598 ( .A(n50388), .B(n42576), .Y(n26358) );
  XNOR2X1 U49599 ( .A(n50389), .B(n42580), .Y(n26388) );
  XNOR2X1 U49600 ( .A(n50381), .B(n34451), .Y(n26539) );
  XNOR2X1 U49601 ( .A(n50384), .B(n42577), .Y(n26419) );
  XNOR2X1 U49602 ( .A(n50385), .B(n34451), .Y(n26449) );
  XOR2X1 U49603 ( .A(n42287), .B(n42486), .Y(n20917) );
  XOR2X1 U49604 ( .A(n42289), .B(n42479), .Y(n20896) );
  XOR2X1 U49605 ( .A(n42292), .B(n42483), .Y(n20854) );
  XOR2X1 U49606 ( .A(n42293), .B(n42479), .Y(n20843) );
  XOR2X1 U49607 ( .A(n42288), .B(n42487), .Y(n20886) );
  XOR2X1 U49608 ( .A(n42294), .B(n42486), .Y(n20874) );
  XOR2X1 U49609 ( .A(n42295), .B(n42479), .Y(n20864) );
  XOR2X1 U49610 ( .A(n42297), .B(n42479), .Y(n20811) );
  XOR2X1 U49611 ( .A(n42298), .B(n42479), .Y(n20832) );
  XOR2X1 U49612 ( .A(n42299), .B(n42479), .Y(n20822) );
  XOR2X1 U49613 ( .A(n42253), .B(n36807), .Y(n24456) );
  XOR2X1 U49614 ( .A(n42253), .B(n42492), .Y(n22062) );
  XOR2X1 U49615 ( .A(n42254), .B(n36811), .Y(n24446) );
  XOR2X1 U49616 ( .A(n42252), .B(n42488), .Y(n22072) );
  XOR2X1 U49617 ( .A(n42254), .B(n42486), .Y(n22052) );
  XOR2X1 U49618 ( .A(n42257), .B(n36814), .Y(n24406) );
  XOR2X1 U49619 ( .A(n42255), .B(n42486), .Y(n22042) );
  XOR2X1 U49620 ( .A(n42258), .B(n36814), .Y(n24396) );
  XOR2X1 U49621 ( .A(n42261), .B(n36809), .Y(n24476) );
  XOR2X1 U49622 ( .A(n42262), .B(n36807), .Y(n24466) );
  XOR2X1 U49623 ( .A(n42262), .B(n42479), .Y(n21992) );
  XOR2X1 U49624 ( .A(n42263), .B(n42491), .Y(n21982) );
  XOR2X1 U49625 ( .A(n42265), .B(n42486), .Y(n21952) );
  XOR2X1 U49626 ( .A(n42268), .B(n36816), .Y(n24274) );
  XOR2X1 U49627 ( .A(n42256), .B(n36817), .Y(n24426) );
  XOR2X1 U49628 ( .A(n42266), .B(n42486), .Y(n21972) );
  XOR2X1 U49629 ( .A(n42269), .B(n36810), .Y(n24264) );
  XOR2X1 U49630 ( .A(n42255), .B(n36810), .Y(n24436) );
  XOR2X1 U49631 ( .A(n42267), .B(n42478), .Y(n21962) );
  XOR2X1 U49632 ( .A(n42270), .B(n36816), .Y(n24254) );
  XOR2X1 U49633 ( .A(n42272), .B(n36813), .Y(n24294) );
  XOR2X1 U49634 ( .A(n42260), .B(n36813), .Y(n24486) );
  XOR2X1 U49635 ( .A(n42266), .B(n36816), .Y(n24354) );
  XOR2X1 U49636 ( .A(n42267), .B(n36816), .Y(n24344) );
  XOR2X1 U49637 ( .A(n42274), .B(n36817), .Y(n24244) );
  XOR2X1 U49638 ( .A(n42273), .B(n42488), .Y(n21860) );
  XOR2X1 U49639 ( .A(n42264), .B(n36807), .Y(n24374) );
  XOR2X1 U49640 ( .A(n42265), .B(n36807), .Y(n24364) );
  XOR2X1 U49641 ( .A(n42256), .B(n42486), .Y(n22022) );
  XOR2X1 U49642 ( .A(n42257), .B(n42479), .Y(n22032) );
  XOR2X1 U49643 ( .A(n42261), .B(n42479), .Y(n22002) );
  XOR2X1 U49644 ( .A(n42260), .B(n42492), .Y(n22012) );
  XOR2X1 U49645 ( .A(n42271), .B(n36815), .Y(n24284) );
  XOR2X1 U49646 ( .A(n42277), .B(n42488), .Y(n21911) );
  XOR2X1 U49647 ( .A(n42280), .B(n36807), .Y(n24334) );
  XOR2X1 U49648 ( .A(n42276), .B(n42488), .Y(n21830) );
  XOR2X1 U49649 ( .A(n42278), .B(n42488), .Y(n21932) );
  XOR2X1 U49650 ( .A(n42281), .B(n36808), .Y(n24324) );
  XOR2X1 U49651 ( .A(n42279), .B(n42488), .Y(n21922) );
  XOR2X1 U49652 ( .A(n42281), .B(n42488), .Y(n21891) );
  XOR2X1 U49653 ( .A(n42282), .B(n36815), .Y(n24304) );
  XOR2X1 U49654 ( .A(n42283), .B(n36815), .Y(n24314) );
  XOR2X1 U49655 ( .A(n42272), .B(n42488), .Y(n21820) );
  XOR2X1 U49656 ( .A(n42275), .B(n42488), .Y(n21840) );
  XOR2X1 U49657 ( .A(n42274), .B(n42488), .Y(n21850) );
  XOR2X1 U49658 ( .A(n42284), .B(n36814), .Y(n24608) );
  XOR2X1 U49659 ( .A(n42285), .B(n36815), .Y(n24618) );
  XOR2X1 U49660 ( .A(n42280), .B(n42488), .Y(n21901) );
  XOR2X1 U49661 ( .A(n42282), .B(n42488), .Y(n21871) );
  XOR2X1 U49662 ( .A(n42287), .B(n36815), .Y(n24588) );
  XOR2X1 U49663 ( .A(n42286), .B(n36810), .Y(n24598) );
  XOR2X1 U49664 ( .A(n42283), .B(n42488), .Y(n21881) );
  XOR2X1 U49665 ( .A(n42288), .B(n36811), .Y(n24568) );
  XOR2X1 U49666 ( .A(n42291), .B(n36816), .Y(n24578) );
  XOR2X1 U49667 ( .A(n42295), .B(n36811), .Y(n24628) );
  XOR2X1 U49668 ( .A(n42289), .B(n36815), .Y(n24546) );
  XOR2X1 U49669 ( .A(n42290), .B(n36807), .Y(n24557) );
  XOR2X1 U49670 ( .A(n42296), .B(n36808), .Y(n24526) );
  XOR2X1 U49671 ( .A(n42297), .B(n36817), .Y(n24536) );
  XOR2X1 U49672 ( .A(n42259), .B(n36816), .Y(n24386) );
  XOR2X1 U49673 ( .A(n42263), .B(n36817), .Y(n24496) );
  XOR2X1 U49674 ( .A(n42299), .B(n36817), .Y(n24506) );
  XOR2X1 U49675 ( .A(n42298), .B(n36815), .Y(n24516) );
  XOR2X1 U49676 ( .A(n42264), .B(n42488), .Y(n21942) );
  XOR2X1 U49677 ( .A(n42260), .B(n36801), .Y(n30118) );
  XOR2X1 U49678 ( .A(n42263), .B(n41321), .Y(n30178) );
  XOR2X1 U49679 ( .A(n42264), .B(n41323), .Y(n30058) );
  XOR2X1 U49680 ( .A(n42265), .B(n36801), .Y(n30028) );
  XOR2X1 U49681 ( .A(n42268), .B(n41323), .Y(n29758) );
  XOR2X1 U49682 ( .A(n42266), .B(n36877), .Y(n29998) );
  XOR2X1 U49683 ( .A(n42271), .B(n41321), .Y(n29788) );
  XOR2X1 U49684 ( .A(n42270), .B(n36873), .Y(n29818) );
  XOR2X1 U49685 ( .A(n42280), .B(n41322), .Y(n29607) );
  XOR2X1 U49686 ( .A(n42261), .B(n41323), .Y(n30088) );
  XOR2X1 U49687 ( .A(n42262), .B(n36801), .Y(n30148) );
  XOR2X1 U49688 ( .A(n42284), .B(n41321), .Y(n26147) );
  XOR2X1 U49689 ( .A(n42286), .B(n41322), .Y(n26087) );
  XOR2X1 U49690 ( .A(n42269), .B(n41323), .Y(n29728) );
  XOR2X1 U49691 ( .A(n42287), .B(n36877), .Y(n26057) );
  XOR2X1 U49692 ( .A(n42274), .B(n41322), .Y(n29848) );
  XOR2X1 U49693 ( .A(n42291), .B(n41323), .Y(n26027) );
  XOR2X1 U49694 ( .A(n42285), .B(n36877), .Y(n26117) );
  XOR2X1 U49695 ( .A(n42275), .B(n36873), .Y(n29908) );
  XOR2X1 U49696 ( .A(n42273), .B(n36877), .Y(n29878) );
  XOR2X1 U49697 ( .A(n42272), .B(n36801), .Y(n29938) );
  XOR2X1 U49698 ( .A(n42277), .B(n36877), .Y(n29547) );
  XOR2X1 U49699 ( .A(n42276), .B(n41323), .Y(n29577) );
  XOR2X1 U49700 ( .A(n42304), .B(n36877), .Y(n26327) );
  XOR2X1 U49701 ( .A(n42303), .B(n36801), .Y(n26177) );
  XOR2X1 U49702 ( .A(n42282), .B(n36801), .Y(n29667) );
  XOR2X1 U49703 ( .A(n42283), .B(n41321), .Y(n29697) );
  XOR2X1 U49704 ( .A(n42281), .B(n36877), .Y(n29637) );
  XOR2X1 U49705 ( .A(n42300), .B(n41322), .Y(n26267) );
  XOR2X1 U49706 ( .A(n42301), .B(n41323), .Y(n26237) );
  XOR2X1 U49707 ( .A(n42302), .B(n36801), .Y(n26207) );
  XOR2X1 U49708 ( .A(n42305), .B(n41321), .Y(n26297) );
  XOR2X1 U49709 ( .A(n42307), .B(n36801), .Y(n26357) );
  XOR2X1 U49710 ( .A(n42030), .B(n36757), .Y(n20895) );
  XNOR2X1 U49711 ( .A(n50609), .B(n42463), .Y(n20894) );
  XNOR2X1 U49712 ( .A(n51037), .B(n36716), .Y(n20893) );
  NOR4X1 U49713 ( .A(n20842), .B(n20841), .C(n20840), .D(n20839), .Y(net211600) );
  XOR2X1 U49714 ( .A(n42034), .B(n36755), .Y(n20842) );
  XNOR2X1 U49715 ( .A(n50605), .B(n42464), .Y(n20841) );
  XNOR2X1 U49716 ( .A(n51033), .B(n36718), .Y(n20840) );
  NOR4X1 U49717 ( .A(n25955), .B(n25956), .C(n25957), .D(n25958), .Y(n44390)
         );
  XNOR2X1 U49718 ( .A(n50194), .B(n42705), .Y(n25955) );
  XNOR2X1 U49719 ( .A(n50409), .B(n42719), .Y(n25956) );
  NOR4X1 U49720 ( .A(n25835), .B(n25836), .C(n25837), .D(n25838), .Y(net215014) );
  NOR4X1 U49721 ( .A(n25895), .B(n25896), .C(n25897), .D(n25898), .Y(n44406)
         );
  XNOR2X1 U49722 ( .A(n50187), .B(n42705), .Y(n25895) );
  XNOR2X1 U49723 ( .A(n50402), .B(n42723), .Y(n25896) );
  NOR4X1 U49724 ( .A(n25715), .B(n25716), .C(n25717), .D(n25718), .Y(net214960) );
  NOR4X1 U49725 ( .A(n25745), .B(n25746), .C(n25747), .D(n25748), .Y(n44417)
         );
  XNOR2X1 U49726 ( .A(n50184), .B(n42711), .Y(n25805) );
  XNOR2X1 U49727 ( .A(n50399), .B(n42720), .Y(n25806) );
  NOR4X1 U49728 ( .A(n25775), .B(n25776), .C(n25777), .D(n25778), .Y(n44412)
         );
  XNOR2X1 U49729 ( .A(n50183), .B(n41642), .Y(n25775) );
  XNOR2X1 U49730 ( .A(n50398), .B(n34435), .Y(n25776) );
  NOR4X1 U49731 ( .A(n26556), .B(n26557), .C(n26558), .D(n26559), .Y(net215194) );
  XNOR2X1 U49732 ( .A(n50168), .B(n42706), .Y(n26556) );
  XNOR2X1 U49733 ( .A(n50383), .B(n41287), .Y(n26557) );
  NOR4X1 U49734 ( .A(n26436), .B(n26437), .C(n26438), .D(n26439), .Y(net214746) );
  XNOR2X1 U49735 ( .A(n50171), .B(n42706), .Y(n26436) );
  XNOR2X1 U49736 ( .A(n50386), .B(n34435), .Y(n26437) );
  XNOR2X1 U49737 ( .A(n51231), .B(n41385), .Y(n26438) );
  NOR4X1 U49738 ( .A(n26616), .B(n26617), .C(n26618), .D(n26619), .Y(net215158) );
  NOR4X1 U49739 ( .A(n26586), .B(n26587), .C(n26588), .D(n26589), .Y(net215203) );
  NOR4X1 U49740 ( .A(n26646), .B(n26647), .C(n26648), .D(n26649), .Y(net215167) );
  NOR4X1 U49741 ( .A(n24702), .B(n24703), .C(n24704), .D(n24705), .Y(net214738) );
  NAND4X1 U49742 ( .A(n11893), .B(n11894), .C(n11895), .D(n11896), .Y(n10136)
         );
  OAI21XL U49743 ( .A0(net171349), .A1(n9715), .B0(n9734), .Y(n9733) );
  NOR3BXL U49744 ( .AN(net210435), .B(net210444), .C(net210445), .Y(n27614) );
  NAND3X1 U49745 ( .A(n11901), .B(n11902), .C(n11897), .Y(n10137) );
  NAND2BX1 U49746 ( .AN(net209395), .B(n12811), .Y(net209977) );
  AND4X1 U49747 ( .A(n_cell_303546_net275987), .B(n_cell_303546_net275967),
        .C(n10480), .D(n30200), .Y(n10140) );
  NOR2X1 U49748 ( .A(net151542), .B(n10610), .Y(n30200) );
  OR2XL U49749 ( .A(n19180), .B(n41796), .Y(net151225) );
  OR4X1 U49750 ( .A(n19506), .B(n19507), .C(n19508), .D(n19509), .Y(n36633) );
  OAI222XL U49751 ( .A0(n49543), .A1(n41797), .B0(n49527), .B1(n42729), .C0(
        n49535), .C1(n42728), .Y(n19508) );
  OAI22XL U49752 ( .A0(n42637), .A1(n42452), .B0(n42698), .B1(n19492), .Y(
        n19509) );
  OAI222XL U49753 ( .A0(n49551), .A1(n19493), .B0(n36831), .B1(n43040), .C0(
        n36744), .C1(n43044), .Y(n19506) );
  OR4X1 U49754 ( .A(n19502), .B(n19503), .C(n19504), .D(n19505), .Y(n36632) );
  OAI222XL U49755 ( .A0(n49544), .A1(n41797), .B0(n49528), .B1(n42729), .C0(
        n49536), .C1(n42728), .Y(n19504) );
  OAI22XL U49756 ( .A0(n34447), .A1(n42452), .B0(n41283), .B1(n19492), .Y(
        n19505) );
  OAI222XL U49757 ( .A0(n49552), .A1(n19493), .B0(n42554), .B1(n43040), .C0(
        n36722), .C1(n43044), .Y(n19502) );
  OR4X1 U49758 ( .A(n19510), .B(n19511), .C(n19512), .D(n19513), .Y(n36634) );
  OAI222XL U49759 ( .A0(n49542), .A1(n41797), .B0(n49526), .B1(n42729), .C0(
        n49534), .C1(n42728), .Y(n19512) );
  OAI22XL U49760 ( .A0(n41286), .A1(n42452), .B0(n36881), .B1(n19492), .Y(
        n19513) );
  OAI222XL U49761 ( .A0(n49550), .A1(n19493), .B0(n36801), .B1(n43040), .C0(
        n42496), .C1(n43044), .Y(n19510) );
  OR4X1 U49762 ( .A(n19514), .B(n19515), .C(n19516), .D(n19517), .Y(n36635) );
  OAI222XL U49763 ( .A0(n49541), .A1(n41797), .B0(n49525), .B1(n42729), .C0(
        n49533), .C1(n42728), .Y(n19516) );
  OAI22XL U49764 ( .A0(n42672), .A1(n42452), .B0(n42705), .B1(n19492), .Y(
        n19517) );
  OAI222XL U49765 ( .A0(n49549), .A1(n19493), .B0(n42569), .B1(n43040), .C0(
        n36734), .C1(n43044), .Y(n19514) );
  NOR2X2 U49766 ( .A(n9734), .B(n50146), .Y(n9679) );
  NOR3X2 U49767 ( .A(n19180), .B(n41736), .C(n19278), .Y(n19185) );
  NOR3X2 U49768 ( .A(n19180), .B(n41736), .C(n19335), .Y(n19186) );
  NAND2X2 U49769 ( .A(n19522), .B(n41796), .Y(n19493) );
  NAND2X2 U49770 ( .A(n32369), .B(n32368), .Y(n19182) );
  NAND2X1 U49771 ( .A(n19376), .B(n9742), .Y(n19335) );
  NAND2X1 U49772 ( .A(n19376), .B(n50141), .Y(n19334) );
  NAND2X1 U49773 ( .A(n19376), .B(n9715), .Y(n19239) );
  INVX1 U49774 ( .A(n41736), .Y(n50144) );
  NOR2X1 U49775 ( .A(n50134), .B(n42316), .Y(n9742) );
  CLKINVX1 U49776 ( .A(n9715), .Y(n50137) );
  CLKINVX1 U49777 ( .A(n9734), .Y(n50141) );
  NOR2XL U49778 ( .A(out_valid), .B(n41796), .Y(n9712) );
  NAND2X1 U49779 ( .A(n42316), .B(n9737), .Y(n9730) );
  AND3XL U49780 ( .A(n19335), .B(n41796), .C(n19334), .Y(n19283) );
  CLKINVX1 U49781 ( .A(n9726), .Y(n50135) );
  NOR3BX2 U49782 ( .AN(n32370), .B(n41736), .C(n19180), .Y(n19181) );
  NAND3BX1 U49783 ( .AN(n32369), .B(n19239), .C(n32368), .Y(n32370) );
  CLKBUFX3 U49784 ( .A(n19458), .Y(n41797) );
  NAND3BXL U49785 ( .AN(n9702), .B(n41796), .C(n50132), .Y(n19458) );
  CLKBUFX3 U49786 ( .A(n37592), .Y(n42321) );
  CLKBUFX3 U49787 ( .A(n37599), .Y(n42320) );
  CLKBUFX3 U49788 ( .A(n37595), .Y(n42319) );
  CLKBUFX3 U49789 ( .A(n37593), .Y(n42318) );
  CLKBUFX3 U49790 ( .A(n37601), .Y(n42317) );
  NOR4X1 U49791 ( .A(n28042), .B(n28041), .C(n28040), .D(n28039), .Y(net215825) );
  NOR4X1 U49792 ( .A(n20279), .B(n20278), .C(n20277), .D(n20276), .Y(net211155) );
  NOR4X1 U49793 ( .A(n23746), .B(n23745), .C(n23744), .D(n23743), .Y(net213350) );
  NOR4X1 U49794 ( .A(n28072), .B(n28071), .C(n28070), .D(n28069), .Y(net215834) );
  XNOR2X1 U49795 ( .A(n34248), .B(n42502), .Y(n44824) );
  NOR2X1 U49796 ( .A(n44817), .B(n44816), .Y(n44823) );
  XNOR2X1 U49797 ( .A(n36847), .B(n34002), .Y(n45668) );
  NOR2X1 U49798 ( .A(n23989), .B(n23988), .Y(n45667) );
  NOR4X1 U49799 ( .A(n23987), .B(n23986), .C(n23985), .D(n23984), .Y(n45666)
         );
  XNOR2X1 U49800 ( .A(n36859), .B(n34224), .Y(n46432) );
  NOR2X1 U49801 ( .A(n46425), .B(n46424), .Y(n46431) );
  NOR4X1 U49802 ( .A(n46429), .B(n46428), .C(n46427), .D(n46426), .Y(n46430)
         );
  NAND4X2 U49803 ( .A(n46304), .B(n46303), .C(n46302), .D(n46301), .Y(
        net209284) );
  XNOR2X1 U49804 ( .A(n36851), .B(n34160), .Y(n46303) );
  NOR2X1 U49805 ( .A(n46296), .B(n46295), .Y(n46302) );
  NOR4X1 U49806 ( .A(n46300), .B(n46299), .C(n46298), .D(n46297), .Y(n46301)
         );
  XNOR2X1 U49807 ( .A(n33938), .B(n42561), .Y(net215353) );
  XNOR2X1 U49808 ( .A(n36844), .B(n34018), .Y(n45663) );
  NOR2X1 U49809 ( .A(n23999), .B(n23998), .Y(n45662) );
  NOR4X1 U49810 ( .A(n23997), .B(n23996), .C(n23995), .D(n23994), .Y(n45661)
         );
  NAND4X2 U49811 ( .A(n44192), .B(n44191), .C(n44190), .D(n44189), .Y(n12085)
         );
  XNOR2X1 U49812 ( .A(n34002), .B(n42561), .Y(n44191) );
  NOR2X1 U49813 ( .A(n27533), .B(n27532), .Y(n44190) );
  NOR4X1 U49814 ( .A(n27531), .B(n27530), .C(n27529), .D(n27528), .Y(n44189)
         );
  NAND4X2 U49815 ( .A(n44233), .B(n44232), .C(n44231), .D(n44230), .Y(n12793)
         );
  XNOR2X1 U49816 ( .A(n33954), .B(n42561), .Y(n44232) );
  NOR2X1 U49817 ( .A(n27292), .B(n27291), .Y(n44231) );
  NOR4X1 U49818 ( .A(n27290), .B(n27289), .C(n27288), .D(n27287), .Y(n44230)
         );
  NOR4X1 U49819 ( .A(n23837), .B(n23836), .C(n23835), .D(n23834), .Y(net212694) );
  XNOR2X1 U49820 ( .A(n36847), .B(n33922), .Y(n46096) );
  NOR2X1 U49821 ( .A(n22461), .B(n22460), .Y(n46095) );
  NOR4X1 U49822 ( .A(n22459), .B(n22458), .C(n22457), .D(n22456), .Y(n46094)
         );
  XNOR2X1 U49823 ( .A(n33946), .B(n42561), .Y(net215362) );
  NOR2X1 U49824 ( .A(n23939), .B(n23938), .Y(net213364) );
  NOR4X1 U49825 ( .A(n23937), .B(n23936), .C(n23935), .D(n23934), .Y(net213365) );
  NOR4X1 U49826 ( .A(n23736), .B(n23735), .C(n23734), .D(n23733), .Y(net213345) );
  NAND4X2 U49827 ( .A(n44852), .B(n44851), .C(n44850), .D(n44849), .Y(
        net209884) );
  XNOR2X1 U49828 ( .A(n34232), .B(n42502), .Y(n44851) );
  NOR2X1 U49829 ( .A(n44844), .B(n44843), .Y(n44850) );
  NOR4X1 U49830 ( .A(n20269), .B(n20268), .C(n20267), .D(n20266), .Y(net211150) );
  NOR2X1 U49831 ( .A(n27684), .B(n27683), .Y(n43839) );
  NOR4X1 U49832 ( .A(n27682), .B(n27681), .C(n27680), .D(n27679), .Y(n43838)
         );
  NOR4X1 U49833 ( .A(n20237), .B(n20236), .C(n20235), .D(n20234), .Y(net211511) );
  NOR2X1 U49834 ( .A(n46378), .B(n46377), .Y(net212476) );
  NOR2X1 U49835 ( .A(n44875), .B(n44874), .Y(net214391) );
  NOR4X1 U49836 ( .A(n44879), .B(n44878), .C(n44877), .D(n44876), .Y(net214392) );
  NOR4X1 U49837 ( .A(n23756), .B(n23755), .C(n23754), .D(n23753), .Y(net213355) );
  XNOR2X1 U49838 ( .A(n36735), .B(n34034), .Y(n47020) );
  NOR2X1 U49839 ( .A(n20189), .B(n20187), .Y(n47019) );
  NOR4X1 U49840 ( .A(n20186), .B(n20185), .C(n20184), .D(n20183), .Y(n47018)
         );
  NOR2X1 U49841 ( .A(n46392), .B(n46391), .Y(n46398) );
  NOR4X1 U49842 ( .A(n46396), .B(n46395), .C(n46394), .D(n46393), .Y(n46397)
         );
  NOR2X1 U49843 ( .A(n44664), .B(n44663), .Y(n44670) );
  XNOR2X1 U49844 ( .A(n34184), .B(n42504), .Y(n44131) );
  NOR2X1 U49845 ( .A(n44124), .B(n44123), .Y(n44130) );
  NOR4X1 U49846 ( .A(n44128), .B(n44127), .C(n44126), .D(n44125), .Y(n44129)
         );
  NOR2X1 U49847 ( .A(n45457), .B(n45456), .Y(n45463) );
  XNOR2X1 U49848 ( .A(n34280), .B(n42505), .Y(n45376) );
  NOR2X1 U49849 ( .A(n43877), .B(n43876), .Y(n43883) );
  XNOR2X1 U49850 ( .A(n36851), .B(n34200), .Y(n46421) );
  NOR2X1 U49851 ( .A(n46414), .B(n46413), .Y(n46420) );
  NOR4X1 U49852 ( .A(n46418), .B(n46417), .C(n46416), .D(n46415), .Y(n46419)
         );
  XNOR2X1 U49853 ( .A(n34240), .B(n36737), .Y(n44793) );
  NOR2X1 U49854 ( .A(n44786), .B(n44785), .Y(n44792) );
  NOR4X1 U49855 ( .A(n44790), .B(n44789), .C(n44788), .D(n44787), .Y(n44791)
         );
  XNOR2X1 U49856 ( .A(n33930), .B(n42568), .Y(n43585) );
  NOR2X1 U49857 ( .A(n29217), .B(n29216), .Y(n43584) );
  NOR4X1 U49858 ( .A(n29215), .B(n29214), .C(n29213), .D(n29212), .Y(n43583)
         );
  NOR2X1 U49859 ( .A(n27503), .B(n27502), .Y(n44195) );
  NOR4X1 U49860 ( .A(n27501), .B(n27500), .C(n27499), .D(n27498), .Y(n44194)
         );
  XNOR2X1 U49861 ( .A(n36839), .B(n34010), .Y(n45658) );
  NOR2X1 U49862 ( .A(n24009), .B(n24008), .Y(n45657) );
  NOR4X1 U49863 ( .A(n24007), .B(n24006), .C(n24005), .D(n24004), .Y(n45656)
         );
  XNOR2X1 U49864 ( .A(n36856), .B(n34208), .Y(n46410) );
  NOR2X1 U49865 ( .A(n46403), .B(n46402), .Y(n46409) );
  NOR4X1 U49866 ( .A(n46407), .B(n46406), .C(n46405), .D(n46404), .Y(n46408)
         );
  XNOR2X1 U49867 ( .A(n33986), .B(n42561), .Y(n44210) );
  NOR2X1 U49868 ( .A(n27232), .B(n27231), .Y(n44209) );
  NOR4X1 U49869 ( .A(n27230), .B(n27229), .C(n27228), .D(n27227), .Y(n44208)
         );
  NOR4X1 U49870 ( .A(n23817), .B(n23816), .C(n23815), .D(n23814), .Y(n46180)
         );
  XNOR2X1 U49871 ( .A(n36840), .B(n33930), .Y(n46091) );
  NOR4X1 U49872 ( .A(n22469), .B(n22468), .C(n22467), .D(n22466), .Y(n46089)
         );
  XNOR2X1 U49873 ( .A(n34200), .B(n42504), .Y(n44731) );
  NOR2X1 U49874 ( .A(n44724), .B(n44723), .Y(n44730) );
  NOR4X1 U49875 ( .A(n44728), .B(n44727), .C(n44726), .D(n44725), .Y(n44729)
         );
  NOR4X1 U49876 ( .A(n23726), .B(n23725), .C(n23724), .D(n23723), .Y(n45696)
         );
  NOR2X1 U49877 ( .A(n45487), .B(n45486), .Y(net213733) );
  NOR4X1 U49878 ( .A(n23807), .B(n23806), .C(n23805), .D(n23804), .Y(n46196)
         );
  XNOR2X1 U49879 ( .A(n36858), .B(n34192), .Y(net212643) );
  XNOR2X1 U49880 ( .A(n34058), .B(n42560), .Y(net215434) );
  NOR2X1 U49881 ( .A(n46447), .B(n46446), .Y(n46453) );
  NOR4X1 U49882 ( .A(n46451), .B(n46450), .C(n46449), .D(n46448), .Y(n46452)
         );
  NOR4X1 U49883 ( .A(n46469), .B(n46468), .C(n46467), .D(n46466), .Y(net212377) );
  XNOR2X1 U49884 ( .A(n36839), .B(n33962), .Y(n47039) );
  NOR2X1 U49885 ( .A(n23718), .B(n23717), .Y(n47038) );
  NOR4X1 U49886 ( .A(n23716), .B(n23715), .C(n23714), .D(n23713), .Y(n47037)
         );
  NOR2X1 U49887 ( .A(n46223), .B(n46222), .Y(n46229) );
  NOR4X1 U49888 ( .A(n46227), .B(n46226), .C(n46225), .D(n46224), .Y(n46228)
         );
  XNOR2X1 U49889 ( .A(n34042), .B(n36846), .Y(n45673) );
  NOR2X1 U49890 ( .A(n23959), .B(n23958), .Y(n45672) );
  NOR4X1 U49891 ( .A(n23957), .B(n23956), .C(n23955), .D(n23954), .Y(n45671)
         );
  XNOR2X1 U49892 ( .A(n33970), .B(n42561), .Y(n44215) );
  NOR2X1 U49893 ( .A(n27172), .B(n27171), .Y(n44214) );
  XNOR2X1 U49894 ( .A(n34050), .B(n42560), .Y(n44185) );
  NOR2X1 U49895 ( .A(n27413), .B(n27412), .Y(n44184) );
  NOR4X1 U49896 ( .A(n27411), .B(n27410), .C(n27409), .D(n27408), .Y(n44183)
         );
  NOR2X1 U49897 ( .A(n45514), .B(n45513), .Y(net213702) );
  NOR2X1 U49898 ( .A(n23859), .B(n23858), .Y(n46191) );
  NOR4X1 U49899 ( .A(n23857), .B(n23856), .C(n23855), .D(n23854), .Y(n46190)
         );
  XNOR2X1 U49900 ( .A(n34018), .B(n42560), .Y(n44167) );
  NOR2X1 U49901 ( .A(n27593), .B(n27592), .Y(n44166) );
  NOR4X1 U49902 ( .A(n27591), .B(n27590), .C(n27589), .D(n27588), .Y(n44165)
         );
  XNOR2X1 U49903 ( .A(n36852), .B(n34288), .Y(n46363) );
  NOR2X1 U49904 ( .A(n46356), .B(n46355), .Y(n46362) );
  NOR4X1 U49905 ( .A(n46360), .B(n46359), .C(n46358), .D(n46357), .Y(n46361)
         );
  NOR4X1 U49906 ( .A(n20257), .B(n20256), .C(n20255), .D(n20254), .Y(net211521) );
  XNOR2X1 U49907 ( .A(n36847), .B(n34074), .Y(n46187) );
  NOR2X1 U49908 ( .A(n23849), .B(n23848), .Y(n46186) );
  NOR4X1 U49909 ( .A(n23847), .B(n23846), .C(n23845), .D(n23844), .Y(n46185)
         );
  NAND4X1 U49910 ( .A(n45709), .B(n45708), .C(n45707), .D(n45706), .Y(n11130)
         );
  XNOR2X1 U49911 ( .A(n36838), .B(n33946), .Y(n45708) );
  NOR2X1 U49912 ( .A(n23698), .B(n23697), .Y(n45707) );
  NOR4X1 U49913 ( .A(n23696), .B(n23695), .C(n23694), .D(n23693), .Y(n45706)
         );
  XNOR2X1 U49914 ( .A(n36746), .B(n33932), .Y(n47241) );
  NOR2X1 U49915 ( .A(n19608), .B(n19607), .Y(n47240) );
  XNOR2X1 U49916 ( .A(n36854), .B(n34232), .Y(n46443) );
  NOR2X1 U49917 ( .A(n46436), .B(n46435), .Y(n46442) );
  NOR4X1 U49918 ( .A(n46440), .B(n46439), .C(n46438), .D(n46437), .Y(n46441)
         );
  XNOR2X1 U49919 ( .A(n36859), .B(n34256), .Y(net212386) );
  NOR2X1 U49920 ( .A(n46458), .B(n46457), .Y(net212387) );
  NOR4X1 U49921 ( .A(n46462), .B(n46461), .C(n46460), .D(n46459), .Y(net212388) );
  NOR2X1 U49922 ( .A(n46334), .B(n46333), .Y(n46340) );
  NOR4X1 U49923 ( .A(n46338), .B(n46337), .C(n46336), .D(n46335), .Y(n46339)
         );
  NOR2X1 U49924 ( .A(n46367), .B(n46366), .Y(n46373) );
  NOR4X1 U49925 ( .A(n46371), .B(n46370), .C(n46369), .D(n46368), .Y(n46372)
         );
  XOR2X1 U49926 ( .A(n36742), .B(n34364), .Y(n47605) );
  XOR2X1 U49927 ( .A(n36918), .B(n34308), .Y(n46314) );
  XOR2X1 U49928 ( .A(n36741), .B(n34300), .Y(n47318) );
  XOR2X1 U49929 ( .A(n36748), .B(n34268), .Y(n47373) );
  XOR2X1 U49930 ( .A(n36717), .B(n34309), .Y(n47310) );
  NOR2X1 U49931 ( .A(n43970), .B(n43969), .Y(n43976) );
  NOR3X1 U49932 ( .A(n46508), .B(n46507), .C(n46506), .Y(n46509) );
  XNOR2X1 U49933 ( .A(n36857), .B(n34304), .Y(n46330) );
  NOR2X1 U49934 ( .A(n46323), .B(n46322), .Y(n46329) );
  XOR2X1 U49935 ( .A(n36907), .B(n34122), .Y(n43861) );
  NOR2X1 U49936 ( .A(n45338), .B(n45337), .Y(n45344) );
  NOR4X1 U49937 ( .A(n45342), .B(n45341), .C(n45340), .D(n45339), .Y(n45343)
         );
  NOR2X1 U49938 ( .A(n46212), .B(n46211), .Y(n46218) );
  NOR4X1 U49939 ( .A(n46216), .B(n46215), .C(n46214), .D(n46213), .Y(n46217)
         );
  NOR2X1 U49940 ( .A(n27142), .B(n27141), .Y(n44219) );
  NOR4X1 U49941 ( .A(n27140), .B(n27139), .C(n27138), .D(n27137), .Y(n44218)
         );
  XOR2X1 U49942 ( .A(n34404), .B(n42699), .Y(n45094) );
  XOR2X1 U49943 ( .A(n41299), .B(n34420), .Y(n46601) );
  NOR2X1 U49944 ( .A(n44001), .B(n44000), .Y(n44007) );
  NOR4X1 U49945 ( .A(n44005), .B(n44004), .C(n44003), .D(n44002), .Y(n44006)
         );
  XOR2X1 U49946 ( .A(n9657), .B(n41641), .Y(n45264) );
  XOR2X1 U49947 ( .A(n9659), .B(n36875), .Y(n45263) );
  XOR2X1 U49948 ( .A(n34429), .B(n42632), .Y(n45262) );
  NOR2X1 U49949 ( .A(n43939), .B(n43938), .Y(n43945) );
  NOR4X1 U49950 ( .A(n43943), .B(n43942), .C(n43941), .D(n43940), .Y(n43944)
         );
  XOR2X1 U49951 ( .A(n42066), .B(n36885), .Y(n44893) );
  XOR2X1 U49952 ( .A(n42073), .B(n36883), .Y(n45181) );
  XNOR2X1 U49953 ( .A(n36847), .B(n34058), .Y(n47000) );
  NOR2X1 U49954 ( .A(n23979), .B(n23978), .Y(n46999) );
  NOR4X1 U49955 ( .A(n23977), .B(n23976), .C(n23975), .D(n23974), .Y(n46998)
         );
  XOR2X1 U49956 ( .A(n41333), .B(n34317), .Y(n46345) );
  XOR2X1 U49957 ( .A(n36715), .B(n34301), .Y(n47316) );
  NOR4X1 U49958 ( .A(n20227), .B(n20226), .C(n20225), .D(n20224), .Y(net211526) );
  NOR2X1 U49959 ( .A(n47512), .B(n47511), .Y(n47518) );
  NOR2X1 U49960 ( .A(n27714), .B(n27713), .Y(n43852) );
  NOR4X1 U49961 ( .A(n27712), .B(n27711), .C(n27710), .D(n27709), .Y(n43851)
         );
  XNOR2X1 U49962 ( .A(n36846), .B(n34106), .Y(n46203) );
  NOR2X1 U49963 ( .A(n23779), .B(n23778), .Y(n46202) );
  NOR4X1 U49964 ( .A(n23777), .B(n23776), .C(n23775), .D(n23774), .Y(n46201)
         );
  XNOR2X1 U49965 ( .A(n36841), .B(n34178), .Y(n46243) );
  NOR4X1 U49966 ( .A(n46389), .B(n46388), .C(n46387), .D(n46386), .Y(net212466) );
  XOR2X1 U49967 ( .A(n9665), .B(net219330), .Y(n45265) );
  NAND4X1 U49968 ( .A(n47016), .B(n47015), .C(n47014), .D(n47013), .Y(n11441)
         );
  XNOR2X1 U49969 ( .A(n36735), .B(n34042), .Y(n47015) );
  NOR2X1 U49970 ( .A(n20199), .B(n20198), .Y(n47014) );
  NOR4X1 U49971 ( .A(n20197), .B(n20196), .C(n20195), .D(n20194), .Y(n47013)
         );
  XNOR2X1 U49972 ( .A(n36860), .B(n34184), .Y(n46240) );
  XNOR2X1 U49973 ( .A(n42471), .B(n34384), .Y(n47659) );
  XNOR2X1 U49974 ( .A(n36734), .B(n34050), .Y(n47005) );
  NOR2X1 U49975 ( .A(n20209), .B(n20208), .Y(n47004) );
  NOR4X1 U49976 ( .A(n20207), .B(n20206), .C(n20205), .D(n20204), .Y(n47003)
         );
  XNOR2X1 U49977 ( .A(n42471), .B(n34360), .Y(n47632) );
  NOR2X1 U49978 ( .A(n47625), .B(n47624), .Y(n47631) );
  NOR4X1 U49979 ( .A(n47629), .B(n47628), .C(n47627), .D(n47626), .Y(n47630)
         );
  XOR2X1 U49980 ( .A(n36918), .B(n34372), .Y(n46475) );
  NAND4X1 U49981 ( .A(n47891), .B(n47890), .C(n47889), .D(n47888), .Y(n12967)
         );
  XNOR2X1 U49982 ( .A(n36734), .B(n33970), .Y(n47890) );
  NOR2X1 U49983 ( .A(n20177), .B(n20176), .Y(n47889) );
  NOR4X1 U49984 ( .A(n20175), .B(n20174), .C(n20173), .D(n20172), .Y(n47888)
         );
  NOR2X1 U49985 ( .A(n44155), .B(n44154), .Y(n44161) );
  NOR4X1 U49986 ( .A(n44159), .B(n44158), .C(n44157), .D(n44156), .Y(n44160)
         );
  NOR2X1 U49987 ( .A(n23708), .B(n23707), .Y(n45702) );
  NOR4X1 U49988 ( .A(n23706), .B(n23705), .C(n23704), .D(n23703), .Y(n45701)
         );
  XNOR2X1 U49989 ( .A(n42473), .B(n34280), .Y(n47356) );
  NOR2X1 U49990 ( .A(n47349), .B(n47348), .Y(n47355) );
  NOR2X1 U49991 ( .A(n47459), .B(n47458), .Y(n47465) );
  NOR3X1 U49992 ( .A(n46476), .B(n46475), .C(n46474), .Y(n46477) );
  NOR2X1 U49993 ( .A(n47603), .B(n47602), .Y(n47609) );
  NOR4X1 U49994 ( .A(n47607), .B(n47606), .C(n47605), .D(n47604), .Y(n47608)
         );
  XNOR2X1 U49995 ( .A(n34034), .B(n36845), .Y(n45683) );
  NOR2X1 U49996 ( .A(n23949), .B(n23948), .Y(n45682) );
  NOR4X1 U49997 ( .A(n23947), .B(n23946), .C(n23945), .D(n23944), .Y(n45681)
         );
  XNOR2X1 U49998 ( .A(n34168), .B(n42504), .Y(n44069) );
  NOR2X1 U49999 ( .A(n44062), .B(n44061), .Y(n44068) );
  NOR2X1 U50000 ( .A(n27262), .B(n27261), .Y(n44204) );
  NOR4X1 U50001 ( .A(n27260), .B(n27259), .C(n27258), .D(n27257), .Y(n44203)
         );
  NOR2X1 U50002 ( .A(n45400), .B(n45399), .Y(n45406) );
  NOR2X1 U50003 ( .A(n44093), .B(n44092), .Y(n44099) );
  NOR4X1 U50004 ( .A(n44097), .B(n44096), .C(n44095), .D(n44094), .Y(n44098)
         );
  NOR2X1 U50005 ( .A(n44695), .B(n44694), .Y(n44701) );
  NOR4X1 U50006 ( .A(n44699), .B(n44698), .C(n44697), .D(n44696), .Y(n44700)
         );
  NOR2X1 U50007 ( .A(n27984), .B(n27983), .Y(n43831) );
  NOR4X1 U50008 ( .A(n27982), .B(n27981), .C(n27980), .D(n27979), .Y(n43830)
         );
  NOR2X1 U50009 ( .A(n44755), .B(n44754), .Y(n44761) );
  NOR4X1 U50010 ( .A(n44759), .B(n44758), .C(n44757), .D(n44756), .Y(n44760)
         );
  NOR2X1 U50011 ( .A(n43908), .B(n43907), .Y(n43914) );
  NOR2X1 U50012 ( .A(n46262), .B(n46261), .Y(n46268) );
  NOR4X1 U50013 ( .A(n46266), .B(n46265), .C(n46264), .D(n46263), .Y(n46267)
         );
  XNOR2X1 U50014 ( .A(n36845), .B(n34050), .Y(n47010) );
  NOR2X1 U50015 ( .A(n23969), .B(n23968), .Y(n47009) );
  NOR4X1 U50016 ( .A(n23967), .B(n23966), .C(n23965), .D(n23964), .Y(n47008)
         );
  NOR2X1 U50017 ( .A(n47636), .B(n47635), .Y(n47642) );
  NOR4X1 U50018 ( .A(n47640), .B(n47639), .C(n47638), .D(n47637), .Y(n47641)
         );
  XNOR2X1 U50019 ( .A(n36850), .B(n34312), .Y(n46319) );
  NOR2X1 U50020 ( .A(n46312), .B(n46311), .Y(n46318) );
  NOR4X1 U50021 ( .A(n46316), .B(n46315), .C(n46314), .D(n46313), .Y(n46317)
         );
  XNOR2X1 U50022 ( .A(n34026), .B(n42560), .Y(n44176) );
  NOR2X1 U50023 ( .A(n27563), .B(n27562), .Y(n44175) );
  NOR4X1 U50024 ( .A(n27561), .B(n27560), .C(n27559), .D(n27558), .Y(n44174)
         );
  NOR2X1 U50025 ( .A(n47426), .B(n47425), .Y(n47432) );
  NOR4X1 U50026 ( .A(n47430), .B(n47429), .C(n47428), .D(n47427), .Y(n47431)
         );
  NOR2X1 U50027 ( .A(n45219), .B(n45218), .Y(n45225) );
  XNOR2X1 U50028 ( .A(n34344), .B(n36737), .Y(n45135) );
  NOR2X1 U50029 ( .A(n45128), .B(n45127), .Y(n45134) );
  NOR2X1 U50030 ( .A(n46524), .B(n46523), .Y(n46530) );
  NOR4X1 U50031 ( .A(n46528), .B(n46527), .C(n46526), .D(n46525), .Y(n46529)
         );
  XOR2X1 U50032 ( .A(n34417), .B(n42718), .Y(n45003) );
  XOR2X1 U50033 ( .A(n34404), .B(n36824), .Y(n44999) );
  XOR2X1 U50034 ( .A(n9662), .B(net219468), .Y(n45244) );
  XOR2X1 U50035 ( .A(n9669), .B(n42638), .Y(n45240) );
  XOR2X1 U50036 ( .A(n34400), .B(n42592), .Y(n45082) );
  XOR2X1 U50037 ( .A(n34320), .B(n34450), .Y(n45437) );
  XOR2X1 U50038 ( .A(n9655), .B(n42660), .Y(n45241) );
  XOR2X1 U50039 ( .A(n9663), .B(n42597), .Y(n45237) );
  XOR2X1 U50040 ( .A(n34316), .B(n36822), .Y(n45410) );
  XOR2X1 U50041 ( .A(n34427), .B(n41323), .Y(n45233) );
  XOR2X1 U50042 ( .A(n34400), .B(n36731), .Y(n45056) );
  XOR2X1 U50043 ( .A(n34408), .B(n36730), .Y(n44996) );
  XOR2X1 U50044 ( .A(n34185), .B(n42577), .Y(n44157) );
  XOR2X1 U50045 ( .A(n34420), .B(n41385), .Y(n45006) );
  XOR2X1 U50046 ( .A(n9655), .B(n36881), .Y(n45259) );
  XOR2X1 U50047 ( .A(n9667), .B(n42628), .Y(n45239) );
  XOR2X1 U50048 ( .A(n34405), .B(n41282), .Y(n45093) );
  XOR2X1 U50049 ( .A(n34393), .B(n36905), .Y(n45089) );
  XOR2X1 U50050 ( .A(n34428), .B(n36822), .Y(n45235) );
  XOR2X1 U50051 ( .A(n34305), .B(n41319), .Y(n45473) );
  XOR2X1 U50052 ( .A(n34325), .B(n41282), .Y(n45448) );
  XOR2X1 U50053 ( .A(n34317), .B(n42628), .Y(n45440) );
  XOR2X1 U50054 ( .A(n34220), .B(n36823), .Y(n44698) );
  XOR2X1 U50055 ( .A(n34204), .B(n36828), .Y(n44758) );
  XOR2X1 U50056 ( .A(n34322), .B(n41630), .Y(n45192) );
  XOR2X1 U50057 ( .A(n9666), .B(net219310), .Y(n45246) );
  XOR2X1 U50058 ( .A(n9665), .B(n42615), .Y(n45238) );
  XOR2X1 U50059 ( .A(n34156), .B(n36828), .Y(n43942) );
  XOR2X1 U50060 ( .A(n34244), .B(n36821), .Y(n44820) );
  XOR2X1 U50061 ( .A(n34228), .B(n36824), .Y(n44847) );
  XOR2X1 U50062 ( .A(n34236), .B(n36822), .Y(n44789) );
  XOR2X1 U50063 ( .A(n34306), .B(n42672), .Y(n45472) );
  XOR2X1 U50064 ( .A(n34310), .B(n41284), .Y(n45468) );
  XOR2X1 U50065 ( .A(n34402), .B(n42557), .Y(n45001) );
  XOR2X1 U50066 ( .A(n34405), .B(n36832), .Y(n44997) );
  NOR4X1 U50067 ( .A(n27200), .B(n27199), .C(n27198), .D(n27197), .Y(net215373) );
  XNOR2X1 U50068 ( .A(n34272), .B(n42505), .Y(n45318) );
  NOR2X1 U50069 ( .A(n45311), .B(n45310), .Y(n45317) );
  NOR4X1 U50070 ( .A(n45315), .B(n45314), .C(n45313), .D(n45312), .Y(n45316)
         );
  NOR2X1 U50071 ( .A(n47470), .B(n47469), .Y(n47476) );
  NOR4X1 U50072 ( .A(n47474), .B(n47473), .C(n47472), .D(n47471), .Y(n47475)
         );
  NOR2X1 U50073 ( .A(n47393), .B(n47392), .Y(n47399) );
  XOR2X1 U50074 ( .A(n9658), .B(n42705), .Y(n45250) );
  XOR2X1 U50075 ( .A(n9656), .B(n36886), .Y(n45249) );
  NOR2X1 U50076 ( .A(n45188), .B(n45187), .Y(n45194) );
  NOR4X2 U50077 ( .A(n45192), .B(n45191), .C(n45190), .D(n45189), .Y(n45193)
         );
  XNOR2X1 U50078 ( .A(n36734), .B(n34082), .Y(n47284) );
  NOR2X1 U50079 ( .A(n20301), .B(n20300), .Y(n47283) );
  NOR4X1 U50080 ( .A(n20299), .B(n20298), .C(n20297), .D(n20296), .Y(n47282)
         );
  XOR2X1 U50081 ( .A(n34401), .B(n34435), .Y(n45097) );
  XOR2X1 U50082 ( .A(n34402), .B(n42704), .Y(n45096) );
  XOR2X1 U50083 ( .A(n42065), .B(n36883), .Y(n45095) );
  XNOR2X1 U50084 ( .A(n34352), .B(n36737), .Y(n45166) );
  NOR2X1 U50085 ( .A(n45159), .B(n45158), .Y(n45165) );
  NOR4X1 U50086 ( .A(n45163), .B(n45162), .C(n45161), .D(n45160), .Y(n45164)
         );
  NOR2X1 U50087 ( .A(n46513), .B(n46512), .Y(n46519) );
  XNOR2X1 U50088 ( .A(n34378), .B(n42560), .Y(n44900) );
  XOR2X1 U50089 ( .A(n42089), .B(n36887), .Y(n44717) );
  XOR2X1 U50090 ( .A(n42083), .B(n36886), .Y(n44808) );
  XOR2X1 U50091 ( .A(n42078), .B(n36882), .Y(n45391) );
  XOR2X1 U50092 ( .A(n42071), .B(n36880), .Y(n45121) );
  XOR2X1 U50093 ( .A(n42079), .B(n36889), .Y(n45360) );
  XOR2X1 U50094 ( .A(n42080), .B(n36879), .Y(n45302) );
  XOR2X1 U50095 ( .A(n42075), .B(n36881), .Y(n45450) );
  XOR2X1 U50096 ( .A(n42085), .B(n36888), .Y(n44839) );
  NOR4X1 U50097 ( .A(n44086), .B(n44085), .C(n44084), .D(n44083), .Y(n44087)
         );
  NOR4X1 U50098 ( .A(n44117), .B(n44116), .C(n44115), .D(n44114), .Y(n44118)
         );
  XOR2X1 U50099 ( .A(n34193), .B(n42717), .Y(n44117) );
  XOR2X1 U50100 ( .A(n34194), .B(n41642), .Y(n44116) );
  XOR2X1 U50101 ( .A(n42091), .B(n36882), .Y(n44115) );
  NOR4X1 U50102 ( .A(n44688), .B(n44687), .C(n44686), .D(n44685), .Y(n44689)
         );
  NOR4X1 U50103 ( .A(n43963), .B(n43962), .C(n43961), .D(n43960), .Y(n43964)
         );
  XOR2X1 U50104 ( .A(n34161), .B(n42717), .Y(n43963) );
  XOR2X1 U50105 ( .A(n34162), .B(n41641), .Y(n43962) );
  XOR2X1 U50106 ( .A(n42095), .B(n36889), .Y(n43961) );
  NOR4X1 U50107 ( .A(n43901), .B(n43900), .C(n43899), .D(n43898), .Y(n43902)
         );
  NOR4X1 U50108 ( .A(n43994), .B(n43993), .C(n43992), .D(n43991), .Y(n43995)
         );
  XOR2X1 U50109 ( .A(n34153), .B(n34435), .Y(n43994) );
  NOR4X1 U50110 ( .A(n43932), .B(n43931), .C(n43930), .D(n43929), .Y(n43933)
         );
  NOR4X1 U50111 ( .A(n44025), .B(n44024), .C(n44023), .D(n44022), .Y(n44026)
         );
  XOR2X1 U50112 ( .A(n34145), .B(n42717), .Y(n44025) );
  XOR2X1 U50113 ( .A(n34146), .B(n41642), .Y(n44024) );
  XOR2X1 U50114 ( .A(n42097), .B(n36889), .Y(n44023) );
  NOR4X1 U50115 ( .A(n44055), .B(n44054), .C(n44053), .D(n44052), .Y(n44056)
         );
  XOR2X1 U50116 ( .A(n34177), .B(n42717), .Y(n44055) );
  XOR2X1 U50117 ( .A(n34178), .B(n42707), .Y(n44054) );
  XOR2X1 U50118 ( .A(n42093), .B(n36886), .Y(n44053) );
  XNOR2X1 U50119 ( .A(n34388), .B(n36822), .Y(n45099) );
  XNOR2X1 U50120 ( .A(n34380), .B(n36825), .Y(n44901) );
  XOR2X1 U50121 ( .A(n34044), .B(n36827), .Y(n45676) );
  XNOR2X1 U50122 ( .A(n34384), .B(n36730), .Y(n44907) );
  XNOR2X1 U50123 ( .A(n34392), .B(n42505), .Y(n45105) );
  XNOR2X1 U50124 ( .A(n36850), .B(n34352), .Y(n46553) );
  NOR2X1 U50125 ( .A(n46546), .B(n46545), .Y(n46552) );
  NOR4X1 U50126 ( .A(n46550), .B(n46549), .C(n46548), .D(n46547), .Y(n46551)
         );
  NOR2X1 U50127 ( .A(n46491), .B(n46490), .Y(n46497) );
  NOR4X1 U50128 ( .A(n46495), .B(n46494), .C(n46493), .D(n46492), .Y(n46496)
         );
  NOR2X1 U50129 ( .A(n47295), .B(n47294), .Y(n47301) );
  NOR4X1 U50130 ( .A(n47299), .B(n47298), .C(n47297), .D(n47296), .Y(n47300)
         );
  XNOR2X1 U50131 ( .A(n36853), .B(n34320), .Y(n46352) );
  NOR2X1 U50132 ( .A(n46345), .B(n46344), .Y(n46351) );
  NOR4X1 U50133 ( .A(n46349), .B(n46348), .C(n46347), .D(n46346), .Y(n46350)
         );
  XNOR2X1 U50134 ( .A(n42471), .B(n34376), .Y(n47621) );
  NOR2X1 U50135 ( .A(n47614), .B(n47613), .Y(n47620) );
  XNOR2X1 U50136 ( .A(n36734), .B(n33978), .Y(n47895) );
  NOR2X1 U50137 ( .A(n20167), .B(n20166), .Y(n47894) );
  NOR4X1 U50138 ( .A(n20165), .B(n20164), .C(n20163), .D(n20162), .Y(n47893)
         );
  NOR4X1 U50139 ( .A(n47320), .B(n47319), .C(n47318), .D(n47317), .Y(n47321)
         );
  NOR2X1 U50140 ( .A(n47592), .B(n47591), .Y(n47598) );
  NOR2X1 U50141 ( .A(n47569), .B(n47568), .Y(n47575) );
  NOR4X1 U50142 ( .A(n47573), .B(n47572), .C(n47571), .D(n47570), .Y(n47574)
         );
  NOR2X1 U50143 ( .A(n47481), .B(n47480), .Y(n47487) );
  XNOR2X1 U50144 ( .A(n36736), .B(n34098), .Y(n47555) );
  NOR2X1 U50145 ( .A(n20393), .B(n20392), .Y(n47554) );
  NOR4X1 U50146 ( .A(n20391), .B(n20390), .C(n20389), .D(n20388), .Y(n47553)
         );
  XNOR2X1 U50147 ( .A(n42472), .B(n34296), .Y(n47334) );
  NOR2X1 U50148 ( .A(n47327), .B(n47326), .Y(n47333) );
  NOR2X1 U50149 ( .A(n47371), .B(n47370), .Y(n47377) );
  NOR4X1 U50150 ( .A(n47375), .B(n47374), .C(n47373), .D(n47372), .Y(n47376)
         );
  NOR2X1 U50151 ( .A(n46535), .B(n46534), .Y(n46541) );
  NOR2X1 U50152 ( .A(n47523), .B(n47522), .Y(n47529) );
  NOR4X1 U50153 ( .A(n47527), .B(n47526), .C(n47525), .D(n47524), .Y(n47528)
         );
  NAND4X1 U50154 ( .A(n47561), .B(n47560), .C(n47559), .D(n47558), .Y(n48037)
         );
  NOR2X1 U50155 ( .A(n20403), .B(n20402), .Y(n47559) );
  NOR4X1 U50156 ( .A(n20401), .B(n20400), .C(n20399), .D(n20398), .Y(n47558)
         );
  XNOR2X1 U50157 ( .A(n36733), .B(n34058), .Y(n46995) );
  NOR2X1 U50158 ( .A(n20219), .B(n20218), .Y(n46994) );
  NOR4X1 U50159 ( .A(n20217), .B(n20216), .C(n20215), .D(n20214), .Y(n46993)
         );
  NOR4X1 U50160 ( .A(n20145), .B(n20144), .C(n20143), .D(n20142), .Y(n47032)
         );
  NOR2X1 U50161 ( .A(n44986), .B(n44985), .Y(n44992) );
  NAND4X1 U50162 ( .A(n47030), .B(n47029), .C(n47028), .D(n47027), .Y(
        net210142) );
  XNOR2X1 U50163 ( .A(n36746), .B(n33988), .Y(n47029) );
  NOR2X1 U50164 ( .A(n20157), .B(n20156), .Y(n47028) );
  NOR4X1 U50165 ( .A(n20155), .B(n20154), .C(n20153), .D(n20152), .Y(n47027)
         );
  NOR2X1 U50166 ( .A(n47581), .B(n47580), .Y(n47587) );
  NOR2X1 U50167 ( .A(n47338), .B(n47337), .Y(n47344) );
  NOR4X1 U50168 ( .A(n47342), .B(n47341), .C(n47340), .D(n47339), .Y(n47343)
         );
  NOR2X1 U50169 ( .A(n47360), .B(n47359), .Y(n47366) );
  XNOR2X1 U50170 ( .A(n36857), .B(n34176), .Y(n46258) );
  NOR2X1 U50171 ( .A(n46251), .B(n46250), .Y(n46257) );
  NOR2X1 U50172 ( .A(n47448), .B(n47447), .Y(n47454) );
  NOR4X1 U50173 ( .A(n47452), .B(n47451), .C(n47450), .D(n47449), .Y(n47453)
         );
  NOR2X1 U50174 ( .A(n47382), .B(n47381), .Y(n47388) );
  NOR4X1 U50175 ( .A(n47386), .B(n47385), .C(n47384), .D(n47383), .Y(n47387)
         );
  NOR2X1 U50176 ( .A(n47404), .B(n47403), .Y(n47410) );
  NOR4X1 U50177 ( .A(n47408), .B(n47407), .C(n47406), .D(n47405), .Y(n47409)
         );
  XNOR2X1 U50178 ( .A(n42472), .B(n34176), .Y(n47499) );
  NOR2X1 U50179 ( .A(n47492), .B(n47491), .Y(n47498) );
  NOR4X1 U50180 ( .A(n47496), .B(n47495), .C(n47494), .D(n47493), .Y(n47497)
         );
  NOR2X1 U50181 ( .A(n47534), .B(n47533), .Y(n47540) );
  NOR4X1 U50182 ( .A(n47538), .B(n47537), .C(n47536), .D(n47535), .Y(n47539)
         );
  NOR4X1 U50183 ( .A(n20289), .B(n20288), .C(n20287), .D(n20286), .Y(n47287)
         );
  XNOR2X1 U50184 ( .A(n42472), .B(n34248), .Y(n47444) );
  NOR2X1 U50185 ( .A(n47437), .B(n47436), .Y(n47443) );
  NOR4X1 U50186 ( .A(n47441), .B(n47440), .C(n47439), .D(n47438), .Y(n47442)
         );
  NOR2X1 U50187 ( .A(n47415), .B(n47414), .Y(n47421) );
  NOR4X1 U50188 ( .A(n45235), .B(n45234), .C(n45233), .D(n45232), .Y(n45255)
         );
  XOR2X1 U50189 ( .A(n34425), .B(n42576), .Y(n45232) );
  NOR4X1 U50190 ( .A(n47704), .B(n47703), .C(n47702), .D(n47701), .Y(n47706)
         );
  NOR4X1 U50191 ( .A(n47508), .B(n47507), .C(n47506), .D(n47505), .Y(n47509)
         );
  XOR2X1 U50192 ( .A(n36736), .B(n34162), .Y(n47503) );
  XOR2X1 U50193 ( .A(n34068), .B(n36821), .Y(n43819) );
  XOR2X1 U50194 ( .A(n41303), .B(n34060), .Y(n46997) );
  NOR2X1 U50195 ( .A(n10393), .B(n44193), .Y(n44197) );
  XOR2X1 U50196 ( .A(n34060), .B(n36828), .Y(n44187) );
  XOR2X1 U50197 ( .A(n34052), .B(n36822), .Y(n44182) );
  XOR2X1 U50198 ( .A(n33993), .B(n36776), .Y(n45692) );
  NOR2X1 U50199 ( .A(n10879), .B(n47024), .Y(net211513) );
  NOR2X1 U50200 ( .A(n10567), .B(n45695), .Y(n45699) );
  NOR2X1 U50201 ( .A(n10382), .B(n44223), .Y(net215361) );
  NOR2X1 U50202 ( .A(n10383), .B(n44217), .Y(n44221) );
  NOR4X1 U50203 ( .A(n46600), .B(n46599), .C(n46598), .D(n46597), .Y(net212212) );
  NOR4X1 U50204 ( .A(n46604), .B(n46603), .C(n46602), .D(n46601), .Y(net212213) );
  NOR2X1 U50205 ( .A(n11770), .B(n44202), .Y(n44206) );
  NOR2X1 U50206 ( .A(n12749), .B(n45665), .Y(n45669) );
  XOR2X1 U50207 ( .A(n34084), .B(n36823), .Y(n43820) );
  NOR2X1 U50208 ( .A(n11131), .B(n47238), .Y(n47242) );
  XOR2X1 U50209 ( .A(n34049), .B(n36782), .Y(n47007) );
  NOR4X1 U50210 ( .A(n46594), .B(n46593), .C(n46592), .D(n46591), .Y(n46596)
         );
  XOR2X1 U50211 ( .A(n36916), .B(n34398), .Y(n46590) );
  XOR2X1 U50212 ( .A(n33972), .B(n36824), .Y(n44212) );
  XOR2X1 U50213 ( .A(n34073), .B(n36786), .Y(n46184) );
  NOR2X1 U50214 ( .A(n12744), .B(n45700), .Y(n45704) );
  XOR2X1 U50215 ( .A(n41305), .B(n33972), .Y(n45700) );
  XOR2X1 U50216 ( .A(n41303), .B(n33956), .Y(n45691) );
  NOR2X1 U50217 ( .A(n47023), .B(net209268), .Y(net211518) );
  NOR2X1 U50218 ( .A(n43818), .B(net210460), .Y(net215831) );
  XOR2X1 U50219 ( .A(n34076), .B(n36824), .Y(n43818) );
  NOR2X1 U50220 ( .A(n46501), .B(n46500), .Y(n46502) );
  XOR2X1 U50221 ( .A(n36913), .B(n34365), .Y(n46501) );
  XOR2X1 U50222 ( .A(n41295), .B(n34366), .Y(n46500) );
  AND2X2 U50223 ( .A(n41792), .B(n41793), .Y(n46470) );
  XNOR2X1 U50224 ( .A(n41328), .B(n34373), .Y(n41792) );
  XNOR2X1 U50225 ( .A(n41290), .B(n34374), .Y(n41793) );
  AND2X2 U50226 ( .A(n41794), .B(n41795), .Y(n46479) );
  NAND3X1 U50227 ( .A(n47691), .B(n47690), .C(n47689), .Y(n47692) );
  XNOR2X1 U50228 ( .A(n36795), .B(n34390), .Y(n47690) );
  XNOR2X1 U50229 ( .A(n42496), .B(n42067), .Y(n47689) );
  XOR2X1 U50230 ( .A(n34404), .B(n42637), .Y(n45067) );
  NOR4X1 U50231 ( .A(n24088), .B(n24087), .C(n24086), .D(n24085), .Y(net212729) );
  XNOR2X1 U50232 ( .A(n33746), .B(n42562), .Y(net215232) );
  NOR2X1 U50233 ( .A(n26660), .B(n26659), .Y(net215233) );
  NOR4X1 U50234 ( .A(n29275), .B(n29274), .C(n29273), .D(n29272), .Y(net216023) );
  NOR4X1 U50235 ( .A(n24160), .B(n24159), .C(n24158), .D(n24157), .Y(net212744) );
  NOR4X1 U50236 ( .A(n26929), .B(n26928), .C(n26927), .D(n26926), .Y(net215292) );
  NOR4X1 U50237 ( .A(n26808), .B(n26807), .C(n26806), .D(n26805), .Y(net215207) );
  NOR4X1 U50238 ( .A(n24078), .B(n24077), .C(n24076), .D(n24075), .Y(net212719) );
  NOR4X1 U50239 ( .A(n22439), .B(n22438), .C(n22437), .D(n22436), .Y(n46104)
         );
  NOR4X1 U50240 ( .A(n26868), .B(n26867), .C(n26866), .D(n26865), .Y(net215225) );
  NOR4X1 U50241 ( .A(n24018), .B(n24017), .C(n24016), .D(n24015), .Y(net213405) );
  NOR4X1 U50242 ( .A(n22389), .B(n22388), .C(n22387), .D(n22386), .Y(n46139)
         );
  XNOR2X1 U50243 ( .A(n36771), .B(n33921), .Y(n47246) );
  NOR2X1 U50244 ( .A(n19598), .B(n19597), .Y(n47245) );
  XNOR2X1 U50245 ( .A(n36746), .B(n33732), .Y(n47157) );
  NOR2X1 U50246 ( .A(n19811), .B(n19810), .Y(n47156) );
  NOR4X1 U50247 ( .A(n24068), .B(n24067), .C(n24066), .D(n24065), .Y(net212714) );
  NOR4X1 U50248 ( .A(n24170), .B(n24169), .C(n24168), .D(n24167), .Y(net212739) );
  XNOR2X1 U50249 ( .A(n33826), .B(n42568), .Y(n43651) );
  NOR2X1 U50250 ( .A(n29096), .B(n29095), .Y(n43650) );
  NOR4X1 U50251 ( .A(n29094), .B(n29093), .C(n29092), .D(n29091), .Y(n43649)
         );
  NOR4X1 U50252 ( .A(n24150), .B(n24149), .C(n24148), .D(n24147), .Y(net212734) );
  NOR4X1 U50253 ( .A(n29245), .B(n29244), .C(n29243), .D(n29242), .Y(net216050) );
  XNOR2X1 U50254 ( .A(n33858), .B(n42568), .Y(n43576) );
  NOR2X1 U50255 ( .A(n29367), .B(n29366), .Y(n43575) );
  NOR4X1 U50256 ( .A(n29365), .B(n29364), .C(n29363), .D(n29362), .Y(n43574)
         );
  NOR4X1 U50257 ( .A(n26959), .B(n26958), .C(n26957), .D(n26956), .Y(net215301) );
  NAND4X2 U50258 ( .A(n44276), .B(n44275), .C(n44274), .D(n44273), .Y(n12150)
         );
  XNOR2X1 U50259 ( .A(n33714), .B(n42562), .Y(n44275) );
  NOR2X1 U50260 ( .A(n26991), .B(n26990), .Y(n44274) );
  NOR4X1 U50261 ( .A(n26989), .B(n26988), .C(n26987), .D(n26986), .Y(n44273)
         );
  NOR4X1 U50262 ( .A(n26899), .B(n26898), .C(n26897), .D(n26896), .Y(net215274) );
  XNOR2X1 U50263 ( .A(n36843), .B(n33810), .Y(n46166) );
  NOR2X1 U50264 ( .A(n22321), .B(n22320), .Y(n46165) );
  NOR4X1 U50265 ( .A(n22319), .B(n22318), .C(n22317), .D(n22316), .Y(n46164)
         );
  NOR4X1 U50266 ( .A(n24119), .B(n24118), .C(n24117), .D(n24116), .Y(n45624)
         );
  NAND4X1 U50267 ( .A(n43563), .B(n43562), .C(n43561), .D(n43560), .Y(n12146)
         );
  XNOR2X1 U50268 ( .A(n33842), .B(n42568), .Y(n43562) );
  NOR2X1 U50269 ( .A(n29427), .B(n29426), .Y(n43561) );
  NOR4X1 U50270 ( .A(n29425), .B(n29424), .C(n29423), .D(n29422), .Y(n43560)
         );
  XNOR2X1 U50271 ( .A(n36847), .B(n33690), .Y(net213423) );
  NOR2X1 U50272 ( .A(n29006), .B(n29005), .Y(n43675) );
  NOR4X1 U50273 ( .A(n29004), .B(n29003), .C(n29002), .D(n29001), .Y(n43674)
         );
  XNOR2X1 U50274 ( .A(n36736), .B(n33762), .Y(net211252) );
  NOR2X1 U50275 ( .A(n19720), .B(n19719), .Y(net211253) );
  NOR4X1 U50276 ( .A(n19718), .B(n19717), .C(n19716), .D(n19715), .Y(net211254) );
  XNOR2X1 U50277 ( .A(n36735), .B(n33842), .Y(n47236) );
  NOR2X1 U50278 ( .A(n19638), .B(n19637), .Y(n47235) );
  NOR4X1 U50279 ( .A(n19636), .B(n19635), .C(n19634), .D(n19633), .Y(n47234)
         );
  NOR4X1 U50280 ( .A(n22329), .B(n22328), .C(n22327), .D(n22326), .Y(n46159)
         );
  XNOR2X1 U50281 ( .A(n33698), .B(n42561), .Y(n44259) );
  NOR2X1 U50282 ( .A(n27111), .B(n27110), .Y(n44258) );
  NOR4X1 U50283 ( .A(n27109), .B(n27108), .C(n27107), .D(n27106), .Y(n44257)
         );
  NAND4X1 U50284 ( .A(n46147), .B(n46146), .C(n46145), .D(n46144), .Y(n12323)
         );
  XNOR2X1 U50285 ( .A(n36840), .B(n33850), .Y(n46146) );
  NOR2X1 U50286 ( .A(n22381), .B(n22380), .Y(n46145) );
  NOR4X1 U50287 ( .A(n22379), .B(n22378), .C(n22377), .D(n22376), .Y(n46144)
         );
  NOR4X1 U50288 ( .A(n22419), .B(n22418), .C(n22417), .D(n22416), .Y(n46114)
         );
  NOR4X1 U50289 ( .A(n22449), .B(n22448), .C(n22447), .D(n22446), .Y(n46099)
         );
  NAND4X1 U50290 ( .A(n43668), .B(n43667), .C(n43666), .D(n43665), .Y(n12064)
         );
  XNOR2X1 U50291 ( .A(n33818), .B(n42569), .Y(n43667) );
  NOR2X1 U50292 ( .A(n29036), .B(n29035), .Y(n43666) );
  NOR4X1 U50293 ( .A(n29034), .B(n29033), .C(n29032), .D(n29031), .Y(n43665)
         );
  NAND4X1 U50294 ( .A(n46157), .B(n46156), .C(n46155), .D(n46154), .Y(n11116)
         );
  XNOR2X1 U50295 ( .A(n36846), .B(n33834), .Y(n46156) );
  NOR2X1 U50296 ( .A(n22341), .B(n22340), .Y(n46155) );
  NOR4X1 U50297 ( .A(n22339), .B(n22338), .C(n22337), .D(n22336), .Y(n46154)
         );
  XNOR2X1 U50298 ( .A(n33850), .B(n42558), .Y(n43553) );
  NOR2X1 U50299 ( .A(n29457), .B(n29456), .Y(n43552) );
  NOR4X1 U50300 ( .A(n29455), .B(n29454), .C(n29453), .D(n29452), .Y(n43551)
         );
  NAND4X1 U50301 ( .A(n45622), .B(n45621), .C(n45620), .D(n45619), .Y(n11205)
         );
  XNOR2X1 U50302 ( .A(n36844), .B(n33738), .Y(n45621) );
  NOR2X1 U50303 ( .A(n24131), .B(n24130), .Y(n45620) );
  NOR4X1 U50304 ( .A(n24129), .B(n24128), .C(n24127), .D(n24126), .Y(n45619)
         );
  XNOR2X1 U50305 ( .A(n36840), .B(n33794), .Y(n47202) );
  NOR2X1 U50306 ( .A(n24050), .B(n24049), .Y(n47201) );
  NOR4X1 U50307 ( .A(n24048), .B(n24047), .C(n24046), .D(n24045), .Y(n47200)
         );
  NAND4X1 U50308 ( .A(n43660), .B(n43659), .C(n43658), .D(n43657), .Y(n12731)
         );
  XNOR2X1 U50309 ( .A(n33834), .B(n42568), .Y(n43659) );
  NOR2X1 U50310 ( .A(n29066), .B(n29065), .Y(n43658) );
  NOR4X1 U50311 ( .A(n29064), .B(n29063), .C(n29062), .D(n29061), .Y(n43657)
         );
  NOR4X1 U50312 ( .A(n20135), .B(n20134), .C(n20133), .D(n20132), .Y(net211481) );
  NAND4X1 U50313 ( .A(n43568), .B(n43567), .C(n43566), .D(n43565), .Y(n12072)
         );
  XNOR2X1 U50314 ( .A(n33866), .B(n42568), .Y(n43567) );
  NOR2X1 U50315 ( .A(n29397), .B(n29396), .Y(n43566) );
  NOR4X1 U50316 ( .A(n29395), .B(n29394), .C(n29393), .D(n29392), .Y(n43565)
         );
  NAND4X1 U50317 ( .A(n47153), .B(n47152), .C(n47151), .D(n47150), .Y(n11417)
         );
  XNOR2X1 U50318 ( .A(n36733), .B(n33826), .Y(n47152) );
  NOR2X1 U50319 ( .A(n19821), .B(n19820), .Y(n47151) );
  NOR4X1 U50320 ( .A(n19819), .B(n19818), .C(n19817), .D(n19816), .Y(n47150)
         );
  XNOR2X1 U50321 ( .A(n36736), .B(n33890), .Y(n47266) );
  NOR4X1 U50322 ( .A(n22349), .B(n22348), .C(n22347), .D(n22346), .Y(n46149)
         );
  NOR4X1 U50323 ( .A(n24099), .B(n24098), .C(n24097), .D(n24096), .Y(n45634)
         );
  XNOR2X1 U50324 ( .A(n33802), .B(n42563), .Y(n44285) );
  NOR2X1 U50325 ( .A(n26780), .B(n26779), .Y(n44284) );
  NOR4X1 U50326 ( .A(n26778), .B(n26777), .C(n26776), .D(n26775), .Y(n44283)
         );
  NAND4X1 U50327 ( .A(n47208), .B(n47207), .C(n47206), .D(n47205), .Y(n11410)
         );
  XNOR2X1 U50328 ( .A(n36736), .B(n33786), .Y(n47207) );
  NOR2X1 U50329 ( .A(n19670), .B(n19669), .Y(n47206) );
  NOR4X1 U50330 ( .A(n19668), .B(n19667), .C(n19666), .D(n19665), .Y(n47205)
         );
  XNOR2X1 U50331 ( .A(n33890), .B(n42568), .Y(n43633) );
  NOR2X1 U50332 ( .A(n29337), .B(n29336), .Y(n43632) );
  NOR4X1 U50333 ( .A(n29335), .B(n29334), .C(n29333), .D(n29332), .Y(n43631)
         );
  NOR4X1 U50334 ( .A(n22369), .B(n22368), .C(n22367), .D(n22366), .Y(n46129)
         );
  XNOR2X1 U50335 ( .A(n36736), .B(n33770), .Y(net211257) );
  NOR2X1 U50336 ( .A(n19731), .B(n19729), .Y(net211258) );
  NOR4X1 U50337 ( .A(n19728), .B(n19727), .C(n19726), .D(n19725), .Y(net211259) );
  XNOR2X1 U50338 ( .A(n36735), .B(n33754), .Y(net211247) );
  NOR2X1 U50339 ( .A(n19710), .B(n19709), .Y(net211248) );
  NOR4X1 U50340 ( .A(n19708), .B(n19707), .C(n19706), .D(n19705), .Y(net211249) );
  NOR2X1 U50341 ( .A(n19648), .B(n19647), .Y(n47230) );
  NOR4X1 U50342 ( .A(n19646), .B(n19645), .C(n19644), .D(n19643), .Y(n47229)
         );
  NAND4X1 U50343 ( .A(n45648), .B(n45647), .C(n45646), .D(n45645), .Y(n12726)
         );
  XNOR2X1 U50344 ( .A(n33786), .B(n42568), .Y(n45647) );
  NOR2X1 U50345 ( .A(n26720), .B(n26719), .Y(n45646) );
  NOR4X1 U50346 ( .A(n26718), .B(n26717), .C(n26716), .D(n26715), .Y(n45645)
         );
  NAND4X1 U50347 ( .A(n46112), .B(n46111), .C(n46110), .D(n46109), .Y(n12329)
         );
  XNOR2X1 U50348 ( .A(n36840), .B(n33882), .Y(n46111) );
  NOR2X1 U50349 ( .A(n22431), .B(n22430), .Y(n46110) );
  NOR4X1 U50350 ( .A(n22429), .B(n22428), .C(n22427), .D(n22426), .Y(n46109)
         );
  NAND4X1 U50351 ( .A(n47213), .B(n47212), .C(n47211), .D(n47210), .Y(n11411)
         );
  XNOR2X1 U50352 ( .A(n36734), .B(n33778), .Y(n47212) );
  NOR2X1 U50353 ( .A(n19660), .B(n19658), .Y(n47211) );
  NOR4X1 U50354 ( .A(n19657), .B(n19656), .C(n19655), .D(n19654), .Y(n47210)
         );
  NAND4X1 U50355 ( .A(n47193), .B(n47192), .C(n47191), .D(n47190), .Y(n12318)
         );
  XNOR2X1 U50356 ( .A(n36845), .B(n33802), .Y(n47192) );
  NOR2X1 U50357 ( .A(n24060), .B(n24059), .Y(n47191) );
  NOR4X1 U50358 ( .A(n24058), .B(n24057), .C(n24056), .D(n24055), .Y(n47190)
         );
  NAND4X1 U50359 ( .A(n45632), .B(n45631), .C(n45630), .D(n45629), .Y(n12311)
         );
  XNOR2X1 U50360 ( .A(n36837), .B(n33722), .Y(n45631) );
  NOR2X1 U50361 ( .A(n24111), .B(n24110), .Y(n45630) );
  NOR4X1 U50362 ( .A(n24109), .B(n24108), .C(n24107), .D(n24106), .Y(n45629)
         );
  NAND4X1 U50363 ( .A(n47257), .B(n47256), .C(n47255), .D(n47254), .Y(n12954)
         );
  XNOR2X1 U50364 ( .A(n36733), .B(n33874), .Y(n47256) );
  NOR2X1 U50365 ( .A(n19558), .B(n19557), .Y(n47255) );
  NOR4X1 U50366 ( .A(n19556), .B(n19555), .C(n19554), .D(n19553), .Y(n47254)
         );
  XNOR2X1 U50367 ( .A(n36841), .B(n33890), .Y(n46121) );
  NOR2X1 U50368 ( .A(n22411), .B(n22410), .Y(n46120) );
  NOR4X1 U50369 ( .A(n22409), .B(n22408), .C(n22407), .D(n22406), .Y(n46119)
         );
  NAND4X1 U50370 ( .A(n44251), .B(n44250), .C(n44249), .D(n44248), .Y(n12717)
         );
  XNOR2X1 U50371 ( .A(n33690), .B(n42561), .Y(n44250) );
  NOR2X1 U50372 ( .A(n27021), .B(n27020), .Y(n44249) );
  NOR4X1 U50373 ( .A(n27019), .B(n27018), .C(n27017), .D(n27016), .Y(n44248)
         );
  NOR4X1 U50374 ( .A(n19829), .B(n19828), .C(n19827), .D(n19826), .Y(n47145)
         );
  NAND4X1 U50375 ( .A(n47198), .B(n47197), .C(n47196), .D(n47195), .Y(n13016)
         );
  XNOR2X1 U50376 ( .A(n36734), .B(n33794), .Y(n47197) );
  NOR2X1 U50377 ( .A(n19680), .B(n19679), .Y(n47196) );
  NOR4X1 U50378 ( .A(n19678), .B(n19677), .C(n19676), .D(n19675), .Y(n47195)
         );
  NAND4X1 U50379 ( .A(n44265), .B(n44264), .C(n44263), .D(n44262), .Y(
        net209817) );
  XNOR2X1 U50380 ( .A(n33706), .B(n42561), .Y(n44264) );
  NOR2X1 U50381 ( .A(n27081), .B(n27080), .Y(n44263) );
  NOR4X1 U50382 ( .A(n27079), .B(n27078), .C(n27077), .D(n27076), .Y(n44262)
         );
  NOR4X1 U50383 ( .A(n19849), .B(n19848), .C(n19847), .D(n19846), .Y(n47135)
         );
  NOR2X1 U50384 ( .A(n29307), .B(n29306), .Y(n43641) );
  NOR4X1 U50385 ( .A(n29305), .B(n29304), .C(n29303), .D(n29302), .Y(n43640)
         );
  NAND4X1 U50386 ( .A(n46137), .B(n46136), .C(n46135), .D(n46134), .Y(n12326)
         );
  XNOR2X1 U50387 ( .A(n36840), .B(n33866), .Y(n46136) );
  NOR2X1 U50388 ( .A(n22361), .B(n22360), .Y(n46135) );
  NOR4X1 U50389 ( .A(n22359), .B(n22358), .C(n22357), .D(n22356), .Y(n46134)
         );
  XNOR2X1 U50390 ( .A(n33778), .B(n36837), .Y(n45652) );
  NOR2X1 U50391 ( .A(n24030), .B(n24029), .Y(n45651) );
  NOR4X1 U50392 ( .A(n24028), .B(n24027), .C(n24026), .D(n24025), .Y(n45650)
         );
  NOR4X1 U50393 ( .A(n43591), .B(n43590), .C(n29186), .D(n29185), .Y(n43592)
         );
  XOR2X1 U50394 ( .A(n33922), .B(n42560), .Y(n43590) );
  XOR2X1 U50395 ( .A(n33924), .B(n36823), .Y(n43591) );
  XOR2X1 U50396 ( .A(n42125), .B(n36877), .Y(n29186) );
  NAND4X1 U50397 ( .A(n47901), .B(n47900), .C(n47899), .D(n47898), .Y(n12959)
         );
  XNOR2X1 U50398 ( .A(n36734), .B(n33906), .Y(n47900) );
  NOR2X1 U50399 ( .A(n19578), .B(n19577), .Y(n47899) );
  NOR4X1 U50400 ( .A(n19576), .B(n19575), .C(n19574), .D(n19573), .Y(n47898)
         );
  XOR2X1 U50401 ( .A(n34036), .B(n36827), .Y(n45686) );
  XOR2X1 U50402 ( .A(n34042), .B(n42558), .Y(n45675) );
  XOR2X1 U50403 ( .A(n34034), .B(n42558), .Y(n45685) );
  NOR4X1 U50404 ( .A(n19789), .B(n19788), .C(n19787), .D(n19786), .Y(n47878)
         );
  NAND4X1 U50405 ( .A(n47906), .B(n47905), .C(n47904), .D(n47903), .Y(n12962)
         );
  XNOR2X1 U50406 ( .A(n36735), .B(n33914), .Y(n47905) );
  NOR2X1 U50407 ( .A(n19588), .B(n19587), .Y(n47904) );
  NOR4X1 U50408 ( .A(n19586), .B(n19585), .C(n19584), .D(n19583), .Y(n47903)
         );
  NAND4X1 U50409 ( .A(n46127), .B(n46126), .C(n46125), .D(n46124), .Y(
        net211197) );
  XNOR2X1 U50410 ( .A(n36843), .B(n33898), .Y(n46126) );
  NOR2X1 U50411 ( .A(n22401), .B(n22400), .Y(n46125) );
  NOR4X1 U50412 ( .A(n22399), .B(n22398), .C(n22397), .D(n22396), .Y(n46124)
         );
  NAND4X1 U50413 ( .A(n45643), .B(n45642), .C(n45641), .D(n45640), .Y(
        net211271) );
  XNOR2X1 U50414 ( .A(n33786), .B(n36846), .Y(n45642) );
  NOR2X1 U50415 ( .A(n24040), .B(n24039), .Y(n45641) );
  NOR4X1 U50416 ( .A(n24038), .B(n24037), .C(n24036), .D(n24035), .Y(n45640)
         );
  NOR4X1 U50417 ( .A(n19546), .B(n19545), .C(n19544), .D(n19543), .Y(n47259)
         );
  XNOR2X1 U50418 ( .A(n36734), .B(n33802), .Y(n47187) );
  NOR2X1 U50419 ( .A(n19690), .B(n19689), .Y(n47186) );
  NOR4X1 U50420 ( .A(n19688), .B(n19687), .C(n19686), .D(n19685), .Y(n47185)
         );
  XNOR2X1 U50421 ( .A(n36764), .B(n33737), .Y(n47162) );
  NOR2X1 U50422 ( .A(n19801), .B(n19800), .Y(n47161) );
  NOR4X1 U50423 ( .A(n19799), .B(n19798), .C(n19797), .D(n19796), .Y(n47160)
         );
  NAND4X1 U50424 ( .A(n47222), .B(n47221), .C(n47220), .D(n47219), .Y(n48057)
         );
  XNOR2X1 U50425 ( .A(n36766), .B(n33857), .Y(n47221) );
  NOR2X1 U50426 ( .A(n19628), .B(n19627), .Y(n47220) );
  NOR4X1 U50427 ( .A(n19626), .B(n19625), .C(n19624), .D(n19623), .Y(n47219)
         );
  XNOR2X1 U50428 ( .A(n36771), .B(n33865), .Y(n47226) );
  NOR2X1 U50429 ( .A(n19618), .B(n19617), .Y(n47225) );
  NAND4X1 U50430 ( .A(n47252), .B(n47251), .C(n47250), .D(n47249), .Y(n12957)
         );
  XNOR2X1 U50431 ( .A(n36735), .B(n33882), .Y(n47251) );
  NOR2X1 U50432 ( .A(n19568), .B(n19567), .Y(n47250) );
  NOR4X1 U50433 ( .A(n19566), .B(n19565), .C(n19564), .D(n19563), .Y(n47249)
         );
  XOR2X1 U50434 ( .A(n33737), .B(n36776), .Y(n45618) );
  XOR2X1 U50435 ( .A(n33764), .B(n36830), .Y(n44308) );
  NOR2X1 U50436 ( .A(n10556), .B(n45654), .Y(net213402) );
  NOR2X1 U50437 ( .A(n12384), .B(n47258), .Y(n47262) );
  XOR2X1 U50438 ( .A(n36774), .B(n33897), .Y(n47258) );
  NOR2X1 U50439 ( .A(n10852), .B(n47159), .Y(n47163) );
  NOR2X1 U50440 ( .A(n11850), .B(n43648), .Y(n43652) );
  NOR2X1 U50441 ( .A(n12385), .B(n47134), .Y(n47138) );
  NOR2X1 U50442 ( .A(n10855), .B(n47214), .Y(net211261) );
  XOR2X1 U50443 ( .A(n36764), .B(n33745), .Y(n47214) );
  NOR2X1 U50444 ( .A(n11741), .B(n44313), .Y(net215213) );
  NOR2X1 U50445 ( .A(n12795), .B(n46148), .Y(n46152) );
  XOR2X1 U50446 ( .A(n36918), .B(n33820), .Y(n46148) );
  NOR2X1 U50447 ( .A(n10424), .B(n44261), .Y(n44265) );
  NOR2X1 U50448 ( .A(n10607), .B(n45633), .Y(n45637) );
  XOR2X1 U50449 ( .A(n41301), .B(n33716), .Y(n45633) );
  NOR2X1 U50450 ( .A(n11204), .B(n47877), .Y(n47881) );
  NOR2X1 U50451 ( .A(n10608), .B(n45623), .Y(n45627) );
  NOR2X1 U50452 ( .A(n11733), .B(n44272), .Y(n44276) );
  XOR2X1 U50453 ( .A(n33716), .B(n36829), .Y(n44272) );
  NOR2X1 U50454 ( .A(n10423), .B(n44266), .Y(net215298) );
  NOR2X1 U50455 ( .A(n11117), .B(n47144), .Y(n47148) );
  NOR2X1 U50456 ( .A(n11744), .B(n45644), .Y(n45648) );
  NOR2X1 U50457 ( .A(n12324), .B(n47223), .Y(n47227) );
  XOR2X1 U50458 ( .A(n33905), .B(n36776), .Y(n46103) );
  NOR2X1 U50459 ( .A(n11752), .B(n43656), .Y(n43660) );
  NAND4X1 U50460 ( .A(n43610), .B(n43609), .C(n37209), .D(n43608), .Y(n43624)
         );
  XNOR2X1 U50461 ( .A(n33906), .B(n42568), .Y(n43609) );
  NOR2X1 U50462 ( .A(n29122), .B(n29133), .Y(n43608) );
  NAND4X1 U50463 ( .A(n43597), .B(n43596), .C(n37254), .D(n43595), .Y(n43607)
         );
  XNOR2X1 U50464 ( .A(n33914), .B(n42568), .Y(n43596) );
  NOR2X1 U50465 ( .A(n29152), .B(n29163), .Y(n43595) );
  NOR2X1 U50466 ( .A(n11848), .B(n43550), .Y(n43554) );
  NOR2X1 U50467 ( .A(n12147), .B(n46138), .Y(n46142) );
  NOR2X1 U50468 ( .A(n12731), .B(n46158), .Y(n46162) );
  NOR2X1 U50469 ( .A(n11114), .B(n47139), .Y(n47143) );
  NOR2X1 U50470 ( .A(n12072), .B(n46128), .Y(n46132) );
  XOR2X1 U50471 ( .A(n33793), .B(n36782), .Y(n47199) );
  XOR2X1 U50472 ( .A(n33820), .B(n36824), .Y(n43664) );
  NOR2X1 U50473 ( .A(n12322), .B(n47228), .Y(n47232) );
  NAND2X1 U50474 ( .A(n44291), .B(n44290), .Y(n44292) );
  XOR2X1 U50475 ( .A(n33796), .B(n36831), .Y(n44289) );
  NOR2X1 U50476 ( .A(n12583), .B(n43639), .Y(n43643) );
  XOR2X1 U50477 ( .A(n36733), .B(n33858), .Y(n47218) );
  NOR2X1 U50478 ( .A(n47042), .B(net209253), .Y(net211483) );
  XOR2X1 U50479 ( .A(n36741), .B(n33964), .Y(n47042) );
  NOR2X1 U50480 ( .A(n46169), .B(net209817), .Y(net212736) );
  XOR2X1 U50481 ( .A(n36772), .B(n33889), .Y(n47263) );
  NOR4X1 U50482 ( .A(n28343), .B(n28342), .C(n28341), .D(n28340), .Y(net215915) );
  NAND4X2 U50483 ( .A(n45782), .B(n45781), .C(n45780), .D(n45779), .Y(n11085)
         );
  XNOR2X1 U50484 ( .A(n36841), .B(n33570), .Y(n45781) );
  NOR2X1 U50485 ( .A(n23463), .B(n23462), .Y(n45780) );
  NOR4X1 U50486 ( .A(n23461), .B(n23460), .C(n23459), .D(n23458), .Y(n45779)
         );
  NOR4X1 U50487 ( .A(n23196), .B(n23195), .C(n23194), .D(n23193), .Y(n45849)
         );
  XNOR2X1 U50488 ( .A(n36846), .B(n33634), .Y(n45751) );
  NOR2X1 U50489 ( .A(n23513), .B(n23512), .Y(n45750) );
  NOR4X1 U50490 ( .A(n23511), .B(n23510), .C(n23509), .D(n23508), .Y(n45749)
         );
  XNOR2X1 U50491 ( .A(n36845), .B(n33490), .Y(n45816) );
  NOR2X1 U50492 ( .A(n23248), .B(n23247), .Y(n45815) );
  NOR4X1 U50493 ( .A(n23246), .B(n23245), .C(n23244), .D(n23243), .Y(n45814)
         );
  XNOR2X1 U50494 ( .A(n36837), .B(n33522), .Y(n45821) );
  NOR2X1 U50495 ( .A(n23238), .B(n23237), .Y(n45820) );
  NOR4X1 U50496 ( .A(n23236), .B(n23235), .C(n23234), .D(n23233), .Y(n45819)
         );
  XNOR2X1 U50497 ( .A(n36839), .B(n33602), .Y(n45731) );
  NOR2X1 U50498 ( .A(n23585), .B(n23583), .Y(n45730) );
  NOR4X1 U50499 ( .A(n23582), .B(n23581), .C(n23580), .D(n23579), .Y(n45729)
         );
  XNOR2X1 U50500 ( .A(n36736), .B(n33650), .Y(net211652) );
  NOR2X1 U50501 ( .A(n21032), .B(n21030), .Y(net211653) );
  NOR4X1 U50502 ( .A(n21029), .B(n21028), .C(n21027), .D(n21026), .Y(net211654) );
  XNOR2X1 U50503 ( .A(n36843), .B(n33506), .Y(n45806) );
  NOR2X1 U50504 ( .A(n23269), .B(n23267), .Y(n45805) );
  NOR4X1 U50505 ( .A(n23266), .B(n23265), .C(n23264), .D(n23263), .Y(n45804)
         );
  XNOR2X1 U50506 ( .A(n33538), .B(n42569), .Y(n43812) );
  NOR2X1 U50507 ( .A(n28105), .B(n28104), .Y(n43811) );
  NOR4X1 U50508 ( .A(n28103), .B(n28102), .C(n28101), .D(n28100), .Y(n43810)
         );
  XNOR2X1 U50509 ( .A(n33410), .B(n36724), .Y(n43226) );
  NOR2X1 U50510 ( .A(n31534), .B(n31533), .Y(n43225) );
  NOR4X1 U50511 ( .A(n31532), .B(n31531), .C(n31530), .D(n31529), .Y(n43224)
         );
  NOR4X1 U50512 ( .A(n22956), .B(n22955), .C(n22954), .D(n22953), .Y(n45916)
         );
  NAND4X2 U50513 ( .A(n44551), .B(n44550), .C(n44549), .D(n44548), .Y(n12035)
         );
  XNOR2X1 U50514 ( .A(n33554), .B(n42559), .Y(n44550) );
  NOR2X1 U50515 ( .A(n24797), .B(n24796), .Y(n44549) );
  NOR4X1 U50516 ( .A(n24795), .B(n24794), .C(n24793), .D(n24792), .Y(n44548)
         );
  XNOR2X1 U50517 ( .A(n33442), .B(n34452), .Y(n43721) );
  NOR2X1 U50518 ( .A(n28435), .B(n28434), .Y(n43720) );
  NOR4X1 U50519 ( .A(n28433), .B(n28432), .C(n28431), .D(n28430), .Y(n43719)
         );
  XNOR2X1 U50520 ( .A(n33426), .B(n34452), .Y(n43739) );
  NOR2X1 U50521 ( .A(n28375), .B(n28374), .Y(n43738) );
  NOR4X1 U50522 ( .A(n28373), .B(n28372), .C(n28371), .D(n28370), .Y(n43737)
         );
  NOR4X1 U50523 ( .A(n25005), .B(n25004), .C(n25003), .D(n25002), .Y(net214882) );
  XNOR2X1 U50524 ( .A(n36845), .B(n33618), .Y(n45761) );
  NOR2X1 U50525 ( .A(n23493), .B(n23492), .Y(n45760) );
  NOR4X1 U50526 ( .A(n23491), .B(n23490), .C(n23489), .D(n23488), .Y(n45759)
         );
  XNOR2X1 U50527 ( .A(n36736), .B(n33522), .Y(n47091) );
  NOR2X1 U50528 ( .A(n19932), .B(n19931), .Y(n47090) );
  NOR4X1 U50529 ( .A(n19930), .B(n19929), .C(n19928), .D(n19927), .Y(n47089)
         );
  XNOR2X1 U50530 ( .A(n33394), .B(n36726), .Y(n43208) );
  NOR2X1 U50531 ( .A(n31594), .B(n31593), .Y(n43207) );
  NOR4X1 U50532 ( .A(n31592), .B(n31591), .C(n31590), .D(n31589), .Y(n43206)
         );
  NAND4X2 U50533 ( .A(n43695), .B(n43694), .C(n43693), .D(n43692), .Y(n12026)
         );
  XNOR2X1 U50534 ( .A(n33490), .B(n42560), .Y(n43694) );
  NOR2X1 U50535 ( .A(n28525), .B(n28524), .Y(n43693) );
  NOR4X1 U50536 ( .A(n28523), .B(n28522), .C(n28521), .D(n28520), .Y(n43692)
         );
  NAND4X1 U50537 ( .A(n46959), .B(n46958), .C(n46957), .D(n46956), .Y(
        net211667) );
  XNOR2X1 U50538 ( .A(n36740), .B(n33676), .Y(n46958) );
  NOR2X1 U50539 ( .A(n21011), .B(n21010), .Y(n46957) );
  NAND4X1 U50540 ( .A(n45757), .B(n45756), .C(n45755), .D(n45754), .Y(n11095)
         );
  XNOR2X1 U50541 ( .A(n36844), .B(n33642), .Y(n45756) );
  NOR2X1 U50542 ( .A(n23503), .B(n23502), .Y(n45755) );
  NOR4X1 U50543 ( .A(n23501), .B(n23500), .C(n23499), .D(n23498), .Y(n45754)
         );
  NAND4X1 U50544 ( .A(n46964), .B(n46963), .C(n46962), .D(n46961), .Y(n12303)
         );
  XNOR2X1 U50545 ( .A(n36837), .B(n33666), .Y(n46963) );
  NOR2X1 U50546 ( .A(n23543), .B(n23542), .Y(n46962) );
  NOR4X1 U50547 ( .A(n23541), .B(n23540), .C(n23539), .D(n23538), .Y(n46961)
         );
  NAND4X1 U50548 ( .A(n44542), .B(n44541), .C(n44540), .D(n44539), .Y(n12034)
         );
  XNOR2X1 U50549 ( .A(n33562), .B(n42558), .Y(n44541) );
  NOR2X1 U50550 ( .A(n24827), .B(n24826), .Y(n44540) );
  NOR4X1 U50551 ( .A(n24825), .B(n24824), .C(n24823), .D(n24822), .Y(n44539)
         );
  XNOR2X1 U50552 ( .A(n36736), .B(n33506), .Y(n47096) );
  NOR2X1 U50553 ( .A(n19922), .B(n19921), .Y(n47095) );
  NOR4X1 U50554 ( .A(n19920), .B(n19919), .C(n19918), .D(n19917), .Y(n47094)
         );
  NOR4X1 U50555 ( .A(n23603), .B(n23602), .C(n23601), .D(n23600), .Y(n45718)
         );
  XNOR2X1 U50556 ( .A(n36841), .B(n33578), .Y(n45776) );
  NOR2X1 U50557 ( .A(n23473), .B(n23472), .Y(n45775) );
  NOR4X1 U50558 ( .A(n23471), .B(n23470), .C(n23469), .D(n23468), .Y(n45774)
         );
  NOR4X1 U50559 ( .A(n23176), .B(n23175), .C(n23174), .D(n23173), .Y(n45839)
         );
  NOR2X1 U50560 ( .A(n28495), .B(n28494), .Y(n43702) );
  NOR4X1 U50561 ( .A(n28493), .B(n28492), .C(n28491), .D(n28490), .Y(n43701)
         );
  NAND4X1 U50562 ( .A(n45857), .B(n45856), .C(n45855), .D(n45854), .Y(n11066)
         );
  XNOR2X1 U50563 ( .A(n36843), .B(n33450), .Y(n45856) );
  NOR2X1 U50564 ( .A(n23188), .B(n23187), .Y(n45855) );
  NOR4X1 U50565 ( .A(n23186), .B(n23185), .C(n23184), .D(n23183), .Y(n45854)
         );
  NAND4X1 U50566 ( .A(n44242), .B(n44241), .C(n44240), .D(n44239), .Y(n12715)
         );
  XNOR2X1 U50567 ( .A(n33682), .B(n42561), .Y(n44241) );
  NOR2X1 U50568 ( .A(n27051), .B(n27050), .Y(n44240) );
  NOR4X1 U50569 ( .A(n27049), .B(n27048), .C(n27047), .D(n27046), .Y(n44239)
         );
  NAND4X1 U50570 ( .A(n43686), .B(n43685), .C(n43684), .D(n43683), .Y(n12025)
         );
  XNOR2X1 U50571 ( .A(n33498), .B(n42569), .Y(n43685) );
  NOR2X1 U50572 ( .A(n28555), .B(n28554), .Y(n43684) );
  NOR4X1 U50573 ( .A(n28553), .B(n28552), .C(n28551), .D(n28550), .Y(n43683)
         );
  XNOR2X1 U50574 ( .A(n36736), .B(n33490), .Y(n47111) );
  NOR2X1 U50575 ( .A(n19892), .B(n19891), .Y(n47110) );
  NOR4X1 U50576 ( .A(n19890), .B(n19889), .C(n19888), .D(n19887), .Y(n47109)
         );
  XNOR2X1 U50577 ( .A(n33666), .B(n42565), .Y(n44483) );
  NOR2X1 U50578 ( .A(n25037), .B(n25036), .Y(n44482) );
  NOR4X1 U50579 ( .A(n25035), .B(n25034), .C(n25033), .D(n25032), .Y(n44481)
         );
  XNOR2X1 U50580 ( .A(n36734), .B(n33634), .Y(n46953) );
  NOR2X1 U50581 ( .A(n20970), .B(n20969), .Y(n46952) );
  NOR4X1 U50582 ( .A(n20968), .B(n20967), .C(n20966), .D(n20965), .Y(n46951)
         );
  NOR4X1 U50583 ( .A(n23226), .B(n23225), .C(n23224), .D(n23223), .Y(n45824)
         );
  NAND4X1 U50584 ( .A(n44569), .B(n44568), .C(n44567), .D(n44566), .Y(n12796)
         );
  XNOR2X1 U50585 ( .A(n33570), .B(n41630), .Y(n44568) );
  NOR2X1 U50586 ( .A(n24737), .B(n24736), .Y(n44567) );
  NOR4X1 U50587 ( .A(n24735), .B(n24734), .C(n24733), .D(n24732), .Y(n44566)
         );
  NOR2X1 U50588 ( .A(n23208), .B(n23207), .Y(n45835) );
  NOR4X1 U50589 ( .A(n23206), .B(n23205), .C(n23204), .D(n23203), .Y(n45834)
         );
  NAND4X1 U50590 ( .A(n45924), .B(n45923), .C(n45922), .D(n45921), .Y(n12280)
         );
  XNOR2X1 U50591 ( .A(n36847), .B(n33402), .Y(n45923) );
  NOR2X1 U50592 ( .A(n22948), .B(n22947), .Y(n45922) );
  NOR4X1 U50593 ( .A(n22946), .B(n22945), .C(n22944), .D(n22943), .Y(n45921)
         );
  NAND4X1 U50594 ( .A(n44475), .B(n44474), .C(n44473), .D(n44472), .Y(n12048)
         );
  XNOR2X1 U50595 ( .A(n33674), .B(n42569), .Y(n44474) );
  NOR2X1 U50596 ( .A(n25067), .B(n25066), .Y(n44473) );
  NOR4X1 U50597 ( .A(n25065), .B(n25064), .C(n25063), .D(n25062), .Y(n44472)
         );
  NOR2X1 U50598 ( .A(n31564), .B(n31563), .Y(n43216) );
  NOR4X1 U50599 ( .A(n31562), .B(n31561), .C(n31560), .D(n31559), .Y(n43215)
         );
  NOR2X1 U50600 ( .A(n23258), .B(n23257), .Y(n45810) );
  NOR4X1 U50601 ( .A(n23256), .B(n23255), .C(n23254), .D(n23253), .Y(n45809)
         );
  XNOR2X1 U50602 ( .A(n33618), .B(n41630), .Y(n44438) );
  NAND4X1 U50603 ( .A(n47178), .B(n47177), .C(n47176), .D(n47175), .Y(n11396)
         );
  XNOR2X1 U50604 ( .A(n36735), .B(n33682), .Y(n47177) );
  NOR2X1 U50605 ( .A(n19751), .B(n19750), .Y(n47176) );
  NOR4X1 U50606 ( .A(n19749), .B(n19748), .C(n19747), .D(n19746), .Y(n47175)
         );
  NOR2X1 U50607 ( .A(n28405), .B(n28404), .Y(n43729) );
  NOR4X1 U50608 ( .A(n28403), .B(n28402), .C(n28401), .D(n28400), .Y(n43728)
         );
  XNOR2X1 U50609 ( .A(n36736), .B(n33666), .Y(net211642) );
  NOR2X1 U50610 ( .A(n21021), .B(n21020), .Y(net211643) );
  NOR4X1 U50611 ( .A(n21019), .B(n21018), .C(n21017), .D(n21016), .Y(net211644) );
  XNOR2X1 U50612 ( .A(n33602), .B(n42569), .Y(n44524) );
  NOR2X1 U50613 ( .A(n24887), .B(n24886), .Y(n44523) );
  NOR4X1 U50614 ( .A(n24885), .B(n24884), .C(n24883), .D(n24882), .Y(n44522)
         );
  NOR2X1 U50615 ( .A(n28465), .B(n28464), .Y(n43711) );
  NOR4X1 U50616 ( .A(n28463), .B(n28462), .C(n28461), .D(n28460), .Y(n43710)
         );
  NOR2X1 U50617 ( .A(n23279), .B(n23278), .Y(n45800) );
  NOR4X1 U50618 ( .A(n23277), .B(n23276), .C(n23275), .D(n23274), .Y(n45799)
         );
  NOR2X1 U50619 ( .A(n23595), .B(n23594), .Y(n45724) );
  NOR4X1 U50620 ( .A(n23593), .B(n23592), .C(n23591), .D(n23590), .Y(n45723)
         );
  NAND4X1 U50621 ( .A(n43795), .B(n43794), .C(n43793), .D(n43792), .Y(n12153)
         );
  XNOR2X1 U50622 ( .A(n33530), .B(n42569), .Y(n43794) );
  NOR2X1 U50623 ( .A(n28165), .B(n28164), .Y(n43793) );
  NOR4X1 U50624 ( .A(n28163), .B(n28162), .C(n28161), .D(n28160), .Y(n43792)
         );
  NAND4X1 U50625 ( .A(n46753), .B(n46752), .C(n46751), .D(n46750), .Y(n12274)
         );
  XNOR2X1 U50626 ( .A(n36837), .B(n33378), .Y(n46752) );
  NOR2X1 U50627 ( .A(n23008), .B(n23007), .Y(n46751) );
  NOR4X1 U50628 ( .A(n23006), .B(n23005), .C(n23004), .D(n23003), .Y(n46750)
         );
  XNOR2X1 U50629 ( .A(n36733), .B(n33658), .Y(net211658) );
  NOR2X1 U50630 ( .A(n21042), .B(n21041), .Y(net211659) );
  NOR4X1 U50631 ( .A(n21040), .B(n21039), .C(n21038), .D(n21037), .Y(net211660) );
  XNOR2X1 U50632 ( .A(n36843), .B(n33418), .Y(n45913) );
  NOR2X1 U50633 ( .A(n22968), .B(n22967), .Y(n45912) );
  NOR4X1 U50634 ( .A(n22966), .B(n22965), .C(n22964), .D(n22963), .Y(n45911)
         );
  NOR2X1 U50635 ( .A(n28135), .B(n28134), .Y(n43802) );
  NOR4X1 U50636 ( .A(n28133), .B(n28132), .C(n28131), .D(n28130), .Y(n43801)
         );
  NAND4X1 U50637 ( .A(n45934), .B(n45933), .C(n45932), .D(n45931), .Y(n11049)
         );
  XNOR2X1 U50638 ( .A(n36838), .B(n33354), .Y(n45933) );
  NOR2X1 U50639 ( .A(n22928), .B(n22927), .Y(n45932) );
  NOR4X1 U50640 ( .A(n22926), .B(n22925), .C(n22924), .D(n22923), .Y(n45931)
         );
  NOR4X1 U50641 ( .A(n22976), .B(n22975), .C(n22974), .D(n22973), .Y(n45906)
         );
  XNOR2X1 U50642 ( .A(n36839), .B(n33466), .Y(net213126) );
  NOR2X1 U50643 ( .A(n23483), .B(n23482), .Y(n45770) );
  NOR4X1 U50644 ( .A(n23481), .B(n23480), .C(n23479), .D(n23478), .Y(n45769)
         );
  XNOR2X1 U50645 ( .A(n33402), .B(n36726), .Y(n43199) );
  NOR2X1 U50646 ( .A(n31624), .B(n31623), .Y(n43198) );
  NOR4X1 U50647 ( .A(n31622), .B(n31621), .C(n31620), .D(n31619), .Y(n43197)
         );
  NOR4X1 U50648 ( .A(n23146), .B(n23145), .C(n23144), .D(n23143), .Y(n45860)
         );
  NAND4X1 U50649 ( .A(n43298), .B(n43297), .C(n43296), .D(n43295), .Y(n12007)
         );
  XNOR2X1 U50650 ( .A(n33362), .B(n42569), .Y(n43297) );
  NOR2X1 U50651 ( .A(n31294), .B(n31293), .Y(n43296) );
  NOR4X1 U50652 ( .A(n31292), .B(n31291), .C(n31290), .D(n31289), .Y(n43295)
         );
  NAND4X1 U50653 ( .A(n47132), .B(n47131), .C(n47130), .D(n47129), .Y(n12287)
         );
  XNOR2X1 U50654 ( .A(n36840), .B(n33474), .Y(n47131) );
  NOR2X1 U50655 ( .A(n23138), .B(n23137), .Y(n47130) );
  NOR4X1 U50656 ( .A(n23136), .B(n23135), .C(n23134), .D(n23133), .Y(n47129)
         );
  XNOR2X1 U50657 ( .A(n36733), .B(n33442), .Y(n47071) );
  NOR2X1 U50658 ( .A(n20003), .B(n20002), .Y(n47070) );
  NOR4X1 U50659 ( .A(n20001), .B(n20000), .C(n19999), .D(n19998), .Y(n47069)
         );
  NOR2X1 U50660 ( .A(n31354), .B(n31353), .Y(n43278) );
  NOR4X1 U50661 ( .A(n31352), .B(n31351), .C(n31350), .D(n31349), .Y(n43277)
         );
  NAND4X1 U50662 ( .A(n43271), .B(n43270), .C(n43269), .D(n43268), .Y(n12799)
         );
  XNOR2X1 U50663 ( .A(n33378), .B(n42569), .Y(n43270) );
  NOR2X1 U50664 ( .A(n31384), .B(n31383), .Y(n43269) );
  NOR4X1 U50665 ( .A(n31382), .B(n31381), .C(n31380), .D(n31379), .Y(n43268)
         );
  NAND4X1 U50666 ( .A(n47087), .B(n47086), .C(n47085), .D(n47084), .Y(n11368)
         );
  XNOR2X1 U50667 ( .A(n36735), .B(n33530), .Y(n47086) );
  NOR2X1 U50668 ( .A(n19942), .B(n19941), .Y(n47085) );
  NOR4X1 U50669 ( .A(n19940), .B(n19939), .C(n19938), .D(n19937), .Y(n47084)
         );
  XNOR2X1 U50670 ( .A(n33626), .B(n42564), .Y(n44430) );
  NOR2X1 U50671 ( .A(n25187), .B(n25186), .Y(n44429) );
  NOR4X1 U50672 ( .A(n25185), .B(n25184), .C(n25183), .D(n25182), .Y(n44428)
         );
  XNOR2X1 U50673 ( .A(n33458), .B(n34452), .Y(n43758) );
  NOR2X1 U50674 ( .A(n28285), .B(n28284), .Y(n43757) );
  NOR4X1 U50675 ( .A(n28283), .B(n28282), .C(n28281), .D(n28280), .Y(n43756)
         );
  NAND4X1 U50676 ( .A(n43307), .B(n43306), .C(n43305), .D(n43304), .Y(n10526)
         );
  XNOR2X1 U50677 ( .A(n33322), .B(n36726), .Y(n43306) );
  NOR2X1 U50678 ( .A(n31264), .B(n31263), .Y(n43305) );
  NOR4X1 U50679 ( .A(n31262), .B(n31261), .C(n31260), .D(n31259), .Y(n43304)
         );
  NAND4X1 U50680 ( .A(n46971), .B(n46970), .C(n46969), .D(n46968), .Y(n12306)
         );
  XNOR2X1 U50681 ( .A(n36841), .B(n33674), .Y(n46970) );
  NOR2X1 U50682 ( .A(n235530), .B(n235520), .Y(n46969) );
  NOR4X1 U50683 ( .A(n235510), .B(n23550), .C(n23549), .D(n23548), .Y(n46968)
         );
  NAND4X1 U50684 ( .A(n47857), .B(n47856), .C(n47855), .D(n47854), .Y(n12929)
         );
  XNOR2X1 U50685 ( .A(n36736), .B(n33586), .Y(n47856) );
  NOR2X1 U50686 ( .A(n21052), .B(n21051), .Y(n47855) );
  NOR4X1 U50687 ( .A(n21050), .B(n21049), .C(n21048), .D(n21047), .Y(n47854)
         );
  NAND4X1 U50688 ( .A(n47102), .B(n47101), .C(n47100), .D(n47099), .Y(n11366)
         );
  XNOR2X1 U50689 ( .A(n36736), .B(n33514), .Y(n47101) );
  NOR2X1 U50690 ( .A(n19912), .B(n19911), .Y(n47100) );
  NOR4X1 U50691 ( .A(n19910), .B(n19909), .C(n19908), .D(n19907), .Y(n47099)
         );
  NAND4X1 U50692 ( .A(n45737), .B(n45736), .C(n45735), .D(n45734), .Y(n12297)
         );
  XNOR2X1 U50693 ( .A(n36839), .B(n33594), .Y(n45736) );
  NOR2X1 U50694 ( .A(n23574), .B(n23572), .Y(n45735) );
  NOR4X1 U50695 ( .A(n23571), .B(n23570), .C(n23569), .D(n23568), .Y(n45734)
         );
  NOR2X1 U50696 ( .A(n21586), .B(n21585), .Y(n46716) );
  NOR4X1 U50697 ( .A(n21584), .B(n21583), .C(n21582), .D(n21581), .Y(n46715)
         );
  NOR4X1 U50698 ( .A(n19960), .B(n19959), .C(n19958), .D(n19957), .Y(n47074)
         );
  NOR2X1 U50699 ( .A(n24767), .B(n24766), .Y(n44558) );
  NOR4X1 U50700 ( .A(n24765), .B(n24764), .C(n24763), .D(n24762), .Y(n44557)
         );
  NAND4X1 U50701 ( .A(n45742), .B(n45741), .C(n45740), .D(n45739), .Y(
        net209225) );
  XNOR2X1 U50702 ( .A(n36838), .B(n33650), .Y(n45741) );
  NOR2X1 U50703 ( .A(n23563), .B(n235620), .Y(n45740) );
  NOR4X1 U50704 ( .A(n235610), .B(n235600), .C(n235590), .D(n235580), .Y(
        n45739) );
  NOR2X1 U50705 ( .A(n19771), .B(n19770), .Y(n47166) );
  NOR4X1 U50706 ( .A(n19769), .B(n19768), .C(n19767), .D(n19766), .Y(n47165)
         );
  NAND4X1 U50707 ( .A(n47127), .B(n47126), .C(n47125), .D(n47124), .Y(n12922)
         );
  XNOR2X1 U50708 ( .A(n36733), .B(n33482), .Y(n47126) );
  NOR2X1 U50709 ( .A(n19862), .B(n19861), .Y(n47125) );
  NOR4X1 U50710 ( .A(n19860), .B(n19859), .C(n19858), .D(n19857), .Y(n47124)
         );
  NAND4X1 U50711 ( .A(n46939), .B(n46938), .C(n46937), .D(n46936), .Y(n11386)
         );
  XNOR2X1 U50712 ( .A(n36733), .B(n33618), .Y(n46938) );
  NOR2X1 U50713 ( .A(n21001), .B(n21000), .Y(n46937) );
  NOR4X1 U50714 ( .A(n20999), .B(n20998), .C(n20997), .D(n20996), .Y(n46936)
         );
  NOR2X1 U50715 ( .A(n24917), .B(n24916), .Y(n44514) );
  NOR4X1 U50716 ( .A(n24915), .B(n24914), .C(n24913), .D(n24912), .Y(n44513)
         );
  NAND4X1 U50717 ( .A(n46768), .B(n46767), .C(n46766), .D(n46765), .Y(n12278)
         );
  XNOR2X1 U50718 ( .A(n36837), .B(n33386), .Y(n46767) );
  NOR2X1 U50719 ( .A(n22998), .B(n22997), .Y(n46766) );
  NOR4X1 U50720 ( .A(n22996), .B(n22995), .C(n22994), .D(n22993), .Y(n46765)
         );
  NAND4X1 U50721 ( .A(n43777), .B(n43776), .C(n43775), .D(n43774), .Y(
        net209960) );
  XNOR2X1 U50722 ( .A(n33514), .B(n42569), .Y(n43776) );
  NOR2X1 U50723 ( .A(n28225), .B(n28224), .Y(n43775) );
  NOR4X1 U50724 ( .A(n28223), .B(n28222), .C(n28221), .D(n28220), .Y(n43774)
         );
  NAND4X1 U50725 ( .A(n45847), .B(n45846), .C(n45845), .D(n45844), .Y(n48521)
         );
  XNOR2X1 U50726 ( .A(n36839), .B(n33434), .Y(n45846) );
  NOR2X1 U50727 ( .A(n23168), .B(n23167), .Y(n45845) );
  NOR4X1 U50728 ( .A(n23166), .B(n23165), .C(n23164), .D(n23163), .Y(n45844)
         );
  NAND4X1 U50729 ( .A(n45899), .B(n45898), .C(n45897), .D(n45896), .Y(n11051)
         );
  XNOR2X1 U50730 ( .A(n36841), .B(n33370), .Y(n45898) );
  NOR2X1 U50731 ( .A(n23018), .B(n23017), .Y(n45897) );
  NOR4X1 U50732 ( .A(n23016), .B(n23015), .C(n23014), .D(n23013), .Y(n45896)
         );
  NAND4X1 U50733 ( .A(n46944), .B(n46943), .C(n46942), .D(n46941), .Y(n11387)
         );
  XNOR2X1 U50734 ( .A(n36735), .B(n33626), .Y(n46943) );
  NOR2X1 U50735 ( .A(n20991), .B(n20990), .Y(n46942) );
  NOR4X1 U50736 ( .A(n20989), .B(n20988), .C(n20987), .D(n20986), .Y(n46941)
         );
  NAND4X1 U50737 ( .A(n46949), .B(n46948), .C(n46947), .D(n46946), .Y(n11388)
         );
  XNOR2X1 U50738 ( .A(n36734), .B(n33642), .Y(n46948) );
  NOR2X1 U50739 ( .A(n20981), .B(n20979), .Y(n46947) );
  NOR4X1 U50740 ( .A(n20978), .B(n20977), .C(n20976), .D(n20975), .Y(n46946)
         );
  NOR2X1 U50741 ( .A(n21102), .B(n21101), .Y(n46917) );
  NOR4X1 U50742 ( .A(n21100), .B(n21099), .C(n21098), .D(n21097), .Y(n46916)
         );
  NOR2X1 U50743 ( .A(n21122), .B(n21121), .Y(n46907) );
  NOR4X1 U50744 ( .A(n21120), .B(n21119), .C(n21118), .D(n21117), .Y(n46906)
         );
  NAND4X1 U50745 ( .A(n47107), .B(n47106), .C(n47105), .D(n47104), .Y(n11510)
         );
  XNOR2X1 U50746 ( .A(n36734), .B(n33498), .Y(n47106) );
  NOR2X1 U50747 ( .A(n19902), .B(n19901), .Y(n47105) );
  NOR4X1 U50748 ( .A(n19900), .B(n19899), .C(n19898), .D(n19897), .Y(n47104)
         );
  NOR2X1 U50749 ( .A(n28315), .B(n28314), .Y(net215905) );
  NOR4X1 U50750 ( .A(n28313), .B(n28312), .C(n28311), .D(n28310), .Y(net215906) );
  NOR4X1 U50751 ( .A(n20011), .B(n20010), .C(n20009), .D(n20008), .Y(n47064)
         );
  NAND4X1 U50752 ( .A(n47057), .B(n47056), .C(n47055), .D(n47054), .Y(n12915)
         );
  XNOR2X1 U50753 ( .A(n36733), .B(n33426), .Y(n47056) );
  NOR2X1 U50754 ( .A(n19993), .B(n19991), .Y(n47055) );
  NOR4X1 U50755 ( .A(n19990), .B(n19989), .C(n19988), .D(n19987), .Y(n47054)
         );
  NAND4X1 U50756 ( .A(n45767), .B(n45766), .C(n45765), .D(n45764), .Y(n11093)
         );
  XNOR2X1 U50757 ( .A(n36838), .B(n33626), .Y(n45766) );
  NOR2X1 U50758 ( .A(n23523), .B(n23522), .Y(n45765) );
  NOR4X1 U50759 ( .A(n23521), .B(n23520), .C(n23519), .D(n23518), .Y(n45764)
         );
  NOR2X1 U50760 ( .A(n28255), .B(n28254), .Y(n43766) );
  NOR4X1 U50761 ( .A(n28253), .B(n28252), .C(n28251), .D(n28250), .Y(n43765)
         );
  NOR2X1 U50762 ( .A(n21506), .B(n21505), .Y(n46761) );
  NOR4X1 U50763 ( .A(n21504), .B(n21503), .C(n21502), .D(n21501), .Y(n46760)
         );
  XOR2X1 U50764 ( .A(n33650), .B(n42560), .Y(n44460) );
  XOR2X1 U50765 ( .A(n33652), .B(n36822), .Y(n44461) );
  XOR2X1 U50766 ( .A(n42159), .B(n36877), .Y(n25096) );
  NAND4X1 U50767 ( .A(n47852), .B(n47851), .C(n47850), .D(n47849), .Y(n12931)
         );
  XNOR2X1 U50768 ( .A(n36734), .B(n33594), .Y(n47851) );
  NOR2X1 U50769 ( .A(n21062), .B(n21061), .Y(n47850) );
  NOR4X1 U50770 ( .A(n21060), .B(n21059), .C(n21058), .D(n21057), .Y(n47849)
         );
  NAND4X1 U50771 ( .A(n47117), .B(n47116), .C(n47115), .D(n47114), .Y(n13017)
         );
  XNOR2X1 U50772 ( .A(n36736), .B(n33474), .Y(n47116) );
  NOR2X1 U50773 ( .A(n19882), .B(n19881), .Y(n47115) );
  NOR4X1 U50774 ( .A(n19880), .B(n19879), .C(n19878), .D(n19877), .Y(n47114)
         );
  NOR2X1 U50775 ( .A(n24857), .B(n24856), .Y(n44531) );
  NOR4X1 U50776 ( .A(n24855), .B(n24854), .C(n24853), .D(n24852), .Y(n44530)
         );
  XNOR2X1 U50777 ( .A(n36839), .B(n33658), .Y(n45746) );
  NOR2X1 U50778 ( .A(n23533), .B(n23532), .Y(n45745) );
  NOR4X1 U50779 ( .A(n23531), .B(n23530), .C(n23529), .D(n23528), .Y(n45744)
         );
  NAND4X1 U50780 ( .A(n46934), .B(n46933), .C(n46932), .D(n46931), .Y(
        net210099) );
  XNOR2X1 U50781 ( .A(n36770), .B(n33601), .Y(n46933) );
  NOR2X1 U50782 ( .A(n21072), .B(n21071), .Y(n46932) );
  NOR4X1 U50783 ( .A(n21070), .B(n21069), .C(n21068), .D(n21067), .Y(n46931)
         );
  NOR2X1 U50784 ( .A(n21607), .B(n21605), .Y(n46706) );
  NOR4X1 U50785 ( .A(n21604), .B(n21603), .C(n21602), .D(n21601), .Y(n46705)
         );
  NOR2X1 U50786 ( .A(n21082), .B(n21081), .Y(n46927) );
  NOR4X1 U50787 ( .A(n21080), .B(n21079), .C(n21078), .D(n21077), .Y(n46926)
         );
  NOR2X1 U50788 ( .A(n19741), .B(n19740), .Y(n47181) );
  NOR4X1 U50789 ( .A(n19739), .B(n19738), .C(n19737), .D(n19736), .Y(n47180)
         );
  NAND4X1 U50790 ( .A(n46783), .B(n46782), .C(n46781), .D(n46780), .Y(
        net210091) );
  XNOR2X1 U50791 ( .A(n36766), .B(n33345), .Y(n46782) );
  NOR2X1 U50792 ( .A(n21456), .B(n21455), .Y(n46781) );
  NOR4X1 U50793 ( .A(n21454), .B(n21453), .C(n21452), .D(n21451), .Y(n46780)
         );
  NOR4X1 U50794 ( .A(n19980), .B(n19979), .C(n19978), .D(n19977), .Y(n47059)
         );
  NOR2X1 U50795 ( .A(n11711), .B(n44503), .Y(n44507) );
  XOR2X1 U50796 ( .A(n33588), .B(n36822), .Y(n44503) );
  NOR2X1 U50797 ( .A(n11085), .B(n46905), .Y(n46909) );
  NOR2X1 U50798 ( .A(n11699), .B(n43782), .Y(n43786) );
  NOR2X1 U50799 ( .A(n12501), .B(n43691), .Y(n43695) );
  NOR2X1 U50800 ( .A(n11065), .B(n47058), .Y(n47062) );
  NOR2X1 U50801 ( .A(n11693), .B(n43745), .Y(net215912) );
  XOR2X1 U50802 ( .A(n33476), .B(n36825), .Y(n43745) );
  NOR2X1 U50803 ( .A(n11706), .B(n43809), .Y(n43813) );
  NOR2X1 U50804 ( .A(n11208), .B(n47848), .Y(n47852) );
  NOR2X1 U50805 ( .A(n12506), .B(n44547), .Y(n44551) );
  XOR2X1 U50806 ( .A(n33529), .B(n36779), .Y(n45833) );
  NOR2X1 U50807 ( .A(n11058), .B(n46714), .Y(n46718) );
  XOR2X1 U50808 ( .A(n33401), .B(n36786), .Y(n45920) );
  NOR2X1 U50809 ( .A(n12035), .B(n45823), .Y(n45827) );
  NOR2X1 U50810 ( .A(n10847), .B(n47164), .Y(n47168) );
  NOR2X1 U50811 ( .A(n11697), .B(n43700), .Y(n43704) );
  XOR2X1 U50812 ( .A(n33308), .B(n36831), .Y(n43330) );
  NOR2X1 U50813 ( .A(n11092), .B(n46925), .Y(n46929) );
  NOR2X1 U50814 ( .A(n12026), .B(n45864), .Y(net213115) );
  NOR2X1 U50815 ( .A(n11694), .B(n43750), .Y(net215903) );
  NOR2X1 U50816 ( .A(n11095), .B(n46950), .Y(n46954) );
  NOR2X1 U50817 ( .A(n12034), .B(n45768), .Y(n45772) );
  NOR2X1 U50818 ( .A(n12387), .B(n46915), .Y(n46919) );
  NOR2X1 U50819 ( .A(n11686), .B(n43727), .Y(n43731) );
  NOR2X1 U50820 ( .A(n11705), .B(n43791), .Y(n43795) );
  XOR2X1 U50821 ( .A(n33532), .B(n36821), .Y(n43791) );
  NOR2X1 U50822 ( .A(n11698), .B(n43682), .Y(n43686) );
  XOR2X1 U50823 ( .A(n33500), .B(n36824), .Y(n43682) );
  NOR2X1 U50824 ( .A(n12797), .B(n45808), .Y(n45812) );
  NOR2X1 U50825 ( .A(n12715), .B(n46967), .Y(n46971) );
  XOR2X1 U50826 ( .A(n36918), .B(n33676), .Y(n46967) );
  NOR2X1 U50827 ( .A(n11687), .B(n43709), .Y(n43713) );
  NOR2X1 U50828 ( .A(n11211), .B(n47078), .Y(n47082) );
  XOR2X1 U50829 ( .A(n36767), .B(n33537), .Y(n47078) );
  NOR2X1 U50830 ( .A(n12049), .B(n45743), .Y(n45747) );
  NOR2X1 U50831 ( .A(n12796), .B(n45783), .Y(n45787) );
  XOR2X1 U50832 ( .A(n41305), .B(n33564), .Y(n45783) );
  NOR2X1 U50833 ( .A(n12154), .B(n45798), .Y(n45802) );
  NOR2X1 U50834 ( .A(n40392), .B(n46960), .Y(n46964) );
  XOR2X1 U50835 ( .A(n33665), .B(n36779), .Y(n46960) );
  NOR2X1 U50836 ( .A(n12014), .B(n45915), .Y(n45919) );
  NOR2X1 U50837 ( .A(n12016), .B(n45838), .Y(n45842) );
  NOR2X1 U50838 ( .A(n11717), .B(n44512), .Y(n44516) );
  NOR2X1 U50839 ( .A(n11709), .B(n44538), .Y(n44542) );
  XOR2X1 U50840 ( .A(n36735), .B(n33602), .Y(n46930) );
  NOR2X1 U50841 ( .A(n12692), .B(n45848), .Y(n45852) );
  NOR2X1 U50842 ( .A(n11712), .B(n44556), .Y(n44560) );
  NOR2X1 U50843 ( .A(n11721), .B(n44427), .Y(n44431) );
  XOR2X1 U50844 ( .A(n33636), .B(n36821), .Y(n44489) );
  NOR2X1 U50845 ( .A(n11083), .B(n46910), .Y(n46914) );
  XOR2X1 U50846 ( .A(n36741), .B(n33556), .Y(n46910) );
  NOR2X1 U50847 ( .A(n11049), .B(n46779), .Y(n46783) );
  XOR2X1 U50848 ( .A(n36736), .B(n33346), .Y(n46779) );
  NOR2X1 U50849 ( .A(n11054), .B(n46759), .Y(n46763) );
  NOR2X1 U50850 ( .A(n12386), .B(n47179), .Y(n47183) );
  XOR2X1 U50851 ( .A(n33537), .B(n36778), .Y(n45828) );
  NOR2X1 U50852 ( .A(n10827), .B(n47118), .Y(n47122) );
  XOR2X1 U50853 ( .A(n36741), .B(n33460), .Y(n47118) );
  NOR2X1 U50854 ( .A(n11082), .B(n47073), .Y(n47077) );
  NOR2X1 U50855 ( .A(n10157), .B(n45945), .Y(n45949) );
  XOR2X1 U50856 ( .A(n41305), .B(n33300), .Y(n45945) );
  NOR2X1 U50857 ( .A(n12157), .B(n45905), .Y(n45909) );
  XOR2X1 U50858 ( .A(n33393), .B(n36784), .Y(n45905) );
  NOR2X1 U50859 ( .A(n12686), .B(n46749), .Y(n46753) );
  NOR2X1 U50860 ( .A(n46704), .B(n48522), .Y(n46708) );
  NOR2X1 U50861 ( .A(n12490), .B(n43196), .Y(n43200) );
  XOR2X1 U50862 ( .A(n33404), .B(n36825), .Y(n43196) );
  NOR2X1 U50863 ( .A(n12587), .B(n43764), .Y(n43768) );
  XOR2X1 U50864 ( .A(n33412), .B(n36821), .Y(n43223) );
  NOR2X1 U50865 ( .A(n12585), .B(n44529), .Y(n44533) );
  XOR2X1 U50866 ( .A(n33612), .B(n36824), .Y(n44529) );
  NOR2X1 U50867 ( .A(n47063), .B(net209202), .Y(n47067) );
  NOR2X1 U50868 ( .A(n12586), .B(n43800), .Y(n43804) );
  XOR2X1 U50869 ( .A(n33548), .B(n36823), .Y(n43800) );
  NOR2X1 U50870 ( .A(n12706), .B(n45717), .Y(n45721) );
  NOR2X1 U50871 ( .A(n12518), .B(n44480), .Y(n44484) );
  NOR2X1 U50872 ( .A(n10530), .B(n45859), .Y(n45863) );
  NOR2X1 U50873 ( .A(n44435), .B(net209503), .Y(n44439) );
  XOR2X1 U50874 ( .A(n33620), .B(n36831), .Y(n44435) );
  NOR2X1 U50875 ( .A(n43214), .B(n48387), .Y(n43218) );
  NOR2X1 U50876 ( .A(n44471), .B(n44598), .Y(n44475) );
  XOR2X1 U50877 ( .A(n33676), .B(n36822), .Y(n44471) );
  NOR2X1 U50878 ( .A(n43276), .B(net214730), .Y(n43280) );
  XNOR2X1 U50879 ( .A(n36843), .B(n33306), .Y(net213023) );
  XNOR2X1 U50880 ( .A(n36843), .B(n33322), .Y(net213017) );
  XNOR2X1 U50881 ( .A(n36845), .B(n33274), .Y(net212982) );
  NOR2X1 U50882 ( .A(n22867), .B(n22866), .Y(net212983) );
  NOR4X1 U50883 ( .A(n22865), .B(n22864), .C(n22863), .D(n22862), .Y(net212984) );
  NOR4X1 U50884 ( .A(n31863), .B(n31862), .C(n31861), .D(n31860), .Y(net214649) );
  NOR4X1 U50885 ( .A(n19970), .B(n19969), .C(n19968), .D(n19967), .Y(net211351) );
  NOR2X1 U50886 ( .A(n31835), .B(n31834), .Y(net214643) );
  NOR4X1 U50887 ( .A(n31833), .B(n31832), .C(n31831), .D(n31830), .Y(net214644) );
  NAND4X1 U50888 ( .A(n43391), .B(n43390), .C(n43389), .D(n43388), .Y(n11984)
         );
  XNOR2X1 U50889 ( .A(n33178), .B(n42569), .Y(n43390) );
  NOR2X1 U50890 ( .A(n30963), .B(n30962), .Y(n43389) );
  NOR4X1 U50891 ( .A(n30961), .B(n30960), .C(n30959), .D(n30958), .Y(n43388)
         );
  NOR4X1 U50892 ( .A(n21747), .B(n21746), .C(n21745), .D(n21744), .Y(net211990) );
  NAND4X1 U50893 ( .A(n43347), .B(n43346), .C(n43345), .D(n43344), .Y(n11991)
         );
  XNOR2X1 U50894 ( .A(n33218), .B(n42569), .Y(n43346) );
  NOR2X1 U50895 ( .A(n31113), .B(n31112), .Y(n43345) );
  NOR4X1 U50896 ( .A(n31111), .B(n31110), .C(n31109), .D(n31108), .Y(n43344)
         );
  NAND4X1 U50897 ( .A(n45884), .B(n45883), .C(n45882), .D(n45881), .Y(n11031)
         );
  XNOR2X1 U50898 ( .A(n36841), .B(n33218), .Y(n45883) );
  NOR2X1 U50899 ( .A(n23068), .B(n23067), .Y(n45882) );
  NOR4X1 U50900 ( .A(n23066), .B(n23065), .C(n23064), .D(n23063), .Y(n45881)
         );
  NAND4X1 U50901 ( .A(n45978), .B(n45977), .C(n45976), .D(n45975), .Y(n11035)
         );
  XNOR2X1 U50902 ( .A(n36844), .B(n33266), .Y(n45977) );
  NOR2X1 U50903 ( .A(n22806), .B(n22805), .Y(n45976) );
  NOR4X1 U50904 ( .A(n22804), .B(n22803), .C(n22802), .D(n22801), .Y(n45975)
         );
  NAND4X1 U50905 ( .A(n45973), .B(n45972), .C(n45971), .D(n45970), .Y(n11040)
         );
  XNOR2X1 U50906 ( .A(n36843), .B(n33282), .Y(n45972) );
  NOR2X1 U50907 ( .A(n22816), .B(n22815), .Y(n45971) );
  NOR4X1 U50908 ( .A(n22814), .B(n22813), .C(n22812), .D(n22811), .Y(n45970)
         );
  NAND4X1 U50909 ( .A(n43316), .B(n43315), .C(n43314), .D(n43313), .Y(n10525)
         );
  XNOR2X1 U50910 ( .A(n33314), .B(n42569), .Y(n43315) );
  NOR2X1 U50911 ( .A(n31234), .B(n31233), .Y(n43314) );
  NOR4X1 U50912 ( .A(n31232), .B(n31231), .C(n31230), .D(n31229), .Y(n43313)
         );
  NAND4X1 U50913 ( .A(n45944), .B(n45943), .C(n45942), .D(n45941), .Y(n12270)
         );
  XNOR2X1 U50914 ( .A(n36840), .B(n33338), .Y(n45943) );
  NOR2X1 U50915 ( .A(n22908), .B(n22907), .Y(n45942) );
  NOR4X1 U50916 ( .A(n22906), .B(n22905), .C(n22904), .D(n22903), .Y(n45941)
         );
  NAND4X1 U50917 ( .A(n43356), .B(n43355), .C(n43354), .D(n43353), .Y(n11988)
         );
  XNOR2X1 U50918 ( .A(n33210), .B(n42569), .Y(n43355) );
  NOR2X1 U50919 ( .A(n31083), .B(n31082), .Y(n43354) );
  NOR4X1 U50920 ( .A(n31081), .B(n31080), .C(n31079), .D(n31078), .Y(n43353)
         );
  NAND4X1 U50921 ( .A(n45889), .B(n45888), .C(n45887), .D(n45886), .Y(n11028)
         );
  XNOR2X1 U50922 ( .A(n36847), .B(n33210), .Y(n45888) );
  NOR2X1 U50923 ( .A(n23058), .B(n23057), .Y(n45887) );
  NOR4X1 U50924 ( .A(n23056), .B(n23055), .C(n23054), .D(n23053), .Y(n45886)
         );
  NOR4X1 U50925 ( .A(n21767), .B(n21766), .C(n21765), .D(n21764), .Y(net212000) );
  NAND4X1 U50926 ( .A(n45983), .B(n45982), .C(n45981), .D(n45980), .Y(n12262)
         );
  XNOR2X1 U50927 ( .A(n36847), .B(n33242), .Y(n45982) );
  NOR2X1 U50928 ( .A(n22877), .B(n22876), .Y(n45981) );
  NOR4X1 U50929 ( .A(n22875), .B(n22874), .C(n22873), .D(n22872), .Y(n45980)
         );
  NOR4X1 U50930 ( .A(n22916), .B(n22915), .C(n22914), .D(n22913), .Y(n45936)
         );
  NAND4X1 U50931 ( .A(n44635), .B(n44634), .C(n44633), .D(n44632), .Y(n11994)
         );
  XNOR2X1 U50932 ( .A(n33234), .B(n42560), .Y(n44634) );
  NOR2X1 U50933 ( .A(n31805), .B(n31804), .Y(n44633) );
  NOR4X1 U50934 ( .A(n31803), .B(n31802), .C(n31801), .D(n31800), .Y(n44632)
         );
  NAND4X1 U50935 ( .A(n43382), .B(n43381), .C(n43380), .D(n43379), .Y(n12800)
         );
  XNOR2X1 U50936 ( .A(n33186), .B(n42569), .Y(n43381) );
  NOR2X1 U50937 ( .A(n30993), .B(n30992), .Y(n43380) );
  NOR4X1 U50938 ( .A(n30991), .B(n30990), .C(n30989), .D(n30988), .Y(n43379)
         );
  NAND4X1 U50939 ( .A(n45929), .B(n45928), .C(n45927), .D(n45926), .Y(n12389)
         );
  XNOR2X1 U50940 ( .A(n36844), .B(n33330), .Y(n45928) );
  NOR2X1 U50941 ( .A(n22938), .B(n22937), .Y(n45927) );
  NOR4X1 U50942 ( .A(n22936), .B(n22935), .C(n22934), .D(n22933), .Y(n45926)
         );
  NAND4X1 U50943 ( .A(n43339), .B(n43338), .C(n43337), .D(n43336), .Y(n11990)
         );
  XNOR2X1 U50944 ( .A(n33226), .B(n42569), .Y(n43338) );
  NOR2X1 U50945 ( .A(n31143), .B(n31142), .Y(n43337) );
  NOR4X1 U50946 ( .A(n31141), .B(n31140), .C(n31139), .D(n31138), .Y(n43336)
         );
  NAND4X1 U50947 ( .A(n45879), .B(n45878), .C(n45877), .D(n45876), .Y(n11030)
         );
  XNOR2X1 U50948 ( .A(n36839), .B(n33226), .Y(n45878) );
  NOR2X1 U50949 ( .A(n23078), .B(n23077), .Y(n45877) );
  NOR4X1 U50950 ( .A(n23076), .B(n23075), .C(n23074), .D(n23073), .Y(n45876)
         );
  NAND4X1 U50951 ( .A(n45968), .B(n45967), .C(n45966), .D(n45965), .Y(n11039)
         );
  XNOR2X1 U50952 ( .A(n36845), .B(n33290), .Y(n45967) );
  NOR2X1 U50953 ( .A(n22826), .B(n22825), .Y(n45966) );
  NOR4X1 U50954 ( .A(n22824), .B(n22823), .C(n22822), .D(n22821), .Y(n45965)
         );
  NOR2X1 U50955 ( .A(n31324), .B(n31323), .Y(n43287) );
  NOR4X1 U50956 ( .A(n31322), .B(n31321), .C(n31320), .D(n31319), .Y(n43286)
         );
  NAND4X1 U50957 ( .A(n45874), .B(n45873), .C(n45872), .D(n45871), .Y(n11024)
         );
  XNOR2X1 U50958 ( .A(n36839), .B(n33186), .Y(n45873) );
  NOR2X1 U50959 ( .A(n23108), .B(n23107), .Y(n45872) );
  NOR4X1 U50960 ( .A(n23106), .B(n23105), .C(n23104), .D(n23103), .Y(n45871)
         );
  NAND4X1 U50961 ( .A(n43364), .B(n43363), .C(n43362), .D(n43361), .Y(n11989)
         );
  XNOR2X1 U50962 ( .A(n33202), .B(n42569), .Y(n43363) );
  NOR2X1 U50963 ( .A(n31053), .B(n31052), .Y(n43362) );
  NOR4X1 U50964 ( .A(n31051), .B(n31050), .C(n31049), .D(n31048), .Y(n43361)
         );
  NAND4X1 U50965 ( .A(n45894), .B(n45893), .C(n45892), .D(n45891), .Y(n11029)
         );
  XNOR2X1 U50966 ( .A(n36837), .B(n33202), .Y(n45893) );
  NOR2X1 U50967 ( .A(n23048), .B(n23047), .Y(n45892) );
  NOR4X1 U50968 ( .A(n23046), .B(n23045), .C(n23044), .D(n23043), .Y(n45891)
         );
  XNOR2X1 U50969 ( .A(n33346), .B(n42569), .Y(n43262) );
  NOR2X1 U50970 ( .A(n31414), .B(n31413), .Y(n43261) );
  NOR4X1 U50971 ( .A(n31412), .B(n31411), .C(n31410), .D(n31409), .Y(n43260)
         );
  NOR4X1 U50972 ( .A(n21697), .B(n21696), .C(n21695), .D(n21694), .Y(net212005) );
  NAND4X1 U50973 ( .A(n46879), .B(n46878), .C(n46877), .D(n46876), .Y(n12255)
         );
  XNOR2X1 U50974 ( .A(n36844), .B(n33178), .Y(n46878) );
  NOR2X1 U50975 ( .A(n23098), .B(n23097), .Y(n46877) );
  NOR4X1 U50976 ( .A(n23096), .B(n23095), .C(n23094), .D(n23093), .Y(n46876)
         );
  NAND4X1 U50977 ( .A(n43325), .B(n43324), .C(n43323), .D(n43322), .Y(n10527)
         );
  XNOR2X1 U50978 ( .A(n33298), .B(n42569), .Y(n43324) );
  NOR2X1 U50979 ( .A(n31204), .B(n31203), .Y(n43323) );
  NOR4X1 U50980 ( .A(n31202), .B(n31201), .C(n31200), .D(n31199), .Y(n43322)
         );
  NAND4X1 U50981 ( .A(n43186), .B(n43185), .C(n43184), .D(n43183), .Y(n12668)
         );
  XNOR2X1 U50982 ( .A(n33250), .B(n36725), .Y(n43185) );
  NOR2X1 U50983 ( .A(n31655), .B(n31654), .Y(n43184) );
  NOR4X1 U50984 ( .A(n31653), .B(n31652), .C(n31651), .D(n31650), .Y(n43183)
         );
  NAND4X1 U50985 ( .A(n45963), .B(n45962), .C(n45961), .D(n45960), .Y(n12260)
         );
  XNOR2X1 U50986 ( .A(n36838), .B(n33250), .Y(n45962) );
  NOR2X1 U50987 ( .A(n22836), .B(n22835), .Y(n45961) );
  NOR4X1 U50988 ( .A(n22834), .B(n22833), .C(n22832), .D(n22831), .Y(n45960)
         );
  NAND4X1 U50989 ( .A(n43172), .B(n43171), .C(n43170), .D(n43169), .Y(n12672)
         );
  XNOR2X1 U50990 ( .A(n33282), .B(n36725), .Y(n43171) );
  NOR2X1 U50991 ( .A(n31745), .B(n31744), .Y(n43170) );
  NOR4X1 U50992 ( .A(n31743), .B(n31742), .C(n31741), .D(n31740), .Y(n43169)
         );
  XNOR2X1 U50993 ( .A(n36774), .B(n33353), .Y(n46777) );
  NOR2X1 U50994 ( .A(n21466), .B(n21465), .Y(n46776) );
  XNOR2X1 U50995 ( .A(n36734), .B(n33282), .Y(net211993) );
  NOR2X1 U50996 ( .A(n21759), .B(n21758), .Y(net211994) );
  NOR4X1 U50997 ( .A(n21757), .B(n21756), .C(n21755), .D(n21754), .Y(net211995) );
  NAND4X1 U50998 ( .A(n43373), .B(n43372), .C(n43371), .D(n43370), .Y(n12665)
         );
  XNOR2X1 U50999 ( .A(n33194), .B(n42569), .Y(n43372) );
  NOR2X1 U51000 ( .A(n31023), .B(n31022), .Y(n43371) );
  NOR4X1 U51001 ( .A(n31021), .B(n31020), .C(n31019), .D(n31018), .Y(n43370)
         );
  NAND4X1 U51002 ( .A(n43236), .B(n43235), .C(n43234), .D(n43233), .Y(
        net209778) );
  XNOR2X1 U51003 ( .A(n33338), .B(n36726), .Y(n43235) );
  NOR2X1 U51004 ( .A(n31504), .B(n31503), .Y(n43234) );
  NOR4X1 U51005 ( .A(n31502), .B(n31501), .C(n31500), .D(n31499), .Y(n43233)
         );
  NAND4X1 U51006 ( .A(n43191), .B(n43190), .C(n43189), .D(n43188), .Y(
        net209767) );
  XNOR2X1 U51007 ( .A(n33242), .B(n36725), .Y(n43190) );
  NOR2X1 U51008 ( .A(n31715), .B(n31714), .Y(n43189) );
  NOR4X1 U51009 ( .A(n31713), .B(n31712), .C(n31711), .D(n31710), .Y(n43188)
         );
  NAND4X1 U51010 ( .A(n46798), .B(n46797), .C(n46796), .D(n46795), .Y(n12251)
         );
  XNOR2X1 U51011 ( .A(n36846), .B(n33170), .Y(n46797) );
  NOR2X1 U51012 ( .A(n23088), .B(n23087), .Y(n46796) );
  NOR4X1 U51013 ( .A(n23086), .B(n23085), .C(n23084), .D(n23083), .Y(n46795)
         );
  NAND4X1 U51014 ( .A(n45869), .B(n45868), .C(n45867), .D(n45866), .Y(n11023)
         );
  XNOR2X1 U51015 ( .A(n36838), .B(n33194), .Y(n45868) );
  NOR2X1 U51016 ( .A(n23118), .B(n23117), .Y(n45867) );
  NOR4X1 U51017 ( .A(n23116), .B(n23115), .C(n23114), .D(n23113), .Y(n45866)
         );
  NAND4X1 U51018 ( .A(n43163), .B(n43162), .C(n43161), .D(n43160), .Y(n12675)
         );
  XNOR2X1 U51019 ( .A(n33290), .B(n36726), .Y(n43162) );
  NOR2X1 U51020 ( .A(n31775), .B(n31774), .Y(n43161) );
  NOR4X1 U51021 ( .A(n31773), .B(n31772), .C(n31771), .D(n31770), .Y(n43160)
         );
  NAND4X1 U51022 ( .A(n43181), .B(n43180), .C(n43179), .D(n43178), .Y(n12671)
         );
  XNOR2X1 U51023 ( .A(n33258), .B(n36726), .Y(n43180) );
  NOR2X1 U51024 ( .A(n31685), .B(n31684), .Y(n43179) );
  NOR4X1 U51025 ( .A(n31683), .B(n31682), .C(n31681), .D(n31680), .Y(n43178)
         );
  NAND4X1 U51026 ( .A(n45958), .B(n45957), .C(n45956), .D(n45955), .Y(n12264)
         );
  XNOR2X1 U51027 ( .A(n36837), .B(n33258), .Y(n45957) );
  NOR2X1 U51028 ( .A(n22846), .B(n22845), .Y(n45956) );
  NOR4X1 U51029 ( .A(n22844), .B(n22843), .C(n22842), .D(n22841), .Y(n45955)
         );
  NOR2X1 U51030 ( .A(n21203), .B(n21202), .Y(n46862) );
  NOR4X1 U51031 ( .A(n21201), .B(n21200), .C(n21199), .D(n21198), .Y(n46861)
         );
  NAND4X1 U51032 ( .A(n45904), .B(n45903), .C(n45902), .D(n45901), .Y(n11052)
         );
  XNOR2X1 U51033 ( .A(n36847), .B(n33362), .Y(n45903) );
  NOR2X1 U51034 ( .A(n22988), .B(n22987), .Y(n45902) );
  NOR4X1 U51035 ( .A(n22986), .B(n22985), .C(n22984), .D(n22983), .Y(n45901)
         );
  NAND4X1 U51036 ( .A(n46884), .B(n46883), .C(n46882), .D(n46881), .Y(n11515)
         );
  XNOR2X1 U51037 ( .A(n36736), .B(n33170), .Y(n46883) );
  NOR2X1 U51038 ( .A(n21173), .B(n21172), .Y(n46882) );
  NOR4X1 U51039 ( .A(n21171), .B(n21170), .C(n21169), .D(n21168), .Y(n46881)
         );
  NOR2X1 U51040 ( .A(n21516), .B(n21515), .Y(n46756) );
  NOR4X1 U51041 ( .A(n21514), .B(n21513), .C(n21512), .D(n21511), .Y(n46755)
         );
  XNOR2X1 U51042 ( .A(n33354), .B(n42558), .Y(n43253) );
  NOR2X1 U51043 ( .A(n31444), .B(n31443), .Y(n43252) );
  NOR4X1 U51044 ( .A(n31442), .B(n31441), .C(n31440), .D(n31439), .Y(n43251)
         );
  XNOR2X1 U51045 ( .A(n36733), .B(n33202), .Y(n46893) );
  NOR2X1 U51046 ( .A(n21153), .B(n21152), .Y(n46892) );
  NOR4X1 U51047 ( .A(n21151), .B(n21150), .C(n21149), .D(n21148), .Y(n46891)
         );
  NAND4X1 U51048 ( .A(n46869), .B(n46868), .C(n46867), .D(n46866), .Y(n11325)
         );
  XNOR2X1 U51049 ( .A(n36735), .B(n33186), .Y(n46868) );
  NOR2X1 U51050 ( .A(n21193), .B(n21192), .Y(n46867) );
  NOR4X1 U51051 ( .A(n21191), .B(n21190), .C(n21189), .D(n21188), .Y(n46866)
         );
  NAND4X1 U51052 ( .A(n46679), .B(n46678), .C(n46677), .D(n46676), .Y(n11334)
         );
  XNOR2X1 U51053 ( .A(n36736), .B(n33258), .Y(n46678) );
  NOR2X1 U51054 ( .A(n21719), .B(n21718), .Y(n46677) );
  NOR4X1 U51055 ( .A(n21717), .B(n21716), .C(n21715), .D(n21714), .Y(n46676)
         );
  NAND4X1 U51056 ( .A(n46899), .B(n46898), .C(n46897), .D(n46896), .Y(n12893)
         );
  XNOR2X1 U51057 ( .A(n36734), .B(n33226), .Y(n46898) );
  NOR2X1 U51058 ( .A(n21143), .B(n21142), .Y(n46897) );
  NOR4X1 U51059 ( .A(n21141), .B(n21140), .C(n21139), .D(n21138), .Y(n46896)
         );
  NAND4X1 U51060 ( .A(n46889), .B(n46888), .C(n46887), .D(n46886), .Y(n11326)
         );
  XNOR2X1 U51061 ( .A(n36735), .B(n33210), .Y(n46888) );
  NOR2X1 U51062 ( .A(n21163), .B(n21162), .Y(n46887) );
  NOR4X1 U51063 ( .A(n21161), .B(n21160), .C(n21159), .D(n21158), .Y(n46886)
         );
  NOR2X1 U51064 ( .A(n21486), .B(n21485), .Y(n47924) );
  NOR4X1 U51065 ( .A(n21484), .B(n21483), .C(n21482), .D(n21481), .Y(n47923)
         );
  NAND4X1 U51066 ( .A(n47921), .B(n47920), .C(n47919), .D(n47918), .Y(n12906)
         );
  XNOR2X1 U51067 ( .A(n36736), .B(n33330), .Y(n47920) );
  NOR2X1 U51068 ( .A(n21476), .B(n21475), .Y(n47919) );
  NOR4X1 U51069 ( .A(n21474), .B(n21473), .C(n21472), .D(n21471), .Y(n47918)
         );
  NAND4X1 U51070 ( .A(n47931), .B(n47930), .C(n47929), .D(n47928), .Y(n12892)
         );
  XNOR2X1 U51071 ( .A(n36733), .B(n33234), .Y(n47930) );
  NOR2X1 U51072 ( .A(n21739), .B(n21738), .Y(n47929) );
  NOR4X1 U51073 ( .A(n21737), .B(n21736), .C(n21735), .D(n21734), .Y(n47928)
         );
  NAND4X1 U51074 ( .A(n43245), .B(n43244), .C(n43243), .D(n43242), .Y(
        net213021) );
  XNOR2X1 U51075 ( .A(n33330), .B(n36726), .Y(n43244) );
  NOR2X1 U51076 ( .A(n31474), .B(n31473), .Y(n43243) );
  NOR4X1 U51077 ( .A(n31472), .B(n31471), .C(n31470), .D(n31469), .Y(n43242)
         );
  NAND4X1 U51078 ( .A(n46743), .B(n46742), .C(n46741), .D(n46740), .Y(n12901)
         );
  XNOR2X1 U51079 ( .A(n36733), .B(n33298), .Y(n46742) );
  NOR2X1 U51080 ( .A(n21536), .B(n21535), .Y(n46741) );
  NOR4X1 U51081 ( .A(n21534), .B(n21533), .C(n21532), .D(n21531), .Y(n46740)
         );
  NAND4X1 U51082 ( .A(n46733), .B(n46732), .C(n46731), .D(n46730), .Y(n48099)
         );
  XNOR2X1 U51083 ( .A(n36768), .B(n33321), .Y(n46732) );
  NOR2X1 U51084 ( .A(n21556), .B(n21555), .Y(n46731) );
  NOR4X1 U51085 ( .A(n21554), .B(n21553), .C(n21552), .D(n21551), .Y(n46730)
         );
  NAND4X1 U51086 ( .A(n47936), .B(n47935), .C(n47934), .D(n47933), .Y(n12896)
         );
  XNOR2X1 U51087 ( .A(n36734), .B(n33242), .Y(n47935) );
  NOR2X1 U51088 ( .A(n21729), .B(n21728), .Y(n47934) );
  NOR4X1 U51089 ( .A(n21727), .B(n21726), .C(n21725), .D(n21724), .Y(n47933)
         );
  NAND4X1 U51090 ( .A(n46738), .B(n46737), .C(n46736), .D(n46735), .Y(n12904)
         );
  XNOR2X1 U51091 ( .A(n36735), .B(n33306), .Y(n46737) );
  NOR2X1 U51092 ( .A(n21546), .B(n21545), .Y(n46736) );
  NOR4X1 U51093 ( .A(n21544), .B(n21543), .C(n21542), .D(n21541), .Y(n46735)
         );
  NAND4X1 U51094 ( .A(n46684), .B(n46683), .C(n46682), .D(n46681), .Y(n11335)
         );
  XNOR2X1 U51095 ( .A(n36733), .B(n33250), .Y(n46683) );
  NOR2X1 U51096 ( .A(n21709), .B(n21708), .Y(n46682) );
  NOR4X1 U51097 ( .A(n21707), .B(n21706), .C(n21705), .D(n21704), .Y(n46681)
         );
  NAND4X1 U51098 ( .A(n46904), .B(n46903), .C(n46902), .D(n46901), .Y(n13019)
         );
  XNOR2X1 U51099 ( .A(n36736), .B(n33218), .Y(n46903) );
  NOR2X1 U51100 ( .A(n21133), .B(n21132), .Y(n46902) );
  NOR4X1 U51101 ( .A(n21131), .B(n21130), .C(n21129), .D(n21128), .Y(n46901)
         );
  NOR2X1 U51102 ( .A(n10232), .B(n46739), .Y(n46743) );
  XOR2X1 U51103 ( .A(n36746), .B(n33300), .Y(n46739) );
  NOR2X1 U51104 ( .A(n10520), .B(n45974), .Y(n45978) );
  XOR2X1 U51105 ( .A(n33265), .B(n36776), .Y(n45974) );
  NOR2X1 U51106 ( .A(n10339), .B(n43182), .Y(n43186) );
  XOR2X1 U51107 ( .A(n33252), .B(n36825), .Y(n43182) );
  NOR2X1 U51108 ( .A(n10519), .B(n45954), .Y(n45958) );
  XOR2X1 U51109 ( .A(n33257), .B(n36780), .Y(n45954) );
  NOR2X1 U51110 ( .A(n10336), .B(n43187), .Y(n43191) );
  XOR2X1 U51111 ( .A(n33244), .B(n36829), .Y(n43187) );
  NOR2X1 U51112 ( .A(n11984), .B(n46794), .Y(n46798) );
  XOR2X1 U51113 ( .A(n41302), .B(n33172), .Y(n46794) );
  NOR2X1 U51114 ( .A(n11658), .B(n43352), .Y(n43356) );
  XOR2X1 U51115 ( .A(n33212), .B(n36828), .Y(n43352) );
  NOR2X1 U51116 ( .A(n11031), .B(n46885), .Y(n46889) );
  NOR2X1 U51117 ( .A(n11657), .B(n43343), .Y(n43347) );
  XOR2X1 U51118 ( .A(n33220), .B(n36831), .Y(n43343) );
  XNOR2X1 U51119 ( .A(n33313), .B(n36774), .Y(n46727) );
  NOR2X1 U51120 ( .A(n21566), .B(n21565), .Y(n46726) );
  NOR2X1 U51121 ( .A(n11040), .B(n46685), .Y(net212002) );
  NOR2X1 U51122 ( .A(n11991), .B(n45885), .Y(n45889) );
  XOR2X1 U51123 ( .A(n33209), .B(n36784), .Y(n45885) );
  NOR2X1 U51124 ( .A(n10525), .B(n45952), .Y(net213022) );
  XOR2X1 U51125 ( .A(n41301), .B(n33308), .Y(n45952) );
  NOR2X1 U51126 ( .A(n40399), .B(n46890), .Y(n46894) );
  XOR2X1 U51127 ( .A(n36767), .B(n33201), .Y(n46890) );
  NOR2X1 U51128 ( .A(n11988), .B(n45890), .Y(n45894) );
  XOR2X1 U51129 ( .A(n33201), .B(n36786), .Y(n45890) );
  NOR2X1 U51130 ( .A(n11673), .B(n43232), .Y(n43236) );
  NOR2X1 U51131 ( .A(n11650), .B(n43387), .Y(n43391) );
  XOR2X1 U51132 ( .A(n33180), .B(n36830), .Y(n43387) );
  NOR2X1 U51133 ( .A(n40390), .B(n47927), .Y(n47931) );
  XOR2X1 U51134 ( .A(n36768), .B(n33233), .Y(n47927) );
  NOR2X1 U51135 ( .A(n11050), .B(n47922), .Y(n47926) );
  NOR2X1 U51136 ( .A(n11672), .B(n43259), .Y(n43263) );
  XOR2X1 U51137 ( .A(n33348), .B(n36825), .Y(n43259) );
  NOR2X1 U51138 ( .A(n11994), .B(n45875), .Y(n45879) );
  XOR2X1 U51139 ( .A(n33225), .B(n36784), .Y(n45875) );
  NOR2X1 U51140 ( .A(n11652), .B(n43369), .Y(n43373) );
  NOR2X1 U51141 ( .A(n12389), .B(n46729), .Y(n46733) );
  NOR2X1 U51142 ( .A(n11030), .B(n46900), .Y(n46904) );
  XOR2X1 U51143 ( .A(n36772), .B(n33217), .Y(n46900) );
  NOR2X1 U51144 ( .A(n11651), .B(n43360), .Y(n43364) );
  XOR2X1 U51145 ( .A(n33204), .B(n36822), .Y(n43360) );
  NOR2X1 U51146 ( .A(n11649), .B(n43378), .Y(n43382) );
  XOR2X1 U51147 ( .A(n33188), .B(n36828), .Y(n43378) );
  NOR2X1 U51148 ( .A(n12800), .B(n46875), .Y(n46879) );
  XOR2X1 U51149 ( .A(n41303), .B(n33180), .Y(n46875) );
  NOR2X1 U51150 ( .A(n11669), .B(n43241), .Y(n43245) );
  XOR2X1 U51151 ( .A(n33332), .B(n36821), .Y(n43241) );
  NOR2X1 U51152 ( .A(n11039), .B(n46687), .Y(net211992) );
  XOR2X1 U51153 ( .A(n36767), .B(n33281), .Y(n46687) );
  NOR2X1 U51154 ( .A(n11990), .B(n45880), .Y(n45884) );
  NOR2X1 U51155 ( .A(n12274), .B(n46754), .Y(n46758) );
  NOR2X1 U51156 ( .A(n12006), .B(n45900), .Y(n45904) );
  NOR2X1 U51157 ( .A(n11989), .B(n45865), .Y(n45869) );
  XOR2X1 U51158 ( .A(n33193), .B(n36777), .Y(n45865) );
  NOR2X1 U51159 ( .A(n10340), .B(n44631), .Y(n44635) );
  XOR2X1 U51160 ( .A(n33236), .B(n36824), .Y(n44631) );
  NOR2X1 U51161 ( .A(n10341), .B(n43335), .Y(n43339) );
  NOR2X1 U51162 ( .A(n12255), .B(n46880), .Y(n46884) );
  XOR2X1 U51163 ( .A(n36747), .B(n33172), .Y(n46880) );
  NOR2X1 U51164 ( .A(n12474), .B(n44640), .Y(net214646) );
  XOR2X1 U51165 ( .A(n33276), .B(n36821), .Y(n44640) );
  NOR2X1 U51166 ( .A(n10527), .B(n45964), .Y(n45968) );
  XOR2X1 U51167 ( .A(n41300), .B(n33292), .Y(n45964) );
  NOR2X1 U51168 ( .A(n12485), .B(n43285), .Y(n43289) );
  NOR2X1 U51169 ( .A(n12260), .B(n47932), .Y(n47936) );
  NOR2X1 U51170 ( .A(n12668), .B(n45979), .Y(n45983) );
  XOR2X1 U51171 ( .A(n33241), .B(n36779), .Y(n45979) );
  NOR2X1 U51172 ( .A(n12672), .B(n45984), .Y(net212981) );
  XOR2X1 U51173 ( .A(n33273), .B(n36779), .Y(n45984) );
  NOR2X1 U51174 ( .A(n12665), .B(n45870), .Y(n45874) );
  NOR2X1 U51175 ( .A(n11023), .B(n46865), .Y(n46869) );
  XOR2X1 U51176 ( .A(n36750), .B(n33188), .Y(n46865) );
  NOR2X1 U51177 ( .A(n11052), .B(n46774), .Y(n46778) );
  NOR2X1 U51178 ( .A(n12675), .B(n45969), .Y(n45973) );
  NOR2X1 U51179 ( .A(n12671), .B(n45959), .Y(n45963) );
  NOR2X1 U51180 ( .A(n12482), .B(n43250), .Y(n43254) );
  NOR2X1 U51181 ( .A(n12476), .B(n43159), .Y(n43163) );
  XOR2X1 U51182 ( .A(n33292), .B(n36827), .Y(n43159) );
  NOR2X1 U51183 ( .A(n11661), .B(n43177), .Y(n43181) );
  NOR2X1 U51184 ( .A(n11662), .B(n44641), .Y(net214641) );
  XOR2X1 U51185 ( .A(n33268), .B(n36822), .Y(n44641) );
  NOR2X1 U51186 ( .A(n12004), .B(n45935), .Y(n45939) );
  XOR2X1 U51187 ( .A(n33345), .B(n36778), .Y(n45935) );
  NOR2X1 U51188 ( .A(n45925), .B(net209778), .Y(n45929) );
  NOR2X1 U51189 ( .A(n45985), .B(net209767), .Y(n45989) );
  XOR2X1 U51190 ( .A(n33233), .B(n36779), .Y(n45985) );
  NOR4X1 U51191 ( .A(n22653), .B(n22652), .C(n22651), .D(n22650), .Y(net212904) );
  XNOR2X1 U51192 ( .A(n36840), .B(n33042), .Y(net212912) );
  NOR2X1 U51193 ( .A(n22675), .B(n22674), .Y(net212913) );
  NOR4X1 U51194 ( .A(n32314), .B(n32313), .C(n32312), .D(n32311), .Y(net216871) );
  XNOR2X1 U51195 ( .A(n33058), .B(n42565), .Y(net216878) );
  NOR2X1 U51196 ( .A(n32346), .B(n32345), .Y(net216879) );
  NOR4X1 U51197 ( .A(n32344), .B(n32343), .C(n32342), .D(n32341), .Y(net216880) );
  NOR4X1 U51198 ( .A(n22612), .B(n22611), .C(n22610), .D(n22609), .Y(net212864) );
  NOR4X1 U51199 ( .A(n22622), .B(n22621), .C(n22620), .D(n22619), .Y(net212869) );
  NOR4X1 U51200 ( .A(n32014), .B(n32013), .C(n32012), .D(n32011), .Y(net216817) );
  NOR4X1 U51201 ( .A(n22663), .B(n22662), .C(n22661), .D(n22660), .Y(net212909) );
  NOR4X1 U51202 ( .A(n22643), .B(n22642), .C(n22641), .D(n22640), .Y(net212899) );
  NAND4X1 U51203 ( .A(n46068), .B(n46067), .C(n46066), .D(n46065), .Y(n10996)
         );
  XNOR2X1 U51204 ( .A(n36847), .B(n33018), .Y(n46067) );
  NOR2X1 U51205 ( .A(n22574), .B(n22573), .Y(n46066) );
  NOR4X1 U51206 ( .A(n22572), .B(n22571), .C(n22570), .D(n22569), .Y(n46065)
         );
  NAND4X1 U51207 ( .A(n43427), .B(n43426), .C(n43425), .D(n43424), .Y(n11955)
         );
  NOR2X1 U51208 ( .A(n30873), .B(n30872), .Y(n43425) );
  NOR4X1 U51209 ( .A(n30871), .B(n30870), .C(n30869), .D(n30868), .Y(n43424)
         );
  NAND4X1 U51210 ( .A(n46044), .B(n46043), .C(n46042), .D(n46041), .Y(n11017)
         );
  XNOR2X1 U51211 ( .A(n36845), .B(n33146), .Y(n46043) );
  NOR2X1 U51212 ( .A(n22695), .B(n22694), .Y(n46042) );
  NOR4X1 U51213 ( .A(n22693), .B(n22692), .C(n22691), .D(n22690), .Y(n46041)
         );
  NAND4X1 U51214 ( .A(n46073), .B(n46072), .C(n46071), .D(n46070), .Y(n10997)
         );
  XNOR2X1 U51215 ( .A(n36838), .B(n33010), .Y(n46072) );
  NOR2X1 U51216 ( .A(n22564), .B(n22563), .Y(n46071) );
  NOR4X1 U51217 ( .A(n22562), .B(n22561), .C(n22560), .D(n22559), .Y(n46070)
         );
  NAND4X1 U51218 ( .A(n46009), .B(n46008), .C(n46007), .D(n46006), .Y(n11006)
         );
  XNOR2X1 U51219 ( .A(n36846), .B(n33082), .Y(n46008) );
  NOR2X1 U51220 ( .A(n22765), .B(n22764), .Y(n46007) );
  NOR4X1 U51221 ( .A(n22763), .B(n22762), .C(n22761), .D(n22760), .Y(n46006)
         );
  NOR4X1 U51222 ( .A(n22632), .B(n22631), .C(n22630), .D(n22629), .Y(net212874) );
  NAND4X1 U51223 ( .A(n43099), .B(n43098), .C(n43097), .D(n43096), .Y(n11979)
         );
  XNOR2X1 U51224 ( .A(n33154), .B(n42565), .Y(n43098) );
  NOR2X1 U51225 ( .A(n32136), .B(n32135), .Y(n43097) );
  NOR4X1 U51226 ( .A(n32134), .B(n32133), .C(n32132), .D(n32131), .Y(n43096)
         );
  NOR4X1 U51227 ( .A(n30751), .B(n30750), .C(n30749), .D(n30748), .Y(net216511) );
  NAND4X1 U51228 ( .A(n43145), .B(n43144), .C(n43143), .D(n43142), .Y(n10501)
         );
  XNOR2X1 U51229 ( .A(n33050), .B(n36726), .Y(n43144) );
  NOR2X1 U51230 ( .A(n31956), .B(n31955), .Y(n43143) );
  NOR4X1 U51231 ( .A(n31954), .B(n31953), .C(n31952), .D(n31951), .Y(n43142)
         );
  NOR4X1 U51232 ( .A(n31984), .B(n31983), .C(n31982), .D(n31981), .Y(net216808) );
  NAND4X1 U51233 ( .A(n43108), .B(n43107), .C(n43106), .D(n43105), .Y(n11976)
         );
  XNOR2X1 U51234 ( .A(n33146), .B(n42565), .Y(n43107) );
  NOR2X1 U51235 ( .A(n32106), .B(n32105), .Y(n43106) );
  NOR4X1 U51236 ( .A(n32104), .B(n32103), .C(n32102), .D(n32101), .Y(n43105)
         );
  NOR4X1 U51237 ( .A(n30721), .B(n30720), .C(n30719), .D(n30718), .Y(net216502) );
  NAND4X1 U51238 ( .A(n43154), .B(n43153), .C(n43152), .D(n43151), .Y(n10506)
         );
  XNOR2X1 U51239 ( .A(n33114), .B(n36725), .Y(n43153) );
  NOR2X1 U51240 ( .A(n31926), .B(n31925), .Y(n43152) );
  NOR4X1 U51241 ( .A(n31924), .B(n31923), .C(n31922), .D(n31921), .Y(n43151)
         );
  NOR2X1 U51242 ( .A(n22725), .B(n22724), .Y(n46027) );
  NOR4X1 U51243 ( .A(n22723), .B(n22722), .C(n22721), .D(n22720), .Y(n46026)
         );
  NAND4X1 U51244 ( .A(n43400), .B(n43399), .C(n43398), .D(n43397), .Y(n11985)
         );
  XNOR2X1 U51245 ( .A(n33170), .B(n42569), .Y(n43399) );
  NOR2X1 U51246 ( .A(n30933), .B(n30932), .Y(n43398) );
  NOR4X1 U51247 ( .A(n30931), .B(n30930), .C(n30929), .D(n30928), .Y(n43397)
         );
  NAND4X1 U51248 ( .A(n46063), .B(n46062), .C(n46061), .D(n46060), .Y(n11002)
         );
  XNOR2X1 U51249 ( .A(n36844), .B(n33026), .Y(n46062) );
  NOR2X1 U51250 ( .A(n22584), .B(n22583), .Y(n46061) );
  NOR4X1 U51251 ( .A(n22582), .B(n22581), .C(n22580), .D(n22579), .Y(n46060)
         );
  NAND4X1 U51252 ( .A(n46004), .B(n46003), .C(n46002), .D(n46001), .Y(n12391)
         );
  XNOR2X1 U51253 ( .A(n36845), .B(n33090), .Y(n46003) );
  NOR2X1 U51254 ( .A(n22775), .B(n22774), .Y(n46002) );
  NOR4X1 U51255 ( .A(n22773), .B(n22772), .C(n22771), .D(n22770), .Y(n46001)
         );
  NOR4X1 U51256 ( .A(n22753), .B(n22752), .C(n22751), .D(n22750), .Y(n46011)
         );
  NAND4X1 U51257 ( .A(n46049), .B(n46048), .C(n46047), .D(n46046), .Y(n11018)
         );
  XNOR2X1 U51258 ( .A(n36837), .B(n33138), .Y(n46048) );
  NOR2X1 U51259 ( .A(n22685), .B(n22684), .Y(n46047) );
  NOR4X1 U51260 ( .A(n22683), .B(n22682), .C(n22681), .D(n22680), .Y(n46046)
         );
  NAND4X1 U51261 ( .A(n43126), .B(n43125), .C(n43124), .D(n43123), .Y(n12801)
         );
  XNOR2X1 U51262 ( .A(n33122), .B(n36725), .Y(n43125) );
  NOR2X1 U51263 ( .A(n32046), .B(n32045), .Y(n43124) );
  NOR4X1 U51264 ( .A(n32044), .B(n32043), .C(n32042), .D(n32041), .Y(n43123)
         );
  NOR2X1 U51265 ( .A(n22705), .B(n22704), .Y(n46037) );
  NOR4X1 U51266 ( .A(n22703), .B(n22702), .C(n22701), .D(n22700), .Y(n46036)
         );
  NAND4X1 U51267 ( .A(n43091), .B(n43090), .C(n43089), .D(n43088), .Y(n11978)
         );
  XNOR2X1 U51268 ( .A(n33162), .B(n42565), .Y(n43090) );
  NOR2X1 U51269 ( .A(n32166), .B(n32165), .Y(n43089) );
  NOR4X1 U51270 ( .A(n32164), .B(n32163), .C(n32162), .D(n32161), .Y(n43088)
         );
  NOR4X1 U51271 ( .A(n30781), .B(n30780), .C(n30779), .D(n30778), .Y(net216520) );
  NAND4X1 U51272 ( .A(n45994), .B(n45993), .C(n45992), .D(n45991), .Y(n11007)
         );
  XNOR2X1 U51273 ( .A(n36844), .B(n33074), .Y(n45993) );
  NOR2X1 U51274 ( .A(n22795), .B(n22794), .Y(n45992) );
  NOR4X1 U51275 ( .A(n22793), .B(n22792), .C(n22791), .D(n22790), .Y(n45991)
         );
  NAND4X1 U51276 ( .A(n43072), .B(n43071), .C(n43070), .D(n43069), .Y(n11970)
         );
  XNOR2X1 U51277 ( .A(n33090), .B(n42565), .Y(n43071) );
  NOR2X1 U51278 ( .A(n32196), .B(n32195), .Y(n43070) );
  NOR4X1 U51279 ( .A(n32194), .B(n32193), .C(n32192), .D(n32191), .Y(n43069)
         );
  NAND4X1 U51280 ( .A(n43117), .B(n43116), .C(n43115), .D(n43114), .Y(n11977)
         );
  XNOR2X1 U51281 ( .A(n33138), .B(n36726), .Y(n43116) );
  NOR2X1 U51282 ( .A(n32076), .B(n32075), .Y(n43115) );
  NOR4X1 U51283 ( .A(n32074), .B(n32073), .C(n32072), .D(n32071), .Y(n43114)
         );
  XNOR2X1 U51284 ( .A(n33010), .B(n42569), .Y(net216491) );
  NOR2X1 U51285 ( .A(n30693), .B(n30692), .Y(net216492) );
  NAND4X1 U51286 ( .A(n46019), .B(n46018), .C(n46017), .D(n46016), .Y(n11015)
         );
  XNOR2X1 U51287 ( .A(n36843), .B(n33130), .Y(n46018) );
  NOR2X1 U51288 ( .A(n22745), .B(n22744), .Y(n46017) );
  NOR4X1 U51289 ( .A(n22743), .B(n22742), .C(n22741), .D(n22740), .Y(n46016)
         );
  NAND4X1 U51290 ( .A(n46058), .B(n46057), .C(n46056), .D(n46055), .Y(n11001)
         );
  XNOR2X1 U51291 ( .A(n36841), .B(n33034), .Y(n46057) );
  NOR2X1 U51292 ( .A(n22594), .B(n22593), .Y(n46056) );
  NOR4X1 U51293 ( .A(n22592), .B(n22591), .C(n22590), .D(n22589), .Y(n46055)
         );
  NOR4X1 U51294 ( .A(n22733), .B(n22732), .C(n22731), .D(n22730), .Y(n46021)
         );
  XNOR2X1 U51295 ( .A(n33082), .B(n42560), .Y(net216914) );
  NOR2X1 U51296 ( .A(n32286), .B(n32285), .Y(net216915) );
  NOR4X1 U51297 ( .A(n32284), .B(n32283), .C(n32282), .D(n32281), .Y(net216916) );
  NAND4X1 U51298 ( .A(n43063), .B(n43062), .C(n43061), .D(n43060), .Y(n11969)
         );
  XNOR2X1 U51299 ( .A(n33098), .B(n42565), .Y(n43062) );
  NOR2X1 U51300 ( .A(n32226), .B(n32225), .Y(n43061) );
  NOR4X1 U51301 ( .A(n32224), .B(n32223), .C(n32222), .D(n32221), .Y(n43060)
         );
  NOR4X1 U51302 ( .A(n21686), .B(n21685), .C(n21684), .D(n21683), .Y(net211965) );
  NOR4X1 U51303 ( .A(n32254), .B(n32253), .C(n32252), .D(n32251), .Y(net216907) );
  XNOR2X1 U51304 ( .A(n36767), .B(n33089), .Y(n46837) );
  NOR2X1 U51305 ( .A(n21345), .B(n21344), .Y(n46836) );
  NAND4X1 U51306 ( .A(n44630), .B(n44629), .C(n44628), .D(n44627), .Y(
        net210704) );
  XNOR2X1 U51307 ( .A(n33066), .B(n42560), .Y(n44629) );
  NOR2X1 U51308 ( .A(n31896), .B(n31895), .Y(n44628) );
  NOR4X1 U51309 ( .A(n31894), .B(n31893), .C(n31892), .D(n31891), .Y(n44627)
         );
  NOR2X1 U51310 ( .A(n21618), .B(n21617), .Y(net211969) );
  NOR4X1 U51311 ( .A(n21616), .B(n21615), .C(n21614), .D(n21613), .Y(net211970) );
  NAND4X1 U51312 ( .A(n43432), .B(n43431), .C(n43430), .D(n43429), .Y(n12651)
         );
  NOR2X1 U51313 ( .A(n30843), .B(n30842), .Y(n43430) );
  NOR4X1 U51314 ( .A(n30841), .B(n30840), .C(n30839), .D(n30838), .Y(n43429)
         );
  NAND4X1 U51315 ( .A(n45999), .B(n45998), .C(n45997), .D(n45996), .Y(n12246)
         );
  XNOR2X1 U51316 ( .A(n36846), .B(n33098), .Y(n45998) );
  NOR2X1 U51317 ( .A(n22785), .B(n22784), .Y(n45997) );
  NOR4X1 U51318 ( .A(n22783), .B(n22782), .C(n22781), .D(n22780), .Y(n45996)
         );
  NAND4X1 U51319 ( .A(n46793), .B(n46792), .C(n46791), .D(n46790), .Y(n11317)
         );
  XNOR2X1 U51320 ( .A(n36734), .B(n33138), .Y(n46792) );
  NOR2X1 U51321 ( .A(n21435), .B(n21434), .Y(n46791) );
  NOR4X1 U51322 ( .A(n21433), .B(n21432), .C(n21431), .D(n21430), .Y(n46790)
         );
  NAND4X1 U51323 ( .A(n46034), .B(n46033), .C(n46032), .D(n46031), .Y(n12252)
         );
  XNOR2X1 U51324 ( .A(n36841), .B(n33162), .Y(n46033) );
  NOR2X1 U51325 ( .A(n22715), .B(n22714), .Y(n46032) );
  NOR4X1 U51326 ( .A(n22713), .B(n22712), .C(n22711), .D(n22710), .Y(n46031)
         );
  NAND4X1 U51327 ( .A(n46803), .B(n46802), .C(n46801), .D(n46800), .Y(n12887)
         );
  XNOR2X1 U51328 ( .A(n36736), .B(n33162), .Y(n46802) );
  NOR2X1 U51329 ( .A(n21425), .B(n21424), .Y(n46801) );
  NOR4X1 U51330 ( .A(n21423), .B(n21422), .C(n21421), .D(n21420), .Y(n46800)
         );
  NOR2X1 U51331 ( .A(n21234), .B(n21233), .Y(net211795) );
  NOR4X1 U51332 ( .A(n21232), .B(n21231), .C(n21230), .D(n21229), .Y(net211796) );
  NOR2X1 U51333 ( .A(n21648), .B(n21647), .Y(net211984) );
  XNOR2X1 U51334 ( .A(n36734), .B(n33018), .Y(net211973) );
  NOR2X1 U51335 ( .A(n21628), .B(n21627), .Y(net211974) );
  NOR4X1 U51336 ( .A(n21626), .B(n21625), .C(n21624), .D(n21623), .Y(net211975) );
  NAND4X1 U51337 ( .A(n46788), .B(n46787), .C(n46786), .D(n46785), .Y(n11316)
         );
  XNOR2X1 U51338 ( .A(n36734), .B(n33146), .Y(n46787) );
  NOR2X1 U51339 ( .A(n21445), .B(n21444), .Y(n46786) );
  NOR4X1 U51340 ( .A(n21443), .B(n21442), .C(n21441), .D(n21440), .Y(n46785)
         );
  NOR4X1 U51341 ( .A(n21403), .B(n21402), .C(n21401), .D(n21400), .Y(net210510) );
  NOR2X1 U51342 ( .A(n21678), .B(n21677), .Y(net211959) );
  XNOR2X1 U51343 ( .A(n36734), .B(n33130), .Y(n46812) );
  NOR2X1 U51344 ( .A(n21395), .B(n21394), .Y(n46811) );
  NOR4X1 U51345 ( .A(n21393), .B(n21392), .C(n21391), .D(n21390), .Y(n46810)
         );
  NOR2X1 U51346 ( .A(n21183), .B(n21182), .Y(n46872) );
  NOR4X1 U51347 ( .A(n21181), .B(n21180), .C(n21179), .D(n21178), .Y(n46871)
         );
  NAND4X1 U51348 ( .A(n47833), .B(n47832), .C(n47831), .D(n47830), .Y(n10013)
         );
  XNOR2X1 U51349 ( .A(n36733), .B(n33114), .Y(n47832) );
  NOR2X1 U51350 ( .A(n21295), .B(n21294), .Y(n47831) );
  NOR4X1 U51351 ( .A(n21293), .B(n21292), .C(n21291), .D(n21290), .Y(n47830)
         );
  NOR2X1 U51352 ( .A(n21325), .B(n21324), .Y(n47939) );
  NOR4X1 U51353 ( .A(n21323), .B(n21322), .C(n21321), .D(n21320), .Y(n47938)
         );
  NAND4X1 U51354 ( .A(n46848), .B(n46847), .C(n46846), .D(n46845), .Y(n12872)
         );
  NOR2X1 U51355 ( .A(n21305), .B(n21304), .Y(n46846) );
  NOR4X1 U51356 ( .A(n21303), .B(n21302), .C(n21301), .D(n21300), .Y(n46845)
         );
  XNOR2X1 U51357 ( .A(n36736), .B(n33154), .Y(n46807) );
  NOR2X1 U51358 ( .A(n21415), .B(n21414), .Y(n46806) );
  NOR4X1 U51359 ( .A(n21413), .B(n21412), .C(n21411), .D(n21410), .Y(n46805)
         );
  NAND4X1 U51360 ( .A(n46694), .B(n46693), .C(n46692), .D(n46691), .Y(n13021)
         );
  NOR2X1 U51361 ( .A(n21638), .B(n21637), .Y(n46692) );
  NOR4X1 U51362 ( .A(n21636), .B(n21635), .C(n21634), .D(n21633), .Y(n46691)
         );
  NAND4X1 U51363 ( .A(n46833), .B(n46832), .C(n46831), .D(n46830), .Y(
        net210047) );
  XNOR2X1 U51364 ( .A(n36773), .B(n33097), .Y(n46832) );
  NOR2X1 U51365 ( .A(n21355), .B(n21354), .Y(n46831) );
  NOR4X1 U51366 ( .A(n21353), .B(n21352), .C(n21351), .D(n21350), .Y(n46830)
         );
  NAND4X1 U51367 ( .A(n46823), .B(n46822), .C(n46821), .D(n46820), .Y(
        net210043) );
  XNOR2X1 U51368 ( .A(n36770), .B(n33065), .Y(n46822) );
  NOR2X1 U51369 ( .A(n21375), .B(n21374), .Y(n46821) );
  NOR4X1 U51370 ( .A(n21373), .B(n21372), .C(n21371), .D(n21370), .Y(n46820)
         );
  XNOR2X1 U51371 ( .A(n36734), .B(n33082), .Y(n47945) );
  NOR2X1 U51372 ( .A(n21335), .B(n21334), .Y(n47944) );
  NOR4X1 U51373 ( .A(n21333), .B(n21332), .C(n21331), .D(n21330), .Y(n47943)
         );
  NAND4X1 U51374 ( .A(n46843), .B(n46842), .C(n46841), .D(n46840), .Y(n12876)
         );
  NOR2X1 U51375 ( .A(n21315), .B(n21314), .Y(n46841) );
  NOR4X1 U51376 ( .A(n21313), .B(n21312), .C(n21311), .D(n21310), .Y(n46840)
         );
  XNOR2X1 U51377 ( .A(n36736), .B(n33122), .Y(n46817) );
  NOR2X1 U51378 ( .A(n21385), .B(n21384), .Y(n46816) );
  NOR4X1 U51379 ( .A(n21383), .B(n21382), .C(n21381), .D(n21380), .Y(n46815)
         );
  NOR2X1 U51380 ( .A(n10274), .B(n46844), .Y(n46848) );
  NOR2X1 U51381 ( .A(n10502), .B(n46054), .Y(n46058) );
  NOR2X1 U51382 ( .A(n10503), .B(n46052), .Y(net212901) );
  NOR2X1 U51383 ( .A(n10425), .B(n43423), .Y(n43427) );
  NOR2X1 U51384 ( .A(n10504), .B(n45995), .Y(n45999) );
  NOR2X1 U51385 ( .A(n10810), .B(n46839), .Y(n46843) );
  NOR2X1 U51386 ( .A(n10996), .B(n46696), .Y(net211967) );
  NOR2X1 U51387 ( .A(n11017), .B(n46789), .Y(n46793) );
  XOR2X1 U51388 ( .A(n36774), .B(n33137), .Y(n46789) );
  NOR2X1 U51389 ( .A(net260251), .B(n46075), .Y(net212866) );
  NOR2X1 U51390 ( .A(n11646), .B(n43104), .Y(n43108) );
  NOR2X1 U51391 ( .A(n11006), .B(n47937), .Y(n47941) );
  NOR2X1 U51392 ( .A(n10806), .B(n46698), .Y(net211957) );
  NOR2X1 U51393 ( .A(n11645), .B(n43095), .Y(n43099) );
  XOR2X1 U51394 ( .A(n33156), .B(n36829), .Y(n43095) );
  XNOR2X1 U51395 ( .A(n36764), .B(n33057), .Y(n46827) );
  NOR2X1 U51396 ( .A(n21365), .B(n21364), .Y(n46826) );
  NOR2X1 U51397 ( .A(n11979), .B(n46040), .Y(n46044) );
  NOR2X1 U51398 ( .A(n11961), .B(n46064), .Y(n46068) );
  NOR2X1 U51399 ( .A(n10501), .B(n46050), .Y(net212911) );
  NOR2X1 U51400 ( .A(n10505), .B(n46025), .Y(n46029) );
  NOR2X1 U51401 ( .A(n11016), .B(n47829), .Y(n47833) );
  NOR2X1 U51402 ( .A(n11976), .B(n46045), .Y(n46049) );
  NOR2X1 U51403 ( .A(n11958), .B(n46069), .Y(n46073) );
  NOR2X1 U51404 ( .A(n11638), .B(n43150), .Y(n43154) );
  NOR2X1 U51405 ( .A(n11625), .B(n43407), .Y(net216499) );
  NOR2X1 U51406 ( .A(n10506), .B(n46020), .Y(n46024) );
  NOR2X1 U51407 ( .A(n11002), .B(n46695), .Y(net211972) );
  NOR2X1 U51408 ( .A(n11985), .B(n46030), .Y(n46034) );
  XOR2X1 U51409 ( .A(n36918), .B(n33164), .Y(n46030) );
  NOR2X1 U51410 ( .A(n12391), .B(n47942), .Y(n47946) );
  NOR2X1 U51411 ( .A(n40395), .B(n47791), .Y(net210507) );
  XOR2X1 U51412 ( .A(n36764), .B(n33105), .Y(n47791) );
  NOR2X1 U51413 ( .A(n12390), .B(n46784), .Y(n46788) );
  NOR2X1 U51414 ( .A(n11626), .B(n43406), .Y(net216508) );
  XOR2X1 U51415 ( .A(n33028), .B(n36829), .Y(n43406) );
  NOR2X1 U51416 ( .A(n11640), .B(n43136), .Y(net216805) );
  NOR2X1 U51417 ( .A(n11622), .B(n43408), .Y(net216490) );
  NOR2X1 U51418 ( .A(n11639), .B(n43113), .Y(n43117) );
  XOR2X1 U51419 ( .A(n33140), .B(n36824), .Y(n43113) );
  NOR2X1 U51420 ( .A(n11637), .B(n43122), .Y(n43126) );
  NOR2X1 U51421 ( .A(n40388), .B(n46010), .Y(n46014) );
  NOR2X1 U51422 ( .A(n11621), .B(n43428), .Y(n43432) );
  NOR2X1 U51423 ( .A(n11960), .B(n46059), .Y(n46063) );
  NOR2X1 U51424 ( .A(n11978), .B(n46035), .Y(n46039) );
  XOR2X1 U51425 ( .A(n33153), .B(n36777), .Y(n46035) );
  NOR2X1 U51426 ( .A(n11024), .B(n46870), .Y(n46874) );
  NOR2X1 U51427 ( .A(net260277), .B(n46005), .Y(n46009) );
  NOR2X1 U51428 ( .A(n11977), .B(n46015), .Y(n46019) );
  NOR2X1 U51429 ( .A(n11959), .B(n46074), .Y(net212871) );
  NOR2X1 U51430 ( .A(n11015), .B(n46814), .Y(n46818) );
  XOR2X1 U51431 ( .A(n36771), .B(n33121), .Y(n46814) );
  NOR2X1 U51432 ( .A(n40400), .B(n46690), .Y(n46694) );
  NOR2X1 U51433 ( .A(n11967), .B(n45990), .Y(n45994) );
  NOR2X1 U51434 ( .A(n11969), .B(n46000), .Y(n46004) );
  NOR2X1 U51435 ( .A(n11968), .B(n46051), .Y(net212906) );
  NOR2X1 U51436 ( .A(n12457), .B(n43049), .Y(net216913) );
  NOR2X1 U51437 ( .A(n12452), .B(n43141), .Y(n43145) );
  NOR2X1 U51438 ( .A(n12459), .B(n43068), .Y(n43072) );
  NOR2X1 U51439 ( .A(n12455), .B(n43077), .Y(net216877) );
  NOR2X1 U51440 ( .A(n12252), .B(n46804), .Y(n46808) );
  XOR2X1 U51441 ( .A(n36766), .B(n33153), .Y(n46804) );
  NOR2X1 U51442 ( .A(n12588), .B(n43087), .Y(n43091) );
  NOR2X1 U51443 ( .A(n12589), .B(n43059), .Y(n43063) );
  NOR2X1 U51444 ( .A(net260427), .B(n46076), .Y(net212861) );
  NOR2X1 U51445 ( .A(n12466), .B(n43396), .Y(n43400) );
  NOR2X1 U51446 ( .A(n12461), .B(n43131), .Y(net216814) );
  NOR2X1 U51447 ( .A(n12449), .B(n43405), .Y(net216517) );
  XOR2X1 U51448 ( .A(n33036), .B(n36830), .Y(n43405) );
  NOR2X1 U51449 ( .A(n12453), .B(n43082), .Y(net216868) );
  NOR2X1 U51450 ( .A(n46053), .B(net261020), .Y(net212896) );
  NOR2X1 U51451 ( .A(n43054), .B(net214724), .Y(net216904) );
  XOR2X1 U51452 ( .A(n33076), .B(n36831), .Y(n43054) );
  NOR2X1 U51453 ( .A(n44626), .B(net214669), .Y(n44630) );
  NOR4X1 U51454 ( .A(n24353), .B(n24352), .C(n24351), .D(n24350), .Y(net213515) );
  NOR4X1 U51455 ( .A(n24343), .B(n24342), .C(n24341), .D(n24340), .Y(net213510) );
  NOR2X1 U51456 ( .A(n23352), .B(n23351), .Y(net213197) );
  NOR4X1 U51457 ( .A(n23350), .B(n23349), .C(n23348), .D(n23347), .Y(net213198) );
  NOR2X1 U51458 ( .A(n23342), .B(n23340), .Y(net213192) );
  NOR4X1 U51459 ( .A(n23339), .B(n23338), .C(n23337), .D(n23336), .Y(net213193) );
  OAI211X1 U51460 ( .A0(n9738), .A1(n41199), .B0(n9740), .C0(n9741), .Y(
        nxt_data_num[1]) );
  AOI33X1 U51461 ( .A0(net171349), .A1(n50141), .A2(n9707), .B0(n50129), .B1(
        n9737), .B2(n41790), .Y(n9740) );
  AOI222XL U51462 ( .A0(n9742), .A1(n9743), .B0(n9744), .B1(n50134), .C0(
        n41789), .C1(n32399), .Y(n9741) );
  NOR4X1 U51463 ( .A(n30630), .B(n30629), .C(n30628), .D(n30627), .Y(net216394) );
  NOR2X1 U51464 ( .A(n23362), .B(n23361), .Y(net213202) );
  NOR4X1 U51465 ( .A(n23360), .B(n23359), .C(n23358), .D(n23357), .Y(net213203) );
  NOR2X1 U51466 ( .A(n29879), .B(n29878), .Y(net214685) );
  NOR4X1 U51467 ( .A(n29877), .B(n29876), .C(n29875), .D(n29874), .Y(net214686) );
  NOR2X1 U51468 ( .A(n24195), .B(n24194), .Y(n46646) );
  NOR4X1 U51469 ( .A(n24193), .B(n24192), .C(n24191), .D(n24190), .Y(n46645)
         );
  NOR4X1 U51470 ( .A(n22541), .B(n22540), .C(n22539), .D(n22538), .Y(net212834) );
  NOR4X1 U51471 ( .A(n22531), .B(n22530), .C(n22529), .D(n22528), .Y(net212829) );
  NOR4X1 U51472 ( .A(n30660), .B(n30659), .C(n30658), .D(n30657), .Y(net216403) );
  NOR2X1 U51473 ( .A(n29939), .B(n29938), .Y(net214674) );
  NOR4X1 U51474 ( .A(n29937), .B(n29936), .C(n29935), .D(n29934), .Y(net214675) );
  NOR2X1 U51475 ( .A(n24185), .B(n24184), .Y(n45614) );
  NOR4X1 U51476 ( .A(n24183), .B(n24182), .C(n24181), .D(n24180), .Y(n45613)
         );
  NOR2X1 U51477 ( .A(n29909), .B(n29908), .Y(net214680) );
  NOR4X1 U51478 ( .A(n29907), .B(n29906), .C(n29905), .D(n29904), .Y(net214681) );
  NOR4X1 U51479 ( .A(n22551), .B(n22550), .C(n22549), .D(n22548), .Y(net212839) );
  NOR2X1 U51480 ( .A(n29638), .B(n29637), .Y(net214690) );
  NOR4X1 U51481 ( .A(n29636), .B(n29635), .C(n29634), .D(n29633), .Y(net214691) );
  NOR4X1 U51482 ( .A(n24455), .B(n24454), .C(n24453), .D(n24452), .Y(net213535) );
  NAND4X1 U51483 ( .A(n47274), .B(n47273), .C(n47272), .D(n47271), .Y(n10448)
         );
  NOR2X1 U51484 ( .A(n26449), .B(n26448), .Y(n47272) );
  NOR4X1 U51485 ( .A(n26447), .B(n26446), .C(n26445), .D(n26444), .Y(n47271)
         );
  NOR2X1 U51486 ( .A(n25908), .B(n25907), .Y(net214999) );
  NOR4X1 U51487 ( .A(n25906), .B(n25905), .C(n25904), .D(n25903), .Y(net215000) );
  NOR4X1 U51488 ( .A(n24445), .B(n24444), .C(n24443), .D(n24442), .Y(net213530) );
  NOR2X1 U51489 ( .A(n23300), .B(n23299), .Y(net213217) );
  NOR4X1 U51490 ( .A(n23298), .B(n23297), .C(n23296), .D(n23295), .Y(net213218) );
  NOR2X1 U51491 ( .A(n24235), .B(n24234), .Y(net213469) );
  NOR4X1 U51492 ( .A(n22521), .B(n22520), .C(n22519), .D(n22518), .Y(net212859) );
  NOR2X1 U51493 ( .A(n30210), .B(n30209), .Y(net216348) );
  NAND4X1 U51494 ( .A(n44619), .B(n44618), .C(n44617), .D(n44616), .Y(n12170)
         );
  NOR2X1 U51495 ( .A(n29668), .B(n29667), .Y(n44617) );
  NOR4X1 U51496 ( .A(n29666), .B(n29665), .C(n29664), .D(n29663), .Y(n44616)
         );
  NOR2X1 U51497 ( .A(n30149), .B(n30148), .Y(net216303) );
  NOR4X1 U51498 ( .A(n30147), .B(n30146), .C(n30145), .D(n30144), .Y(net216304) );
  NOR4X1 U51499 ( .A(n24363), .B(n24362), .C(n24361), .D(n24360), .Y(net213520) );
  NOR2X1 U51500 ( .A(n26298), .B(n26297), .Y(net215116) );
  NOR4X1 U51501 ( .A(n26296), .B(n26295), .C(n26294), .D(n26293), .Y(net215117) );
  NOR2X1 U51502 ( .A(n24245), .B(n24244), .Y(net213474) );
  NOR4X1 U51503 ( .A(n24243), .B(n24242), .C(n24241), .D(n24240), .Y(net213475) );
  NOR4X1 U51504 ( .A(n22511), .B(n22510), .C(n22509), .D(n22508), .Y(net212854) );
  NOR4X1 U51505 ( .A(n24475), .B(n24474), .C(n24473), .D(n24472), .Y(net213565) );
  NOR2X1 U51506 ( .A(n23311), .B(n23309), .Y(net213227) );
  NOR4X1 U51507 ( .A(n23308), .B(n23307), .C(n23306), .D(n23305), .Y(net213228) );
  NOR4X1 U51508 ( .A(n22501), .B(n22500), .C(n22499), .D(n22498), .Y(net212849) );
  NOR2X1 U51509 ( .A(n21274), .B(n21273), .Y(net211775) );
  NOR4X1 U51510 ( .A(n24323), .B(n24322), .C(n24321), .D(n24320), .Y(net213490) );
  NAND4X1 U51511 ( .A(n44325), .B(n44324), .C(n44323), .D(n44322), .Y(n10447)
         );
  NOR2X1 U51512 ( .A(n26509), .B(n26508), .Y(n44323) );
  NOR4X1 U51513 ( .A(n26507), .B(n26506), .C(n26505), .D(n26504), .Y(n44322)
         );
  NOR4X1 U51514 ( .A(n24465), .B(n24464), .C(n24463), .D(n24462), .Y(net213560) );
  NOR2X1 U51515 ( .A(n21882), .B(n21881), .Y(net212096) );
  NOR4X1 U51516 ( .A(n24435), .B(n24434), .C(n24433), .D(n24432), .Y(net213555) );
  XNOR2X1 U51517 ( .A(n36734), .B(n32810), .Y(net212120) );
  NOR2X1 U51518 ( .A(n21943), .B(n21942), .Y(net212121) );
  NOR4X1 U51519 ( .A(n21941), .B(n21940), .C(n21939), .D(n21938), .Y(net212122) );
  NOR2X1 U51520 ( .A(n26388), .B(n26387), .Y(net215143) );
  NOR4X1 U51521 ( .A(n26386), .B(n26385), .C(n26384), .D(n26383), .Y(net215144) );
  AOI222XL U51522 ( .A0(net221892), .A1(n51092), .B0(n40192), .B1(n51091),
        .C0(n40377), .C1(n51090), .Y(n15017) );
  AOI222XL U51523 ( .A0(net221892), .A1(n50878), .B0(net218074), .B1(n50877),
        .C0(n40356), .C1(n50876), .Y(n15020) );
  AOI222XL U51524 ( .A0(net221892), .A1(n50664), .B0(net218118), .B1(n50663),
        .C0(n40377), .C1(n50662), .Y(n15026) );
  AOI222XL U51525 ( .A0(net221892), .A1(n50455), .B0(net217988), .B1(n50454),
        .C0(n40363), .C1(n50453), .Y(n15005) );
  OA22X1 U51526 ( .A0(net263805), .A1(n32929), .B0(n32937), .B1(n40050), .Y(
        n14764) );
  AOI222XL U51527 ( .A0(net266081), .A1(n50451), .B0(n40186), .B1(n50450),
        .C0(net216992), .C1(n50449), .Y(n14765) );
  AOI222XL U51528 ( .A0(net265891), .A1(n36930), .B0(net217968), .B1(n50455),
        .C0(net217016), .C1(n50454), .Y(n15029) );
  NOR2X1 U51529 ( .A(n29999), .B(n29998), .Y(net216258) );
  NOR4X1 U51530 ( .A(n29997), .B(n29996), .C(n29995), .D(n29994), .Y(net216259) );
  NOR2X1 U51531 ( .A(n30089), .B(n30088), .Y(net216285) );
  NOR4X1 U51532 ( .A(n30087), .B(n30086), .C(n30085), .D(n30084), .Y(net216286) );
  NOR2X1 U51533 ( .A(n30029), .B(n30028), .Y(net216267) );
  NOR4X1 U51534 ( .A(n30027), .B(n30026), .C(n30025), .D(n30024), .Y(net216268) );
  NAND4X1 U51535 ( .A(n44614), .B(n44613), .C(n44612), .D(n44611), .Y(n12169)
         );
  NOR2X1 U51536 ( .A(n29698), .B(n29697), .Y(n44612) );
  NOR4X1 U51537 ( .A(n29696), .B(n29695), .C(n29694), .D(n29693), .Y(n44611)
         );
  NOR2X1 U51538 ( .A(n26088), .B(n26087), .Y(net215071) );
  NOR4X1 U51539 ( .A(n26086), .B(n26085), .C(n26084), .D(n26083), .Y(net215072) );
  NAND4X1 U51540 ( .A(n43472), .B(n43471), .C(n43470), .D(n43469), .Y(n12802)
         );
  NOR2X1 U51541 ( .A(n30602), .B(n30601), .Y(n43470) );
  NOR4X1 U51542 ( .A(n30600), .B(n30599), .C(n30598), .D(n30597), .Y(n43469)
         );
  NAND4X1 U51543 ( .A(n43452), .B(n43451), .C(n43450), .D(n43449), .Y(n10483)
         );
  NOR2X1 U51544 ( .A(n30452), .B(n30451), .Y(n43450) );
  NOR4X1 U51545 ( .A(n30450), .B(n30449), .C(n30448), .D(n30447), .Y(n43449)
         );
  NOR4X1 U51546 ( .A(n30238), .B(n30237), .C(n30236), .D(n30235), .Y(net216358) );
  NOR2X1 U51547 ( .A(n26328), .B(n26327), .Y(net215125) );
  NOR4X1 U51548 ( .A(n26326), .B(n26325), .C(n26324), .D(n26323), .Y(net215126) );
  NAND4X1 U51549 ( .A(n43422), .B(n43421), .C(n43420), .D(n43419), .Y(n11954)
         );
  NOR2X1 U51550 ( .A(n30903), .B(n30902), .Y(n43420) );
  NOR4X1 U51551 ( .A(n30901), .B(n30900), .C(n30899), .D(n30898), .Y(n43419)
         );
  NOR2X1 U51552 ( .A(n30270), .B(n30269), .Y(net216366) );
  NOR4X1 U51553 ( .A(n30268), .B(n30267), .C(n30266), .D(n30265), .Y(net216367) );
  NOR2X1 U51554 ( .A(n26118), .B(n26117), .Y(net215080) );
  NOR4X1 U51555 ( .A(n26116), .B(n26115), .C(n26114), .D(n26113), .Y(net215081) );
  NOR4X1 U51556 ( .A(n24373), .B(n24372), .C(n24371), .D(n24370), .Y(net213525) );
  NOR4X1 U51557 ( .A(n24485), .B(n24484), .C(n24483), .D(n24482), .Y(net213570) );
  NAND4X1 U51558 ( .A(n47757), .B(n47756), .C(n47755), .D(n47754), .Y(n10801)
         );
  NOR2X1 U51559 ( .A(n22483), .B(n22482), .Y(n47755) );
  NOR4X1 U51560 ( .A(n22481), .B(n22480), .C(n22479), .D(n22478), .Y(n47754)
         );
  NOR2X1 U51561 ( .A(n30179), .B(n30178), .Y(net216312) );
  NOR4X1 U51562 ( .A(n30177), .B(n30176), .C(n30175), .D(n30174), .Y(net216313) );
  NOR2X1 U51563 ( .A(n24225), .B(n24224), .Y(net213464) );
  NOR2X1 U51564 ( .A(n20802), .B(n20801), .Y(net211581) );
  NOR4X1 U51565 ( .A(n20800), .B(n20799), .C(n20798), .D(n20797), .Y(net211582) );
  NOR2X1 U51566 ( .A(n30330), .B(n30329), .Y(net212156) );
  NOR4X1 U51567 ( .A(n30328), .B(n30327), .C(n30326), .D(n30325), .Y(net212157) );
  NOR4X1 U51568 ( .A(n24597), .B(n24596), .C(n24595), .D(n24594), .Y(net213626) );
  XNOR2X1 U51569 ( .A(n36734), .B(n32666), .Y(net212090) );
  NOR2X1 U51570 ( .A(n21872), .B(n21871), .Y(net212091) );
  NOR4X1 U51571 ( .A(n21870), .B(n21869), .C(n21868), .D(n21867), .Y(net212092) );
  NOR2X1 U51572 ( .A(n21264), .B(n21263), .Y(net211770) );
  NOR2X1 U51573 ( .A(n26358), .B(n26357), .Y(net215134) );
  NOR4X1 U51574 ( .A(n26356), .B(n26355), .C(n26354), .D(n26353), .Y(net215135) );
  NOR2X1 U51575 ( .A(n30059), .B(n30058), .Y(net216276) );
  NOR4X1 U51576 ( .A(n30057), .B(n30056), .C(n30055), .D(n30054), .Y(net216277) );
  NOR4X1 U51577 ( .A(n24495), .B(n24494), .C(n24493), .D(n24492), .Y(net213575) );
  NOR2X1 U51578 ( .A(n26058), .B(n26057), .Y(net215062) );
  NOR4X1 U51579 ( .A(n26056), .B(n26055), .C(n26054), .D(n26053), .Y(net215063) );
  NOR4X1 U51580 ( .A(n24556), .B(n24555), .C(n24554), .D(n24553), .Y(net213606) );
  NOR2X1 U51581 ( .A(n29969), .B(n29968), .Y(net216249) );
  NOR4X1 U51582 ( .A(n29967), .B(n29966), .C(n29965), .D(n29964), .Y(net216250) );
  NOR2X1 U51583 ( .A(n21284), .B(n21283), .Y(net211780) );
  NAND4X1 U51584 ( .A(n46632), .B(n46631), .C(n46630), .D(n46629), .Y(n10793)
         );
  NOR2X1 U51585 ( .A(n24387), .B(n24386), .Y(n46630) );
  NOR4X1 U51586 ( .A(n24385), .B(n24384), .C(n24383), .D(n24382), .Y(n46629)
         );
  XNOR2X1 U51587 ( .A(n36734), .B(n32682), .Y(net212074) );
  NOR2X1 U51588 ( .A(n21902), .B(n21901), .Y(net212075) );
  NOR4X1 U51589 ( .A(n21900), .B(n21899), .C(n21898), .D(n21897), .Y(net212076) );
  XNOR2X1 U51590 ( .A(n32994), .B(n42567), .Y(n43412) );
  NOR2X1 U51591 ( .A(n30813), .B(n30812), .Y(n43411) );
  NOR4X1 U51592 ( .A(n30811), .B(n30810), .C(n30809), .D(n30808), .Y(n43410)
         );
  NAND4BX1 U51593 ( .AN(n47952), .B(n49335), .C(n47951), .D(n9756), .Y(n34508)
         );
  NAND3X1 U51594 ( .A(n9773), .B(n9772), .C(n9771), .Y(n47951) );
  AOI31X1 U51595 ( .A0(n9757), .A1(n50105), .A2(n9759), .B0(n9760), .Y(n9756)
         );
  NOR4X1 U51596 ( .A(n24587), .B(n24586), .C(n24585), .D(n24584), .Y(net213621) );
  NOR4X1 U51597 ( .A(n24293), .B(n24292), .C(n24291), .D(n24290), .Y(net213450) );
  NOR4X1 U51598 ( .A(n24567), .B(n24566), .C(n24565), .D(n24564), .Y(net213611) );
  XNOR2X1 U51599 ( .A(n32397), .B(nxt_data_num[3]), .Y(n9695) );
  NOR2X1 U51600 ( .A(n20065), .B(n20064), .Y(net211450) );
  NOR2X1 U51601 ( .A(n21892), .B(n21891), .Y(net212101) );
  NOR4X1 U51602 ( .A(n24577), .B(n24576), .C(n24575), .D(n24574), .Y(net213616) );
  XNOR2X1 U51603 ( .A(n32399), .B(nxt_data_num[1]), .Y(n9697) );
  NAND4X1 U51604 ( .A(n47796), .B(n47795), .C(n47794), .D(n47793), .Y(n12238)
         );
  NOR2X1 U51605 ( .A(n22604), .B(n22603), .Y(n47794) );
  NOR4X1 U51606 ( .A(n22602), .B(n22601), .C(n22600), .D(n22599), .Y(n47793)
         );
  NAND4X1 U51607 ( .A(n46614), .B(n46613), .C(n46612), .D(n46611), .Y(n12228)
         );
  NOR2X1 U51608 ( .A(n24397), .B(n24396), .Y(n46612) );
  NOR4X1 U51609 ( .A(n24395), .B(n24394), .C(n24393), .D(n24392), .Y(n46611)
         );
  NOR2X1 U51610 ( .A(n24255), .B(n24254), .Y(net212024) );
  NOR4X1 U51611 ( .A(n24253), .B(n24252), .C(n24251), .D(n24250), .Y(net212025) );
  NAND4X1 U51612 ( .A(n47871), .B(n47870), .C(n47869), .D(n47868), .Y(n12186)
         );
  NOR2X1 U51613 ( .A(n23616), .B(n23615), .Y(n47869) );
  NOR4X1 U51614 ( .A(n23614), .B(n23613), .C(n23612), .D(n23611), .Y(n47868)
         );
  NOR2X1 U51615 ( .A(n26208), .B(n26207), .Y(net213222) );
  NOR4X1 U51616 ( .A(n26206), .B(n26205), .C(n26204), .D(n26203), .Y(net213223) );
  NOR4X1 U51617 ( .A(n23329), .B(n23328), .C(n23327), .D(n23326), .Y(net213239) );
  NAND4X1 U51618 ( .A(n46084), .B(n46083), .C(n46082), .D(n46081), .Y(n10906)
         );
  NOR2X1 U51619 ( .A(n22493), .B(n22492), .Y(n46082) );
  NOR4X1 U51620 ( .A(n22491), .B(n22490), .C(n22489), .D(n22488), .Y(n46081)
         );
  NOR2X1 U51621 ( .A(n25998), .B(n25997), .Y(net215044) );
  NOR4X1 U51622 ( .A(n25996), .B(n25995), .C(n25994), .D(n25993), .Y(net215045) );
  NAND4X1 U51623 ( .A(n45596), .B(n45595), .C(n45594), .D(n45593), .Y(n12213)
         );
  XNOR2X1 U51624 ( .A(n36837), .B(n32682), .Y(n45595) );
  NOR2X1 U51625 ( .A(n24335), .B(n24334), .Y(n45594) );
  NOR4X1 U51626 ( .A(n24333), .B(n24332), .C(n24331), .D(n24330), .Y(n45593)
         );
  NAND4X1 U51627 ( .A(n44334), .B(n44333), .C(n44332), .D(n44331), .Y(n10446)
         );
  NOR2X1 U51628 ( .A(n26479), .B(n26478), .Y(n44332) );
  NOR4X1 U51629 ( .A(n26477), .B(n26476), .C(n26475), .D(n26474), .Y(n44331)
         );
  NOR2X1 U51630 ( .A(n20908), .B(n20906), .Y(net211637) );
  OAI211X1 U51631 ( .A0(n34420), .A1(n42911), .B0(n13040), .C0(n50077), .Y(
        n34522) );
  OAI222XL U51632 ( .A0(net266654), .A1(n9670), .B0(n40159), .B1(n9669), .C0(
        n40292), .C1(n34428), .Y(n13042) );
  CLKINVX1 U51633 ( .A(n19167), .Y(n49562) );
  OAI222XL U51634 ( .A0(net266381), .A1(n9669), .B0(n40174), .B1(n34428), .C0(
        n40303), .C1(n34420), .Y(n19167) );
  AOI222XL U51635 ( .A0(net265302), .A1(n51438), .B0(net218034), .B1(n51437),
        .C0(net217108), .C1(n51436), .Y(n18206) );
  AOI222XL U51636 ( .A0(net265283), .A1(n51437), .B0(n40213), .B1(n51436),
        .C0(n40318), .C1(n51435), .Y(n18182) );
  AOI222XL U51637 ( .A0(net265283), .A1(n51436), .B0(n40236), .B1(n51435),
        .C0(n40318), .C1(n51434), .Y(n18158) );
  AOI222XL U51638 ( .A0(net265283), .A1(n51435), .B0(n40236), .B1(n51434),
        .C0(n40318), .C1(n51433), .Y(n18134) );
  AOI222XL U51639 ( .A0(net265264), .A1(n51434), .B0(n40236), .B1(n51433),
        .C0(n40319), .C1(n51432), .Y(n18110) );
  AOI222XL U51640 ( .A0(net265264), .A1(n51433), .B0(n40237), .B1(n51432),
        .C0(n40319), .C1(n51431), .Y(n18086) );
  OAI211X1 U51641 ( .A0(n34044), .A1(n42802), .B0(n18061), .C0(n18062), .Y(
        n36193) );
  OA22X1 U51642 ( .A0(net262912), .A1(n34028), .B0(n34036), .B1(n40101), .Y(
        n18061) );
  AOI222XL U51643 ( .A0(net265264), .A1(n51432), .B0(n40237), .B1(n51431),
        .C0(n40320), .C1(n51430), .Y(n18062) );
  OAI211X1 U51644 ( .A0(n34036), .A1(n42803), .B0(n18037), .C0(n18038), .Y(
        n36185) );
  OA22X1 U51645 ( .A0(net262912), .A1(n34020), .B0(n34028), .B1(n40101), .Y(
        n18037) );
  AOI222XL U51646 ( .A0(net265245), .A1(n51431), .B0(n40238), .B1(n51430),
        .C0(n40320), .C1(n51429), .Y(n18038) );
  AOI222XL U51647 ( .A0(net265245), .A1(n51430), .B0(n40238), .B1(n51429),
        .C0(n40320), .C1(n51428), .Y(n18014) );
  AOI222XL U51648 ( .A0(net265245), .A1(n51429), .B0(n40238), .B1(n51428),
        .C0(n40321), .C1(n51427), .Y(n17990) );
  AOI222XL U51649 ( .A0(net265226), .A1(n51428), .B0(n40239), .B1(n51427),
        .C0(n40321), .C1(n51426), .Y(n17966) );
  AOI222XL U51650 ( .A0(net265226), .A1(n51427), .B0(n40239), .B1(n51426),
        .C0(n40321), .C1(n51425), .Y(n17942) );
  AOI222XL U51651 ( .A0(net265226), .A1(n51426), .B0(n40240), .B1(n51425),
        .C0(n40322), .C1(n51424), .Y(n17918) );
  AOI222XL U51652 ( .A0(net265207), .A1(n51425), .B0(n40240), .B1(n51424),
        .C0(n40322), .C1(n51423), .Y(n17894) );
  AOI222XL U51653 ( .A0(net265207), .A1(n51424), .B0(n40240), .B1(n51423),
        .C0(n40322), .C1(n51422), .Y(n17870) );
  AOI222XL U51654 ( .A0(net265207), .A1(n51423), .B0(n40241), .B1(n51422),
        .C0(n40323), .C1(n51421), .Y(n17846) );
  OAI211X1 U51655 ( .A0(n33964), .A1(n42814), .B0(n17821), .C0(n17822), .Y(
        n36113) );
  AOI222XL U51656 ( .A0(net265188), .A1(n51422), .B0(n40241), .B1(n51421),
        .C0(n40323), .C1(n51420), .Y(n17822) );
  OAI211X1 U51657 ( .A0(n33956), .A1(n42847), .B0(n17797), .C0(n17798), .Y(
        n36105) );
  AOI222XL U51658 ( .A0(net265188), .A1(n51421), .B0(n40242), .B1(n51420),
        .C0(n40323), .C1(n51419), .Y(n17798) );
  AOI222XL U51659 ( .A0(net265188), .A1(n51420), .B0(n40242), .B1(n51419),
        .C0(n40324), .C1(n51418), .Y(n17774) );
  AOI222XL U51660 ( .A0(net265169), .A1(n51419), .B0(n40242), .B1(n51418),
        .C0(n40324), .C1(n51417), .Y(n17750) );
  AOI222XL U51661 ( .A0(net265169), .A1(n51418), .B0(n40243), .B1(n51417),
        .C0(n40324), .C1(n51416), .Y(n17726) );
  OAI211X1 U51662 ( .A0(n33924), .A1(n42852), .B0(n17701), .C0(n17702), .Y(
        n36073) );
  OA22X1 U51663 ( .A0(net262779), .A1(n33908), .B0(n33916), .B1(n40107), .Y(
        n17701) );
  AOI222XL U51664 ( .A0(net265169), .A1(n51417), .B0(n40243), .B1(n51416),
        .C0(n40325), .C1(n51415), .Y(n17702) );
  OAI211X1 U51665 ( .A0(n33916), .A1(n42853), .B0(n17677), .C0(n17678), .Y(
        n36065) );
  OA22X1 U51666 ( .A0(net262779), .A1(n33900), .B0(n33908), .B1(n40107), .Y(
        n17677) );
  AOI222XL U51667 ( .A0(net265150), .A1(n51416), .B0(n40244), .B1(n51415),
        .C0(n40325), .C1(n51414), .Y(n17678) );
  OAI211X1 U51668 ( .A0(n33908), .A1(n42854), .B0(n17653), .C0(n17654), .Y(
        n36057) );
  OA22X1 U51669 ( .A0(net262779), .A1(n33892), .B0(n33900), .B1(n40106), .Y(
        n17653) );
  AOI222XL U51670 ( .A0(net265150), .A1(n51415), .B0(n40244), .B1(n51414),
        .C0(n40348), .C1(n51413), .Y(n17654) );
  AOI222XL U51671 ( .A0(net265150), .A1(n51414), .B0(n40244), .B1(n51413),
        .C0(n40349), .C1(n51412), .Y(n17630) );
  AOI222XL U51672 ( .A0(net265131), .A1(n51413), .B0(n40245), .B1(n51412),
        .C0(net217092), .C1(n51411), .Y(n17606) );
  AOI222XL U51673 ( .A0(net265473), .A1(n51412), .B0(n40225), .B1(n51411),
        .C0(n40326), .C1(n51410), .Y(n17582) );
  AOI222XL U51674 ( .A0(net265454), .A1(n51411), .B0(n40225), .B1(n51410),
        .C0(n40326), .C1(n51409), .Y(n17558) );
  AOI222XL U51675 ( .A0(net265454), .A1(n51410), .B0(n40226), .B1(n51409),
        .C0(n40326), .C1(n51408), .Y(n17534) );
  AOI222XL U51676 ( .A0(net265454), .A1(n51409), .B0(n40226), .B1(n51408),
        .C0(n40327), .C1(n51407), .Y(n17510) );
  AOI222XL U51677 ( .A0(net265435), .A1(n51408), .B0(n40226), .B1(n51407),
        .C0(n40327), .C1(n51406), .Y(n17486) );
  AOI222XL U51678 ( .A0(net265435), .A1(n51407), .B0(n40227), .B1(n51406),
        .C0(n40327), .C1(n51405), .Y(n17462) );
  AOI222XL U51679 ( .A0(net265435), .A1(n51406), .B0(n40227), .B1(n51405),
        .C0(n40328), .C1(n51404), .Y(n17438) );
  AOI222XL U51680 ( .A0(net265416), .A1(n51405), .B0(n40228), .B1(n51404),
        .C0(n40328), .C1(n51403), .Y(n17414) );
  AOI222XL U51681 ( .A0(net265416), .A1(n51404), .B0(n40228), .B1(n51403),
        .C0(n40328), .C1(n51402), .Y(n17390) );
  AOI222XL U51682 ( .A0(net265416), .A1(n51403), .B0(n40228), .B1(n51402),
        .C0(n40329), .C1(n51401), .Y(n17366) );
  AOI222XL U51683 ( .A0(net265397), .A1(n51402), .B0(n40229), .B1(n51401),
        .C0(n40329), .C1(n51400), .Y(n17342) );
  AOI222XL U51684 ( .A0(net265397), .A1(n51401), .B0(n40229), .B1(n51400),
        .C0(n40329), .C1(n51399), .Y(n17318) );
  AOI222XL U51685 ( .A0(net265397), .A1(n51400), .B0(n40230), .B1(n51399),
        .C0(n40330), .C1(n51398), .Y(n17294) );
  AOI222XL U51686 ( .A0(net265378), .A1(n51399), .B0(n40230), .B1(n51398),
        .C0(n40330), .C1(n51397), .Y(n17270) );
  AOI222XL U51687 ( .A0(net265378), .A1(n51398), .B0(n40231), .B1(n51397),
        .C0(n40331), .C1(n51396), .Y(n17246) );
  AOI222XL U51688 ( .A0(net265378), .A1(n51397), .B0(n40231), .B1(n51396),
        .C0(n40331), .C1(n51395), .Y(n17222) );
  AOI222XL U51689 ( .A0(net265359), .A1(n51396), .B0(n40231), .B1(n51395),
        .C0(n40331), .C1(n51394), .Y(n17198) );
  AOI222XL U51690 ( .A0(net265359), .A1(n51395), .B0(n40232), .B1(n51394),
        .C0(n40332), .C1(n51393), .Y(n17174) );
  AOI222XL U51691 ( .A0(net265359), .A1(n51394), .B0(n40232), .B1(n51393),
        .C0(n40332), .C1(n51392), .Y(n17150) );
  AOI222XL U51692 ( .A0(net265340), .A1(n51393), .B0(n40233), .B1(n51392),
        .C0(n40332), .C1(n51391), .Y(n17126) );
  AOI222XL U51693 ( .A0(net265340), .A1(n51392), .B0(n40233), .B1(n51391),
        .C0(n40333), .C1(n51390), .Y(n17102) );
  AOI222XL U51694 ( .A0(net265340), .A1(n51391), .B0(n40233), .B1(n51390),
        .C0(n40333), .C1(n51389), .Y(n17078) );
  AOI222XL U51695 ( .A0(net265321), .A1(n51390), .B0(n40234), .B1(n51389),
        .C0(n40333), .C1(n51388), .Y(n17054) );
  OAI211X1 U51696 ( .A0(n33700), .A1(n42755), .B0(n17029), .C0(n17030), .Y(
        n35849) );
  AOI222XL U51697 ( .A0(net265321), .A1(n51389), .B0(n40234), .B1(n51388),
        .C0(n40334), .C1(n51387), .Y(n17030) );
  AOI222XL U51698 ( .A0(net265321), .A1(n51388), .B0(n40235), .B1(n51387),
        .C0(n40334), .C1(n51386), .Y(n17006) );
  AOI222XL U51699 ( .A0(net265302), .A1(n51387), .B0(n40235), .B1(n51386),
        .C0(n40334), .C1(n51385), .Y(n16982) );
  AOI222XL U51700 ( .A0(net265302), .A1(n51386), .B0(n40235), .B1(n51385),
        .C0(n40335), .C1(n51384), .Y(n16958) );
  AOI222XL U51701 ( .A0(net264960), .A1(n51385), .B0(n40256), .B1(n51384),
        .C0(n40335), .C1(n51383), .Y(n16934) );
  AOI222XL U51702 ( .A0(net264960), .A1(n51384), .B0(n40256), .B1(n51383),
        .C0(n40335), .C1(n51382), .Y(n16910) );
  OAI211X1 U51703 ( .A0(n33652), .A1(n42762), .B0(n16885), .C0(n16886), .Y(
        n35801) );
  OA22X1 U51704 ( .A0(net261981), .A1(n33636), .B0(n33644), .B1(n40144), .Y(
        n16885) );
  AOI222XL U51705 ( .A0(net264941), .A1(n51383), .B0(n40257), .B1(n51382),
        .C0(n40336), .C1(n51381), .Y(n16886) );
  AOI222XL U51706 ( .A0(net264941), .A1(n51382), .B0(n40257), .B1(n51381),
        .C0(n40336), .C1(n51380), .Y(n16862) );
  AOI222XL U51707 ( .A0(net264941), .A1(n51381), .B0(n40258), .B1(n51380),
        .C0(n40337), .C1(n51379), .Y(n16838) );
  AOI222XL U51708 ( .A0(net264922), .A1(n51380), .B0(n40258), .B1(n51379),
        .C0(n40337), .C1(n51378), .Y(n16814) );
  AOI222XL U51709 ( .A0(net264922), .A1(n51379), .B0(n40258), .B1(n51378),
        .C0(n40337), .C1(n51377), .Y(n16790) );
  AOI222XL U51710 ( .A0(net264922), .A1(n51378), .B0(n40259), .B1(n51377),
        .C0(n40338), .C1(n51376), .Y(n16766) );
  AOI222XL U51711 ( .A0(net264903), .A1(n51377), .B0(n40259), .B1(n51376),
        .C0(n40338), .C1(n51375), .Y(n16742) );
  AOI222XL U51712 ( .A0(net264903), .A1(n51376), .B0(n40260), .B1(n51375),
        .C0(n40338), .C1(n51374), .Y(n16718) );
  AOI222XL U51713 ( .A0(net264903), .A1(n51375), .B0(n40260), .B1(n51374),
        .C0(n40339), .C1(n51373), .Y(n16694) );
  AOI222XL U51714 ( .A0(net264884), .A1(n51374), .B0(n40260), .B1(n51373),
        .C0(n40339), .C1(n51372), .Y(n16670) );
  AOI222XL U51715 ( .A0(net264884), .A1(n51373), .B0(n40261), .B1(n51372),
        .C0(n40339), .C1(n51371), .Y(n16646) );
  AOI222XL U51716 ( .A0(net265207), .A1(n51372), .B0(n40266), .B1(n51371),
        .C0(n40340), .C1(n51370), .Y(n16622) );
  AOI222XL U51717 ( .A0(net264808), .A1(n51371), .B0(n40266), .B1(n51370),
        .C0(n40340), .C1(n51369), .Y(n16598) );
  OAI211X1 U51718 ( .A0(n33548), .A1(n42745), .B0(n16573), .C0(n16574), .Y(
        n35697) );
  OA22X1 U51719 ( .A0(net262361), .A1(n33532), .B0(n33540), .B1(n40125), .Y(
        n16573) );
  AOI222XL U51720 ( .A0(net264808), .A1(n51370), .B0(n40265), .B1(n51369),
        .C0(n40340), .C1(n51368), .Y(n16574) );
  OAI211X1 U51721 ( .A0(n33540), .A1(n42746), .B0(n16549), .C0(n16550), .Y(
        n35689) );
  OA22X1 U51722 ( .A0(net262361), .A1(n33524), .B0(n33532), .B1(n40124), .Y(
        n16549) );
  AOI222XL U51723 ( .A0(net264808), .A1(n51369), .B0(n40265), .B1(n51368),
        .C0(n40341), .C1(n51367), .Y(n16550) );
  OAI211X1 U51724 ( .A0(n33532), .A1(n42747), .B0(n16525), .C0(n16526), .Y(
        n35681) );
  OA22X1 U51725 ( .A0(net262380), .A1(n33516), .B0(n33524), .B1(n40124), .Y(
        n16525) );
  AOI222XL U51726 ( .A0(net264827), .A1(n51368), .B0(n40265), .B1(n51367),
        .C0(n40341), .C1(n51366), .Y(n16526) );
  OAI211X1 U51727 ( .A0(n33524), .A1(n42748), .B0(n16501), .C0(n16502), .Y(
        n35673) );
  OA22X1 U51728 ( .A0(net262380), .A1(n33508), .B0(n33516), .B1(n40123), .Y(
        n16501) );
  AOI222XL U51729 ( .A0(net264827), .A1(n51367), .B0(n40264), .B1(n51366),
        .C0(n40341), .C1(n51365), .Y(n16502) );
  AOI222XL U51730 ( .A0(net264827), .A1(n51366), .B0(n40264), .B1(n51365),
        .C0(n40342), .C1(n51364), .Y(n16478) );
  AOI222XL U51731 ( .A0(net264846), .A1(n51365), .B0(n40263), .B1(n51364),
        .C0(n40342), .C1(n51363), .Y(n16454) );
  AOI222XL U51732 ( .A0(net264846), .A1(n51364), .B0(n40263), .B1(n51363),
        .C0(n40343), .C1(n51362), .Y(n16430) );
  AOI222XL U51733 ( .A0(net264846), .A1(n51363), .B0(n40263), .B1(n51362),
        .C0(n40343), .C1(n51361), .Y(n16406) );
  AOI222XL U51734 ( .A0(net264865), .A1(n51362), .B0(n40262), .B1(n51361),
        .C0(n40343), .C1(n51360), .Y(n16382) );
  AOI222XL U51735 ( .A0(net264865), .A1(n51361), .B0(n40262), .B1(n51360),
        .C0(n40344), .C1(n51359), .Y(n16358) );
  AOI222XL U51736 ( .A0(net264865), .A1(n51360), .B0(n40261), .B1(n51359),
        .C0(n40344), .C1(n51358), .Y(n16334) );
  OAI211X1 U51737 ( .A0(n33460), .A1(n42789), .B0(n16309), .C0(n16310), .Y(
        n35609) );
  AOI222XL U51738 ( .A0(net265036), .A1(n51359), .B0(n40245), .B1(n51358),
        .C0(n40344), .C1(n51357), .Y(n16310) );
  OAI211X1 U51739 ( .A0(n33452), .A1(n42791), .B0(n16285), .C0(n16286), .Y(
        n35601) );
  AOI222XL U51740 ( .A0(net265131), .A1(n51358), .B0(n40246), .B1(n51357),
        .C0(n40345), .C1(n51356), .Y(n16286) );
  OAI211X1 U51741 ( .A0(n33444), .A1(n42792), .B0(n16261), .C0(n16262), .Y(
        n35593) );
  AOI222XL U51742 ( .A0(net265112), .A1(n51357), .B0(n40246), .B1(n51356),
        .C0(n40345), .C1(n51355), .Y(n16262) );
  AOI222XL U51743 ( .A0(net265112), .A1(n51356), .B0(n40246), .B1(n51355),
        .C0(n40345), .C1(n51354), .Y(n16238) );
  OAI211X1 U51744 ( .A0(n33428), .A1(n42794), .B0(n16213), .C0(n16214), .Y(
        n35577) );
  OA22X1 U51745 ( .A0(net262209), .A1(n33412), .B0(n33420), .B1(n40132), .Y(
        n16213) );
  AOI222XL U51746 ( .A0(net265112), .A1(n51355), .B0(n40247), .B1(n51354),
        .C0(n40346), .C1(n51353), .Y(n16214) );
  OAI211X1 U51747 ( .A0(n33420), .A1(n42795), .B0(n16189), .C0(n16190), .Y(
        n35569) );
  OA22X1 U51748 ( .A0(net262228), .A1(n33404), .B0(n33412), .B1(n40132), .Y(
        n16189) );
  AOI222XL U51749 ( .A0(net221814), .A1(n51354), .B0(n40247), .B1(n51353),
        .C0(n40346), .C1(n51352), .Y(n16190) );
  OAI211X1 U51750 ( .A0(n33412), .A1(n42796), .B0(n16165), .C0(n16166), .Y(
        n35561) );
  OA22X1 U51751 ( .A0(net262228), .A1(n33396), .B0(n33404), .B1(n40131), .Y(
        n16165) );
  AOI222XL U51752 ( .A0(net221808), .A1(n51353), .B0(n40248), .B1(n51352),
        .C0(n40346), .C1(n51351), .Y(n16166) );
  OAI211X1 U51753 ( .A0(n33404), .A1(n42797), .B0(n16141), .C0(n16142), .Y(
        n35553) );
  OA22X1 U51754 ( .A0(net262247), .A1(n33388), .B0(n33396), .B1(n40131), .Y(
        n16141) );
  AOI222XL U51755 ( .A0(net221818), .A1(n51352), .B0(n40248), .B1(n51351),
        .C0(n40347), .C1(n51350), .Y(n16142) );
  OAI211X1 U51756 ( .A0(n33396), .A1(n42774), .B0(n16117), .C0(n16118), .Y(
        n35545) );
  OA22X1 U51757 ( .A0(net262247), .A1(n33380), .B0(n33388), .B1(n40130), .Y(
        n16117) );
  AOI222XL U51758 ( .A0(net265074), .A1(n51351), .B0(n40248), .B1(n51350),
        .C0(n40347), .C1(n51349), .Y(n16118) );
  AOI222XL U51759 ( .A0(net265074), .A1(n51350), .B0(n40249), .B1(n51349),
        .C0(n40347), .C1(n51348), .Y(n16094) );
  AOI222XL U51760 ( .A0(net265074), .A1(n51349), .B0(n40249), .B1(n51348),
        .C0(n40348), .C1(n51347), .Y(n16070) );
  AOI222XL U51761 ( .A0(net265055), .A1(n51348), .B0(n40250), .B1(n51347),
        .C0(n40348), .C1(n51346), .Y(n16046) );
  AOI222XL U51762 ( .A0(net265055), .A1(n51347), .B0(n40250), .B1(n51346),
        .C0(n40349), .C1(n51345), .Y(n16022) );
  AOI222XL U51763 ( .A0(net265055), .A1(n51346), .B0(n40250), .B1(n51345),
        .C0(n40349), .C1(n51344), .Y(n15998) );
  AOI222XL U51764 ( .A0(net265036), .A1(n51345), .B0(n40251), .B1(n51344),
        .C0(n40349), .C1(n51343), .Y(n15974) );
  AOI222XL U51765 ( .A0(net265036), .A1(n51344), .B0(n40251), .B1(n51343),
        .C0(n40382), .C1(n51342), .Y(n15950) );
  AOI222XL U51766 ( .A0(net265036), .A1(n51343), .B0(n40252), .B1(n51342),
        .C0(n40382), .C1(n51341), .Y(n15926) );
  AOI222XL U51767 ( .A0(net265017), .A1(n51342), .B0(n40252), .B1(n51341),
        .C0(n40382), .C1(n51340), .Y(n15902) );
  AOI222XL U51768 ( .A0(net265017), .A1(n51341), .B0(n40252), .B1(n51340),
        .C0(n40350), .C1(n51339), .Y(n15878) );
  AOI222XL U51769 ( .A0(net265017), .A1(n51340), .B0(n40253), .B1(n51339),
        .C0(n40350), .C1(n51338), .Y(n15854) );
  AOI222XL U51770 ( .A0(net264998), .A1(n51339), .B0(n40253), .B1(n51338),
        .C0(n40350), .C1(n51337), .Y(n15830) );
  AOI222XL U51771 ( .A0(net264998), .A1(n51338), .B0(n40254), .B1(n51337),
        .C0(net217036), .C1(n51336), .Y(n15806) );
  OAI211X1 U51772 ( .A0(n33284), .A1(n42782), .B0(n15781), .C0(n15782), .Y(
        n35433) );
  OA22X1 U51773 ( .A0(net263710), .A1(n33268), .B0(n33276), .B1(n40056), .Y(
        n15781) );
  AOI222XL U51774 ( .A0(net264998), .A1(n51337), .B0(n40254), .B1(n51336),
        .C0(n40346), .C1(n51335), .Y(n15782) );
  OAI211X1 U51775 ( .A0(n33276), .A1(n42944), .B0(n15757), .C0(n15758), .Y(
        n35425) );
  OA22X1 U51776 ( .A0(net263064), .A1(n33260), .B0(n33268), .B1(n40055), .Y(
        n15757) );
  AOI222XL U51777 ( .A0(net264979), .A1(n51336), .B0(n40254), .B1(n51335),
        .C0(n40343), .C1(n51334), .Y(n15758) );
  OAI211X1 U51778 ( .A0(n33268), .A1(n42945), .B0(n15733), .C0(n15734), .Y(
        n35417) );
  OA22X1 U51779 ( .A0(net263976), .A1(n33252), .B0(n33260), .B1(n40055), .Y(
        n15733) );
  AOI222XL U51780 ( .A0(net264979), .A1(n51335), .B0(n40255), .B1(n51334),
        .C0(n40351), .C1(n51333), .Y(n15734) );
  AOI222XL U51781 ( .A0(net264979), .A1(n51334), .B0(n40255), .B1(n51333),
        .C0(n40351), .C1(n51332), .Y(n15710) );
  AOI222XL U51782 ( .A0(net264960), .A1(n51333), .B0(n40256), .B1(n51332),
        .C0(n40351), .C1(n51331), .Y(n15686) );
  AOI222XL U51783 ( .A0(net265967), .A1(n51332), .B0(n40193), .B1(n51331),
        .C0(n40352), .C1(n51330), .Y(n15662) );
  AOI222XL U51784 ( .A0(net265967), .A1(n51331), .B0(n40193), .B1(n51330),
        .C0(n40352), .C1(n51329), .Y(n15638) );
  AOI222XL U51785 ( .A0(net265967), .A1(n51330), .B0(n40194), .B1(n51329),
        .C0(n40353), .C1(n51328), .Y(n15614) );
  AOI222XL U51786 ( .A0(net265948), .A1(n51329), .B0(n40194), .B1(n51328),
        .C0(n40353), .C1(n51327), .Y(n15590) );
  AOI222XL U51787 ( .A0(net265948), .A1(n51328), .B0(n40194), .B1(n51327),
        .C0(n40353), .C1(n51326), .Y(n15566) );
  AOI222XL U51788 ( .A0(net265948), .A1(n51327), .B0(n40195), .B1(n51326),
        .C0(n40354), .C1(n51325), .Y(n15542) );
  AOI222XL U51789 ( .A0(net265929), .A1(n51326), .B0(n40195), .B1(n51325),
        .C0(n40354), .C1(n51324), .Y(n15518) );
  AOI222XL U51790 ( .A0(net265929), .A1(n51325), .B0(n40196), .B1(n51324),
        .C0(n40354), .C1(n51323), .Y(n15494) );
  AOI222XL U51791 ( .A0(net265929), .A1(n51324), .B0(n40196), .B1(n51323),
        .C0(n40355), .C1(n51322), .Y(n15470) );
  AOI222XL U51792 ( .A0(net265910), .A1(n51323), .B0(n40196), .B1(n51322),
        .C0(n40355), .C1(n51321), .Y(n15446) );
  OAI211X1 U51793 ( .A0(n33164), .A1(n42928), .B0(n15421), .C0(n15422), .Y(
        n35313) );
  OA22X1 U51794 ( .A0(net263577), .A1(n33148), .B0(n33156), .B1(n40063), .Y(
        n15421) );
  AOI222XL U51795 ( .A0(net265910), .A1(n51322), .B0(n40197), .B1(n51321),
        .C0(n40355), .C1(n51320), .Y(n15422) );
  OAI211X1 U51796 ( .A0(n33156), .A1(n42929), .B0(n15397), .C0(n15398), .Y(
        n35305) );
  OA22X1 U51797 ( .A0(net263577), .A1(n33140), .B0(n33148), .B1(n40062), .Y(
        n15397) );
  AOI222XL U51798 ( .A0(net265910), .A1(n51321), .B0(n40197), .B1(n51320),
        .C0(n40356), .C1(n51319), .Y(n15398) );
  OAI211X1 U51799 ( .A0(n33148), .A1(n42930), .B0(n15373), .C0(n15374), .Y(
        n35297) );
  OA22X1 U51800 ( .A0(net263596), .A1(n33132), .B0(n33140), .B1(n40062), .Y(
        n15373) );
  AOI222XL U51801 ( .A0(net265891), .A1(n51320), .B0(n40198), .B1(n51319),
        .C0(n40356), .C1(n51318), .Y(n15374) );
  OAI211X1 U51802 ( .A0(n33140), .A1(n42932), .B0(n15349), .C0(n15350), .Y(
        n35289) );
  OA22X1 U51803 ( .A0(net263596), .A1(n33124), .B0(n33132), .B1(n40061), .Y(
        n15349) );
  AOI222XL U51804 ( .A0(net265891), .A1(n51319), .B0(n40198), .B1(n51318),
        .C0(n40356), .C1(n51317), .Y(n15350) );
  AOI222XL U51805 ( .A0(net265891), .A1(n51318), .B0(n40199), .B1(n51317),
        .C0(n40357), .C1(n51316), .Y(n15326) );
  AOI222XL U51806 ( .A0(net265872), .A1(n51317), .B0(n40199), .B1(n51316),
        .C0(n40357), .C1(n51315), .Y(n15302) );
  AOI222XL U51807 ( .A0(net265872), .A1(n51316), .B0(n40199), .B1(n51315),
        .C0(n40357), .C1(n51314), .Y(n15278) );
  AOI222XL U51808 ( .A0(net265872), .A1(n51315), .B0(n40200), .B1(n51314),
        .C0(n40358), .C1(n51313), .Y(n15254) );
  AOI222XL U51809 ( .A0(net265853), .A1(n51314), .B0(n40200), .B1(n51313),
        .C0(n40358), .C1(n51312), .Y(n15230) );
  AOI222XL U51810 ( .A0(net265853), .A1(n51313), .B0(n40201), .B1(n51312),
        .C0(n40359), .C1(n51311), .Y(n15206) );
  AOI222XL U51811 ( .A0(net265853), .A1(n51312), .B0(n40201), .B1(n51311),
        .C0(n40359), .C1(n51310), .Y(n15182) );
  AOI222XL U51812 ( .A0(net265834), .A1(n51311), .B0(n40201), .B1(n51310),
        .C0(n40359), .C1(n51309), .Y(n15158) );
  AOI222XL U51813 ( .A0(net265834), .A1(n51310), .B0(n40202), .B1(n51309),
        .C0(n40360), .C1(n51308), .Y(n15134) );
  AOI222XL U51814 ( .A0(net265834), .A1(n51309), .B0(n40202), .B1(n51308),
        .C0(n40360), .C1(n51307), .Y(n15110) );
  AOI222XL U51815 ( .A0(net265815), .A1(n51308), .B0(n40203), .B1(n51307),
        .C0(n40360), .C1(n51306), .Y(n15086) );
  AOI222XL U51816 ( .A0(net265815), .A1(n51307), .B0(n40203), .B1(n51306),
        .C0(net217018), .C1(n37242), .Y(n15062) );
  AOI222XL U51817 ( .A0(net265815), .A1(n51306), .B0(n40203), .B1(n37242),
        .C0(n40357), .C1(n51305), .Y(n15038) );
  AOI222XL U51818 ( .A0(net221892), .A1(n37242), .B0(net217954), .B1(n51305),
        .C0(net217020), .C1(n51304), .Y(n15014) );
  AOI222XL U51819 ( .A0(net221892), .A1(n51305), .B0(n40184), .B1(n51304),
        .C0(n40361), .C1(n51303), .Y(n14990) );
  OAI211X1 U51820 ( .A0(n33012), .A1(n42982), .B0(n14965), .C0(n14966), .Y(
        n35161) );
  OA22X1 U51821 ( .A0(net263995), .A1(n32996), .B0(n33004), .B1(net218866),
        .Y(n14965) );
  AOI222XL U51822 ( .A0(net221892), .A1(n51304), .B0(n40184), .B1(n51303),
        .C0(n40361), .C1(n51302), .Y(n14966) );
  AOI222XL U51823 ( .A0(net266119), .A1(n51303), .B0(n40185), .B1(n51302),
        .C0(n40361), .C1(n51301), .Y(n14942) );
  AOI222XL U51824 ( .A0(net266119), .A1(n51302), .B0(n40185), .B1(n51301),
        .C0(n40362), .C1(n51300), .Y(n14918) );
  AOI222XL U51825 ( .A0(net266119), .A1(n51301), .B0(n40185), .B1(n51300),
        .C0(n40362), .C1(n51299), .Y(n14894) );
  AOI222XL U51826 ( .A0(net266100), .A1(n51300), .B0(n40197), .B1(n51299),
        .C0(n40362), .C1(n51298), .Y(n14870) );
  AOI222XL U51827 ( .A0(net266100), .A1(n51299), .B0(n40197), .B1(n51298),
        .C0(n40363), .C1(n51297), .Y(n14846) );
  AOI222XL U51828 ( .A0(net266100), .A1(n51298), .B0(n40186), .B1(n51297),
        .C0(n40363), .C1(n51296), .Y(n14822) );
  OA22X1 U51829 ( .A0(net218474), .A1(n32940), .B0(n32948), .B1(n40051), .Y(
        n14797) );
  AOI222XL U51830 ( .A0(net266081), .A1(n51297), .B0(n40186), .B1(n51296),
        .C0(net217000), .C1(n51295), .Y(n14798) );
  OAI211X1 U51831 ( .A0(n32940), .A1(n42960), .B0(n14749), .C0(n14750), .Y(
        n35089) );
  AOI222XL U51832 ( .A0(net266081), .A1(n51295), .B0(n40187), .B1(n51294),
        .C0(n40372), .C1(n51293), .Y(n14750) );
  OAI211X1 U51833 ( .A0(n32932), .A1(n42961), .B0(n14725), .C0(n14726), .Y(
        n35081) );
  AOI222XL U51834 ( .A0(net266062), .A1(n51294), .B0(n40187), .B1(n51293),
        .C0(n40364), .C1(n51292), .Y(n14726) );
  OAI211X1 U51835 ( .A0(n32924), .A1(n42963), .B0(n14701), .C0(n14702), .Y(
        n35073) );
  AOI222XL U51836 ( .A0(net266062), .A1(n51293), .B0(n40188), .B1(n51292),
        .C0(n40364), .C1(n51291), .Y(n14702) );
  OA22X1 U51837 ( .A0(net263843), .A1(n32900), .B0(n32908), .B1(n40048), .Y(
        n14677) );
  AOI222XL U51838 ( .A0(net266043), .A1(n51292), .B0(n40188), .B1(n51291),
        .C0(n40364), .C1(n51290), .Y(n14678) );
  OAI211X1 U51839 ( .A0(n32908), .A1(n42965), .B0(n14653), .C0(n14654), .Y(
        n35057) );
  OA22X1 U51840 ( .A0(net263843), .A1(n32892), .B0(n32900), .B1(n40048), .Y(
        n14653) );
  AOI222XL U51841 ( .A0(net266043), .A1(n51291), .B0(n40188), .B1(n51290),
        .C0(n40365), .C1(n51289), .Y(n14654) );
  OAI211X1 U51842 ( .A0(n32900), .A1(n42966), .B0(n14629), .C0(n14630), .Y(
        n35049) );
  OA22X1 U51843 ( .A0(net263843), .A1(n32884), .B0(n32892), .B1(n40047), .Y(
        n14629) );
  AOI222XL U51844 ( .A0(net266043), .A1(n51290), .B0(n40189), .B1(n51289),
        .C0(n40365), .C1(n51288), .Y(n14630) );
  OAI211X1 U51845 ( .A0(n32892), .A1(n42967), .B0(n14605), .C0(n14606), .Y(
        n35041) );
  OA22X1 U51846 ( .A0(net263862), .A1(n32876), .B0(n32884), .B1(n40047), .Y(
        n14605) );
  AOI222XL U51847 ( .A0(net266024), .A1(n51289), .B0(n40189), .B1(n51288),
        .C0(n40365), .C1(n51287), .Y(n14606) );
  OAI211X1 U51848 ( .A0(n32884), .A1(n42968), .B0(n14581), .C0(n14582), .Y(
        n35033) );
  OA22X1 U51849 ( .A0(net263862), .A1(n32868), .B0(n32876), .B1(n40046), .Y(
        n14581) );
  AOI222XL U51850 ( .A0(net266024), .A1(n51288), .B0(n40190), .B1(n51287),
        .C0(n40366), .C1(n51286), .Y(n14582) );
  OA22X1 U51851 ( .A0(net263064), .A1(n32860), .B0(n32868), .B1(n40092), .Y(
        n14557) );
  AOI222XL U51852 ( .A0(net266024), .A1(n51287), .B0(n40190), .B1(n51286),
        .C0(n40366), .C1(n51285), .Y(n14558) );
  OA22X1 U51853 ( .A0(net263064), .A1(n32852), .B0(n32860), .B1(n40092), .Y(
        n14533) );
  AOI222XL U51854 ( .A0(net266005), .A1(n51286), .B0(n40190), .B1(n51285),
        .C0(n40366), .C1(n51284), .Y(n14534) );
  OA22X1 U51855 ( .A0(net263083), .A1(n32844), .B0(n32852), .B1(n40091), .Y(
        n14509) );
  AOI222XL U51856 ( .A0(net266005), .A1(n51285), .B0(n40191), .B1(n51284),
        .C0(n40367), .C1(n51283), .Y(n14510) );
  OAI211X1 U51857 ( .A0(n32852), .A1(n42973), .B0(n14485), .C0(n14486), .Y(
        n35001) );
  OA22X1 U51858 ( .A0(net263083), .A1(n32836), .B0(n32844), .B1(n40091), .Y(
        n14485) );
  AOI222XL U51859 ( .A0(net266005), .A1(n51284), .B0(n40191), .B1(n51283),
        .C0(n40367), .C1(n51282), .Y(n14486) );
  OAI211X1 U51860 ( .A0(n32844), .A1(n42974), .B0(n14461), .C0(n14462), .Y(
        n34993) );
  OA22X1 U51861 ( .A0(net263102), .A1(n32828), .B0(n32836), .B1(n40090), .Y(
        n14461) );
  AOI222XL U51862 ( .A0(net265511), .A1(n51283), .B0(n40192), .B1(n51282),
        .C0(n40367), .C1(n51281), .Y(n14462) );
  OAI211X1 U51863 ( .A0(n32836), .A1(n42975), .B0(n14437), .C0(n14438), .Y(
        n34985) );
  OA22X1 U51864 ( .A0(net263102), .A1(n32820), .B0(n32828), .B1(n40090), .Y(
        n14437) );
  AOI222XL U51865 ( .A0(net265606), .A1(n51282), .B0(n40192), .B1(n51281),
        .C0(n40368), .C1(n51280), .Y(n14438) );
  OAI211X1 U51866 ( .A0(n32828), .A1(n42879), .B0(n14413), .C0(n14414), .Y(
        n34977) );
  OA22X1 U51867 ( .A0(net263121), .A1(n32812), .B0(n32820), .B1(n40089), .Y(
        n14413) );
  AOI222XL U51868 ( .A0(net265625), .A1(n51281), .B0(n40192), .B1(n51280),
        .C0(n40368), .C1(n51279), .Y(n14414) );
  OAI211X1 U51869 ( .A0(n32820), .A1(n42880), .B0(n14389), .C0(n14390), .Y(
        n34969) );
  OA22X1 U51870 ( .A0(net263121), .A1(n32804), .B0(n32812), .B1(n40089), .Y(
        n14389) );
  AOI222XL U51871 ( .A0(net266062), .A1(n51280), .B0(n40214), .B1(n51279),
        .C0(n40369), .C1(n51278), .Y(n14390) );
  OAI211X1 U51872 ( .A0(n32812), .A1(n42882), .B0(n14365), .C0(n14366), .Y(
        n34961) );
  OA22X1 U51873 ( .A0(net263140), .A1(n32796), .B0(n32804), .B1(n40088), .Y(
        n14365) );
  AOI222XL U51874 ( .A0(net265625), .A1(n51279), .B0(n40214), .B1(n51278),
        .C0(n40369), .C1(n51277), .Y(n14366) );
  AOI222XL U51875 ( .A0(net265625), .A1(n51278), .B0(n40215), .B1(n51277),
        .C0(n40369), .C1(n51276), .Y(n14342) );
  AOI222XL U51876 ( .A0(net265625), .A1(n51277), .B0(n40215), .B1(n51276),
        .C0(n40370), .C1(n51275), .Y(n14318) );
  OA22X1 U51877 ( .A0(net263159), .A1(n32772), .B0(n32780), .B1(n40086), .Y(
        n14293) );
  AOI222XL U51878 ( .A0(net265606), .A1(n51276), .B0(n40216), .B1(n51275),
        .C0(n40370), .C1(n51274), .Y(n14294) );
  OA22X1 U51879 ( .A0(net263159), .A1(n32764), .B0(n32772), .B1(n40086), .Y(
        n14269) );
  AOI222XL U51880 ( .A0(net265606), .A1(n51275), .B0(n40216), .B1(n51274),
        .C0(n40370), .C1(n51273), .Y(n14270) );
  OAI211X1 U51881 ( .A0(n32772), .A1(n42887), .B0(n14245), .C0(n14246), .Y(
        n34921) );
  OA22X1 U51882 ( .A0(net263178), .A1(n32756), .B0(n32764), .B1(n40085), .Y(
        n14245) );
  AOI222XL U51883 ( .A0(net265606), .A1(n51274), .B0(n40216), .B1(n51273),
        .C0(n40371), .C1(n51272), .Y(n14246) );
  OAI211X1 U51884 ( .A0(n32764), .A1(n42889), .B0(n14221), .C0(n14222), .Y(
        n34913) );
  OA22X1 U51885 ( .A0(net263178), .A1(n32748), .B0(n32756), .B1(n40085), .Y(
        n14221) );
  AOI222XL U51886 ( .A0(net265587), .A1(n51273), .B0(n40217), .B1(n51272),
        .C0(n40371), .C1(n51271), .Y(n14222) );
  OAI211X1 U51887 ( .A0(n32756), .A1(n42890), .B0(n14197), .C0(n14198), .Y(
        n34905) );
  OA22X1 U51888 ( .A0(net261924), .A1(n32740), .B0(n32748), .B1(n40084), .Y(
        n14197) );
  AOI222XL U51889 ( .A0(net265587), .A1(n51272), .B0(n40217), .B1(n51271),
        .C0(n40371), .C1(n51270), .Y(n14198) );
  OAI211X1 U51890 ( .A0(n32748), .A1(n42891), .B0(n14173), .C0(n14174), .Y(
        n34897) );
  OA22X1 U51891 ( .A0(net262931), .A1(n32732), .B0(n32740), .B1(n40100), .Y(
        n14173) );
  AOI222XL U51892 ( .A0(net265587), .A1(n51271), .B0(n40218), .B1(n51270),
        .C0(n40372), .C1(n51269), .Y(n14174) );
  OA22X1 U51893 ( .A0(net262931), .A1(n32724), .B0(n32732), .B1(n40099), .Y(
        n14149) );
  AOI222XL U51894 ( .A0(net265568), .A1(n51270), .B0(n40218), .B1(n51269),
        .C0(n40372), .C1(n51268), .Y(n14150) );
  OA22X1 U51895 ( .A0(net262950), .A1(n32716), .B0(n32724), .B1(n40099), .Y(
        n14125) );
  AOI222XL U51896 ( .A0(net265568), .A1(n51269), .B0(n40218), .B1(n51268),
        .C0(n40372), .C1(n51267), .Y(n14126) );
  OA22X1 U51897 ( .A0(net262950), .A1(n32708), .B0(n32716), .B1(n40098), .Y(
        n14101) );
  AOI222XL U51898 ( .A0(net265568), .A1(n51268), .B0(n40219), .B1(n51267),
        .C0(n40373), .C1(n51266), .Y(n14102) );
  AOI222XL U51899 ( .A0(net265549), .A1(n51267), .B0(n40219), .B1(n51266),
        .C0(n40373), .C1(n51265), .Y(n14078) );
  AOI222XL U51900 ( .A0(net265549), .A1(n51266), .B0(n40220), .B1(n51265),
        .C0(n40373), .C1(n51264), .Y(n14054) );
  OA22X1 U51901 ( .A0(net262988), .A1(n32684), .B0(n32692), .B1(n40097), .Y(
        n14029) );
  AOI222XL U51902 ( .A0(net265549), .A1(n51265), .B0(n40220), .B1(n51264),
        .C0(n40374), .C1(n51263), .Y(n14030) );
  OA22X1 U51903 ( .A0(net262988), .A1(n32676), .B0(n32684), .B1(n40096), .Y(
        n14005) );
  AOI222XL U51904 ( .A0(net265530), .A1(n51264), .B0(n40221), .B1(n51263),
        .C0(n40374), .C1(n51262), .Y(n14006) );
  OAI211X1 U51905 ( .A0(n32684), .A1(n42868), .B0(n13981), .C0(n13982), .Y(
        n34833) );
  AOI222XL U51906 ( .A0(net265530), .A1(n51263), .B0(n40221), .B1(n51262),
        .C0(n40375), .C1(n51261), .Y(n13982) );
  OAI211X1 U51907 ( .A0(n32676), .A1(n42869), .B0(n13957), .C0(n13958), .Y(
        n34825) );
  AOI222XL U51908 ( .A0(net265530), .A1(n51262), .B0(n40221), .B1(n51261),
        .C0(n40375), .C1(n51260), .Y(n13958) );
  OAI211X1 U51909 ( .A0(n32668), .A1(n42870), .B0(n13933), .C0(n13934), .Y(
        n34817) );
  AOI222XL U51910 ( .A0(net265511), .A1(n51261), .B0(n40222), .B1(n51260),
        .C0(n40375), .C1(n51259), .Y(n13934) );
  OA22X1 U51911 ( .A0(net263026), .A1(n32644), .B0(n32652), .B1(n40094), .Y(
        n13909) );
  AOI222XL U51912 ( .A0(net265511), .A1(n51260), .B0(n40222), .B1(n51259),
        .C0(n40376), .C1(n51258), .Y(n13910) );
  OAI211X1 U51913 ( .A0(n32652), .A1(n42873), .B0(n13885), .C0(n13886), .Y(
        n34801) );
  OA22X1 U51914 ( .A0(net263026), .A1(n32636), .B0(n32644), .B1(n40094), .Y(
        n13885) );
  AOI222XL U51915 ( .A0(net265511), .A1(n51259), .B0(n40223), .B1(n51258),
        .C0(n40376), .C1(n51257), .Y(n13886) );
  OAI211X1 U51916 ( .A0(n32644), .A1(n42874), .B0(n13861), .C0(n13862), .Y(
        n34793) );
  OA22X1 U51917 ( .A0(net263045), .A1(n32628), .B0(n32636), .B1(n40093), .Y(
        n13861) );
  AOI222XL U51918 ( .A0(net265492), .A1(n51258), .B0(n40223), .B1(n51257),
        .C0(n40376), .C1(n51256), .Y(n13862) );
  OAI211X1 U51919 ( .A0(n32636), .A1(n42875), .B0(n13837), .C0(n13838), .Y(
        n34785) );
  OA22X1 U51920 ( .A0(net263045), .A1(n32620), .B0(n32628), .B1(n40093), .Y(
        n13837) );
  AOI222XL U51921 ( .A0(net265492), .A1(n51257), .B0(n40223), .B1(n51256),
        .C0(n40377), .C1(n51255), .Y(n13838) );
  OAI211X1 U51922 ( .A0(n32628), .A1(n42876), .B0(n13813), .C0(n13814), .Y(
        n34777) );
  OA22X1 U51923 ( .A0(net263064), .A1(n32612), .B0(n32620), .B1(n40092), .Y(
        n13813) );
  AOI222XL U51924 ( .A0(net265492), .A1(n51256), .B0(n40224), .B1(n51255),
        .C0(n40377), .C1(n51254), .Y(n13814) );
  OA22X1 U51925 ( .A0(net263330), .A1(n32604), .B0(n32612), .B1(n40077), .Y(
        n13789) );
  AOI222XL U51926 ( .A0(net265473), .A1(n51255), .B0(n40224), .B1(n51254),
        .C0(n40377), .C1(n51253), .Y(n13790) );
  OAI211X1 U51927 ( .A0(n32612), .A1(n42878), .B0(n13765), .C0(n13766), .Y(
        n34761) );
  OA22X1 U51928 ( .A0(net263349), .A1(n32596), .B0(n32604), .B1(n40076), .Y(
        n13765) );
  AOI222XL U51929 ( .A0(net265473), .A1(n51254), .B0(n40225), .B1(n51253),
        .C0(n40378), .C1(n51252), .Y(n13766) );
  OA22X1 U51930 ( .A0(net263349), .A1(n32588), .B0(n32596), .B1(n40076), .Y(
        n13741) );
  AOI222XL U51931 ( .A0(net265815), .A1(n51253), .B0(n40204), .B1(n51252),
        .C0(n40378), .C1(n51251), .Y(n13742) );
  OA22X1 U51932 ( .A0(net263368), .A1(n32580), .B0(n32588), .B1(n40075), .Y(
        n13717) );
  AOI222XL U51933 ( .A0(net265796), .A1(n51252), .B0(n40204), .B1(n51251),
        .C0(n40378), .C1(n51250), .Y(n13718) );
  OA22X1 U51934 ( .A0(net263368), .A1(n32572), .B0(n32580), .B1(n40075), .Y(
        n13693) );
  AOI222XL U51935 ( .A0(net265796), .A1(n51251), .B0(n40204), .B1(n51250),
        .C0(n40379), .C1(n51249), .Y(n13694) );
  OA22X1 U51936 ( .A0(net263387), .A1(n32564), .B0(n32572), .B1(n40074), .Y(
        n13669) );
  AOI222XL U51937 ( .A0(net265796), .A1(n51250), .B0(n40205), .B1(n51249),
        .C0(n40379), .C1(n51248), .Y(n13670) );
  OA22X1 U51938 ( .A0(net263387), .A1(n32556), .B0(n32564), .B1(n40074), .Y(
        n13645) );
  AOI222XL U51939 ( .A0(net265777), .A1(n51249), .B0(n40205), .B1(n51248),
        .C0(n40379), .C1(n51247), .Y(n13646) );
  OA22X1 U51940 ( .A0(net263387), .A1(n32548), .B0(n32556), .B1(n40073), .Y(
        n13621) );
  AOI222XL U51941 ( .A0(net265777), .A1(n51248), .B0(n40206), .B1(n51247),
        .C0(n40380), .C1(n51246), .Y(n13622) );
  OAI211X1 U51942 ( .A0(n32556), .A1(n42918), .B0(n13597), .C0(n13598), .Y(
        n34705) );
  OA22X1 U51943 ( .A0(net263406), .A1(n32540), .B0(n32548), .B1(n40073), .Y(
        n13597) );
  AOI222XL U51944 ( .A0(net265777), .A1(n51247), .B0(n40206), .B1(n51246),
        .C0(n40380), .C1(n51245), .Y(n13598) );
  AOI222XL U51945 ( .A0(net265758), .A1(n51246), .B0(n40206), .B1(n51245),
        .C0(n40381), .C1(n51244), .Y(n13574) );
  AOI222XL U51946 ( .A0(net265758), .A1(n51245), .B0(n40207), .B1(n51244),
        .C0(n40381), .C1(n51243), .Y(n13550) );
  OA22X1 U51947 ( .A0(net218496), .A1(n32516), .B0(n32524), .B1(n40071), .Y(
        n13525) );
  AOI222XL U51948 ( .A0(net265758), .A1(n51244), .B0(n40207), .B1(n51243),
        .C0(n40381), .C1(n51242), .Y(n13526) );
  OA22X1 U51949 ( .A0(net263444), .A1(n32508), .B0(n32516), .B1(n40071), .Y(
        n13501) );
  AOI222XL U51950 ( .A0(net265739), .A1(n51243), .B0(n40208), .B1(n51242),
        .C0(n40382), .C1(n51241), .Y(n13502) );
  OAI211X1 U51951 ( .A0(n32516), .A1(n42924), .B0(n13477), .C0(n13478), .Y(
        n34665) );
  OA22X1 U51952 ( .A0(net263444), .A1(n32500), .B0(n32508), .B1(n40070), .Y(
        n13477) );
  AOI222XL U51953 ( .A0(net265739), .A1(n51242), .B0(n40208), .B1(n51241),
        .C0(n40382), .C1(n51240), .Y(n13478) );
  OAI211X1 U51954 ( .A0(n32508), .A1(n42925), .B0(n13453), .C0(n13454), .Y(
        n34657) );
  OA22X1 U51955 ( .A0(net263463), .A1(n32492), .B0(n32500), .B1(n40070), .Y(
        n13453) );
  AOI222XL U51956 ( .A0(net265739), .A1(n51241), .B0(n40208), .B1(n51240),
        .C0(n40382), .C1(n51239), .Y(n13454) );
  OAI211X1 U51957 ( .A0(n32500), .A1(n42926), .B0(n13429), .C0(n13430), .Y(
        n34649) );
  OA22X1 U51958 ( .A0(net263463), .A1(n32484), .B0(n32492), .B1(n40069), .Y(
        n13429) );
  AOI222XL U51959 ( .A0(net265720), .A1(n51240), .B0(n40209), .B1(n51239),
        .C0(n40383), .C1(n51238), .Y(n13430) );
  OA22X1 U51960 ( .A0(net218388), .A1(n32476), .B0(n32484), .B1(n40084), .Y(
        n13405) );
  AOI222XL U51961 ( .A0(net265720), .A1(n51239), .B0(n40209), .B1(n51238),
        .C0(n40383), .C1(n51237), .Y(n13406) );
  AOI222XL U51962 ( .A0(net265701), .A1(n51238), .B0(n40210), .B1(n51237),
        .C0(n40383), .C1(n51236), .Y(n13382) );
  AOI222XL U51963 ( .A0(net265701), .A1(n51237), .B0(n40210), .B1(n51236),
        .C0(n40384), .C1(n51235), .Y(n13358) );
  OA22X1 U51964 ( .A0(net263235), .A1(n32452), .B0(n32460), .B1(n40082), .Y(
        n13333) );
  AOI222XL U51965 ( .A0(net265701), .A1(n51236), .B0(n40210), .B1(n51235),
        .C0(n40384), .C1(n51234), .Y(n13334) );
  OA22X1 U51966 ( .A0(net263235), .A1(n32444), .B0(n32452), .B1(n40082), .Y(
        n13309) );
  AOI222XL U51967 ( .A0(net265682), .A1(n51235), .B0(n40211), .B1(n51234),
        .C0(n40384), .C1(n51233), .Y(n13310) );
  OAI211X1 U51968 ( .A0(n32452), .A1(n42901), .B0(n13285), .C0(n13286), .Y(
        n34601) );
  OA22X1 U51969 ( .A0(net263235), .A1(n32436), .B0(n32444), .B1(n40081), .Y(
        n13285) );
  AOI222XL U51970 ( .A0(net265682), .A1(n51234), .B0(n40211), .B1(n51233),
        .C0(n40385), .C1(n51232), .Y(n13286) );
  OAI211X1 U51971 ( .A0(n32444), .A1(n42902), .B0(n13261), .C0(n13262), .Y(
        n34593) );
  OA22X1 U51972 ( .A0(net263254), .A1(n32428), .B0(n32436), .B1(n40081), .Y(
        n13261) );
  AOI222XL U51973 ( .A0(net265682), .A1(n51233), .B0(n40212), .B1(n51232),
        .C0(n40385), .C1(n51231), .Y(n13262) );
  OAI211X1 U51974 ( .A0(n32436), .A1(n42903), .B0(n13237), .C0(n13238), .Y(
        n34585) );
  OA22X1 U51975 ( .A0(net263254), .A1(n32420), .B0(n32428), .B1(n40080), .Y(
        n13237) );
  AOI222XL U51976 ( .A0(net221826), .A1(n51232), .B0(n40212), .B1(n51231),
        .C0(n40385), .C1(n51230), .Y(n13238) );
  OA22X1 U51977 ( .A0(net218300), .A1(n32412), .B0(n32420), .B1(n40080), .Y(
        n13213) );
  AOI222XL U51978 ( .A0(net221806), .A1(n51231), .B0(n40212), .B1(n51230),
        .C0(net217108), .C1(n51229), .Y(n13214) );
  OAI211X1 U51979 ( .A0(n32420), .A1(n42906), .B0(n13189), .C0(n13190), .Y(
        n34569) );
  AOI222XL U51980 ( .A0(net221828), .A1(n51230), .B0(n40213), .B1(n51229),
        .C0(net216982), .C1(n51228), .Y(n13190) );
  AOI222XL U51981 ( .A0(net265644), .A1(n51229), .B0(n40213), .B1(n51228),
        .C0(net216978), .C1(n51227), .Y(n13166) );
  AOI222XL U51982 ( .A0(net265644), .A1(n51228), .B0(n40214), .B1(n51227),
        .C0(net216970), .C1(n51226), .Y(n13142) );
  OAI211X1 U51983 ( .A0(n34421), .A1(n42911), .B0(n13037), .C0(n50078), .Y(
        n34521) );
  OAI222XL U51984 ( .A0(net266654), .A1(n9668), .B0(n40159), .B1(n9667), .C0(
        n40292), .C1(n34429), .Y(n13039) );
  CLKINVX1 U51985 ( .A(n19170), .Y(n49561) );
  OAI222XL U51986 ( .A0(net266381), .A1(n9667), .B0(n40174), .B1(n34429), .C0(
        n40303), .C1(n34421), .Y(n19170) );
  AOI222XL U51987 ( .A0(net265302), .A1(n49516), .B0(net218038), .B1(n51224),
        .C0(net217108), .C1(n51223), .Y(n18209) );
  AOI222XL U51988 ( .A0(net265283), .A1(n51224), .B0(n40198), .B1(n51223),
        .C0(n40318), .C1(n51222), .Y(n18185) );
  AOI222XL U51989 ( .A0(net265283), .A1(n51223), .B0(n40235), .B1(n51222),
        .C0(n40318), .C1(n51221), .Y(n18161) );
  AOI222XL U51990 ( .A0(net265283), .A1(n51222), .B0(n40236), .B1(n51221),
        .C0(n40318), .C1(n51220), .Y(n18137) );
  AOI222XL U51991 ( .A0(net265264), .A1(n51221), .B0(n40236), .B1(n51220),
        .C0(n40319), .C1(n51219), .Y(n18113) );
  AOI222XL U51992 ( .A0(net265264), .A1(n51220), .B0(n40237), .B1(n51219),
        .C0(n40319), .C1(n51218), .Y(n18089) );
  AOI222XL U51993 ( .A0(net265264), .A1(n51219), .B0(n40237), .B1(n51218),
        .C0(n40319), .C1(n51217), .Y(n18065) );
  AOI222XL U51994 ( .A0(net265245), .A1(n51218), .B0(n40237), .B1(n51217),
        .C0(n40320), .C1(n51216), .Y(n18041) );
  AOI222XL U51995 ( .A0(net265245), .A1(n51217), .B0(n40238), .B1(n51216),
        .C0(n40320), .C1(n51215), .Y(n18017) );
  AOI222XL U51996 ( .A0(net265245), .A1(n51216), .B0(n40238), .B1(n51215),
        .C0(n40321), .C1(n51214), .Y(n17993) );
  AOI222XL U51997 ( .A0(net265226), .A1(n51215), .B0(n40239), .B1(n51214),
        .C0(n40321), .C1(n51213), .Y(n17969) );
  AOI222XL U51998 ( .A0(net265226), .A1(n51214), .B0(n40239), .B1(n51213),
        .C0(n40321), .C1(n51212), .Y(n17945) );
  AOI222XL U51999 ( .A0(net265226), .A1(n51213), .B0(n40239), .B1(n51212),
        .C0(n40322), .C1(n51211), .Y(n17921) );
  AOI222XL U52000 ( .A0(net265207), .A1(n51212), .B0(n40240), .B1(n51211),
        .C0(n40322), .C1(n51210), .Y(n17897) );
  AOI222XL U52001 ( .A0(net265207), .A1(n51211), .B0(n40240), .B1(n51210),
        .C0(n40322), .C1(n51209), .Y(n17873) );
  AOI222XL U52002 ( .A0(net265207), .A1(n51210), .B0(n40241), .B1(n51209),
        .C0(n40323), .C1(n51208), .Y(n17849) );
  AOI222XL U52003 ( .A0(net265188), .A1(n51209), .B0(n40241), .B1(n51208),
        .C0(n40323), .C1(n51207), .Y(n17825) );
  AOI222XL U52004 ( .A0(net265188), .A1(n51208), .B0(n40242), .B1(n51207),
        .C0(n40323), .C1(n51206), .Y(n17801) );
  AOI222XL U52005 ( .A0(net265188), .A1(n51207), .B0(n40242), .B1(n51206),
        .C0(n40324), .C1(n51205), .Y(n17777) );
  AOI222XL U52006 ( .A0(net265169), .A1(n51206), .B0(n40242), .B1(n51205),
        .C0(n40324), .C1(n51204), .Y(n17753) );
  AOI222XL U52007 ( .A0(net265169), .A1(n51205), .B0(n40243), .B1(n51204),
        .C0(n40324), .C1(n51203), .Y(n17729) );
  AOI222XL U52008 ( .A0(net265169), .A1(n51204), .B0(n40243), .B1(n51203),
        .C0(n40325), .C1(n51202), .Y(n17705) );
  AOI222XL U52009 ( .A0(net265150), .A1(n51203), .B0(n40244), .B1(n51202),
        .C0(n40325), .C1(n51201), .Y(n17681) );
  AOI222XL U52010 ( .A0(net265150), .A1(n51202), .B0(n40244), .B1(n51201),
        .C0(n40325), .C1(n51200), .Y(n17657) );
  AOI222XL U52011 ( .A0(net265150), .A1(n51201), .B0(n40244), .B1(n51200),
        .C0(net217098), .C1(n51199), .Y(n17633) );
  AOI222XL U52012 ( .A0(net265131), .A1(n51200), .B0(n40245), .B1(n51199),
        .C0(n40349), .C1(n51198), .Y(n17609) );
  AOI222XL U52013 ( .A0(net265473), .A1(n51199), .B0(n40225), .B1(n51198),
        .C0(n40326), .C1(n51197), .Y(n17585) );
  AOI222XL U52014 ( .A0(net265454), .A1(n51198), .B0(n40225), .B1(n51197),
        .C0(n40326), .C1(n51196), .Y(n17561) );
  AOI222XL U52015 ( .A0(net265454), .A1(n51197), .B0(n40226), .B1(n51196),
        .C0(n40326), .C1(n51195), .Y(n17537) );
  AOI222XL U52016 ( .A0(net265454), .A1(n51196), .B0(n40226), .B1(n51195),
        .C0(n40327), .C1(n51194), .Y(n17513) );
  AOI222XL U52017 ( .A0(net265435), .A1(n51195), .B0(n40226), .B1(n51194),
        .C0(n40327), .C1(n51193), .Y(n17489) );
  AOI222XL U52018 ( .A0(net265435), .A1(n51194), .B0(n40227), .B1(n51193),
        .C0(n40327), .C1(n51192), .Y(n17465) );
  AOI222XL U52019 ( .A0(net265435), .A1(n51193), .B0(n40227), .B1(n51192),
        .C0(n40328), .C1(n51191), .Y(n17441) );
  AOI222XL U52020 ( .A0(net265416), .A1(n51192), .B0(n40228), .B1(n51191),
        .C0(n40328), .C1(n51190), .Y(n17417) );
  AOI222XL U52021 ( .A0(net265416), .A1(n51191), .B0(n40228), .B1(n51190),
        .C0(n40328), .C1(n51189), .Y(n17393) );
  AOI222XL U52022 ( .A0(net265416), .A1(n51190), .B0(n40228), .B1(n51189),
        .C0(n40329), .C1(n51188), .Y(n17369) );
  AOI222XL U52023 ( .A0(net265397), .A1(n51189), .B0(n40229), .B1(n51188),
        .C0(n40329), .C1(n51187), .Y(n17345) );
  AOI222XL U52024 ( .A0(net265397), .A1(n51188), .B0(n40229), .B1(n51187),
        .C0(n40329), .C1(n51186), .Y(n17321) );
  AOI222XL U52025 ( .A0(net265397), .A1(n51187), .B0(n40230), .B1(n51186),
        .C0(n40330), .C1(n51185), .Y(n17297) );
  AOI222XL U52026 ( .A0(net265378), .A1(n51186), .B0(n40230), .B1(n51185),
        .C0(n40330), .C1(n51184), .Y(n17273) );
  AOI222XL U52027 ( .A0(net265378), .A1(n51185), .B0(n40230), .B1(n51184),
        .C0(n40330), .C1(n51183), .Y(n17249) );
  AOI222XL U52028 ( .A0(net265378), .A1(n51184), .B0(n40231), .B1(n51183),
        .C0(n40331), .C1(n51182), .Y(n17225) );
  AOI222XL U52029 ( .A0(net265359), .A1(n51183), .B0(n40231), .B1(n51182),
        .C0(n40331), .C1(n51181), .Y(n17201) );
  AOI222XL U52030 ( .A0(net265359), .A1(n51182), .B0(n40232), .B1(n51181),
        .C0(n40332), .C1(n51180), .Y(n17177) );
  AOI222XL U52031 ( .A0(net265359), .A1(n51181), .B0(n40232), .B1(n51180),
        .C0(n40332), .C1(n51179), .Y(n17153) );
  AOI222XL U52032 ( .A0(net265340), .A1(n51180), .B0(n40232), .B1(n51179),
        .C0(n40332), .C1(n51178), .Y(n17129) );
  AOI222XL U52033 ( .A0(net265340), .A1(n51179), .B0(n40233), .B1(n51178),
        .C0(n40333), .C1(n51177), .Y(n17105) );
  AOI222XL U52034 ( .A0(net265340), .A1(n51178), .B0(n40233), .B1(n51177),
        .C0(n40333), .C1(n51176), .Y(n17081) );
  AOI222XL U52035 ( .A0(net265321), .A1(n51177), .B0(n40234), .B1(n51176),
        .C0(n40333), .C1(n51175), .Y(n17057) );
  AOI222XL U52036 ( .A0(net265321), .A1(n51176), .B0(n40234), .B1(n51175),
        .C0(n40334), .C1(n51174), .Y(n17033) );
  AOI222XL U52037 ( .A0(net265321), .A1(n51175), .B0(n40234), .B1(n51174),
        .C0(n40334), .C1(n51173), .Y(n17009) );
  AOI222XL U52038 ( .A0(net265302), .A1(n51174), .B0(n40235), .B1(n51173),
        .C0(n40334), .C1(n51172), .Y(n16985) );
  AOI222XL U52039 ( .A0(net265302), .A1(n51173), .B0(n40235), .B1(n51172),
        .C0(n40335), .C1(n51171), .Y(n16961) );
  AOI222XL U52040 ( .A0(net264960), .A1(n51172), .B0(n40256), .B1(n51171),
        .C0(n40335), .C1(n51170), .Y(n16937) );
  AOI222XL U52041 ( .A0(net264960), .A1(n51171), .B0(n40256), .B1(n51170),
        .C0(n40335), .C1(n51169), .Y(n16913) );
  AOI222XL U52042 ( .A0(net264941), .A1(n51170), .B0(n40257), .B1(n51169),
        .C0(n40336), .C1(n51168), .Y(n16889) );
  AOI222XL U52043 ( .A0(net264941), .A1(n51169), .B0(n40257), .B1(n51168),
        .C0(n40336), .C1(n51167), .Y(n16865) );
  AOI222XL U52044 ( .A0(net264941), .A1(n51168), .B0(n40258), .B1(n51167),
        .C0(n40336), .C1(n51166), .Y(n16841) );
  AOI222XL U52045 ( .A0(net264922), .A1(n51167), .B0(n40258), .B1(n51166),
        .C0(n40337), .C1(n51165), .Y(n16817) );
  AOI222XL U52046 ( .A0(net264922), .A1(n51166), .B0(n40258), .B1(n51165),
        .C0(n40337), .C1(n51164), .Y(n16793) );
  AOI222XL U52047 ( .A0(net264922), .A1(n51165), .B0(n40259), .B1(n51164),
        .C0(n40338), .C1(n51163), .Y(n16769) );
  AOI222XL U52048 ( .A0(net264903), .A1(n51164), .B0(n40259), .B1(n51163),
        .C0(n40338), .C1(n51162), .Y(n16745) );
  AOI222XL U52049 ( .A0(net264903), .A1(n51163), .B0(n40260), .B1(n51162),
        .C0(n40338), .C1(n51161), .Y(n16721) );
  AOI222XL U52050 ( .A0(net264903), .A1(n51162), .B0(n40260), .B1(n51161),
        .C0(n40339), .C1(n51160), .Y(n16697) );
  AOI222XL U52051 ( .A0(net264884), .A1(n51161), .B0(n40260), .B1(n51160),
        .C0(n40339), .C1(n51159), .Y(n16673) );
  AOI222XL U52052 ( .A0(net264884), .A1(n51160), .B0(n40261), .B1(n51159),
        .C0(n40339), .C1(n51158), .Y(n16649) );
  AOI222XL U52053 ( .A0(net264827), .A1(n51159), .B0(n40266), .B1(n51158),
        .C0(n40340), .C1(n51157), .Y(n16625) );
  AOI222XL U52054 ( .A0(net265036), .A1(n51158), .B0(n40264), .B1(n51157),
        .C0(n40340), .C1(n51156), .Y(n16601) );
  AOI222XL U52055 ( .A0(net264808), .A1(n51157), .B0(n40266), .B1(n51156),
        .C0(n40340), .C1(n51155), .Y(n16577) );
  AOI222XL U52056 ( .A0(net264808), .A1(n51156), .B0(n40265), .B1(n51155),
        .C0(n40341), .C1(n51154), .Y(n16553) );
  AOI222XL U52057 ( .A0(net264827), .A1(n51155), .B0(n40265), .B1(n51154),
        .C0(n40341), .C1(n51153), .Y(n16529) );
  AOI222XL U52058 ( .A0(net264827), .A1(n51154), .B0(n40264), .B1(n51153),
        .C0(n40341), .C1(n51152), .Y(n16505) );
  AOI222XL U52059 ( .A0(net264827), .A1(n51153), .B0(n40264), .B1(n51152),
        .C0(n40342), .C1(n51151), .Y(n16481) );
  AOI222XL U52060 ( .A0(net264846), .A1(n51152), .B0(n40263), .B1(n51151),
        .C0(n40342), .C1(n51150), .Y(n16457) );
  AOI222XL U52061 ( .A0(net264846), .A1(n51151), .B0(n40263), .B1(n51150),
        .C0(n40342), .C1(n51149), .Y(n16433) );
  AOI222XL U52062 ( .A0(net264846), .A1(n51150), .B0(n40263), .B1(n51149),
        .C0(n40343), .C1(n51148), .Y(n16409) );
  AOI222XL U52063 ( .A0(net264865), .A1(n51149), .B0(n40262), .B1(n51148),
        .C0(n40343), .C1(n51147), .Y(n16385) );
  AOI222XL U52064 ( .A0(net264865), .A1(n51148), .B0(n40262), .B1(n51147),
        .C0(n40344), .C1(n51146), .Y(n16361) );
  AOI222XL U52065 ( .A0(net264865), .A1(n51147), .B0(n40261), .B1(n51146),
        .C0(n40344), .C1(n51145), .Y(n16337) );
  AOI222XL U52066 ( .A0(net264884), .A1(n51146), .B0(n40261), .B1(n51145),
        .C0(n40344), .C1(n51144), .Y(n16313) );
  AOI222XL U52067 ( .A0(net265131), .A1(n51145), .B0(n40245), .B1(n51144),
        .C0(n40345), .C1(n51143), .Y(n16289) );
  AOI222XL U52068 ( .A0(net265112), .A1(n51144), .B0(n40246), .B1(n51143),
        .C0(n40345), .C1(n51142), .Y(n16265) );
  AOI222XL U52069 ( .A0(net265112), .A1(n51143), .B0(n40246), .B1(n51142),
        .C0(n40345), .C1(n51141), .Y(n16241) );
  AOI222XL U52070 ( .A0(net265112), .A1(n51142), .B0(n40247), .B1(n51141),
        .C0(n40346), .C1(n51140), .Y(n16217) );
  AOI222XL U52071 ( .A0(net221804), .A1(n51141), .B0(n40247), .B1(n51140),
        .C0(n40346), .C1(n51139), .Y(n16193) );
  AOI222XL U52072 ( .A0(net221808), .A1(n51140), .B0(n40247), .B1(n51139),
        .C0(n40346), .C1(n51138), .Y(n16169) );
  AOI222XL U52073 ( .A0(net221822), .A1(n51139), .B0(n40248), .B1(n51138),
        .C0(n40347), .C1(n51137), .Y(n16145) );
  AOI222XL U52074 ( .A0(net265074), .A1(n51138), .B0(n40248), .B1(n51137),
        .C0(n40347), .C1(n51136), .Y(n16121) );
  AOI222XL U52075 ( .A0(net265074), .A1(n51137), .B0(n40249), .B1(n51136),
        .C0(n40347), .C1(n51135), .Y(n16097) );
  AOI222XL U52076 ( .A0(net265074), .A1(n51136), .B0(n40249), .B1(n51135),
        .C0(n40348), .C1(n51134), .Y(n16073) );
  AOI222XL U52077 ( .A0(net265055), .A1(n51135), .B0(n40249), .B1(n51134),
        .C0(n40348), .C1(n51133), .Y(n16049) );
  AOI222XL U52078 ( .A0(net265055), .A1(n51134), .B0(n40250), .B1(n51133),
        .C0(n40348), .C1(n51132), .Y(n16025) );
  AOI222XL U52079 ( .A0(net265055), .A1(n51133), .B0(n40250), .B1(n51132),
        .C0(n40349), .C1(n51131), .Y(n16001) );
  AOI222XL U52080 ( .A0(net265036), .A1(n51132), .B0(n40251), .B1(n51131),
        .C0(n40349), .C1(n51130), .Y(n15977) );
  AOI222XL U52081 ( .A0(net265036), .A1(n51131), .B0(n40251), .B1(n51130),
        .C0(n40382), .C1(n51129), .Y(n15953) );
  AOI222XL U52082 ( .A0(net265036), .A1(n51130), .B0(n40252), .B1(n51129),
        .C0(n40383), .C1(n51128), .Y(n15929) );
  AOI222XL U52083 ( .A0(net265017), .A1(n51129), .B0(n40252), .B1(n51128),
        .C0(n40383), .C1(n51127), .Y(n15905) );
  AOI222XL U52084 ( .A0(net265017), .A1(n51128), .B0(n40252), .B1(n51127),
        .C0(n40350), .C1(n51126), .Y(n15881) );
  AOI222XL U52085 ( .A0(net265017), .A1(n51127), .B0(n40253), .B1(n51126),
        .C0(n40350), .C1(n51125), .Y(n15857) );
  AOI222XL U52086 ( .A0(net264998), .A1(n51126), .B0(n40253), .B1(n51125),
        .C0(n40350), .C1(n51124), .Y(n15833) );
  AOI222XL U52087 ( .A0(net264998), .A1(n51125), .B0(n40254), .B1(n51124),
        .C0(n40344), .C1(n51123), .Y(n15809) );
  AOI222XL U52088 ( .A0(net264998), .A1(n51124), .B0(n40254), .B1(n51123),
        .C0(n40344), .C1(n51122), .Y(n15785) );
  AOI222XL U52089 ( .A0(net264979), .A1(n51123), .B0(n40254), .B1(n51122),
        .C0(n40345), .C1(n51121), .Y(n15761) );
  AOI222XL U52090 ( .A0(net264979), .A1(n51122), .B0(n40255), .B1(n51121),
        .C0(n40351), .C1(n51120), .Y(n15737) );
  AOI222XL U52091 ( .A0(net264979), .A1(n51121), .B0(n40255), .B1(n51120),
        .C0(n40351), .C1(n51119), .Y(n15713) );
  AOI222XL U52092 ( .A0(net264960), .A1(n51120), .B0(n40256), .B1(n51119),
        .C0(n40351), .C1(n51118), .Y(n15689) );
  AOI222XL U52093 ( .A0(net265967), .A1(n51119), .B0(n40193), .B1(n51118),
        .C0(n40352), .C1(n51117), .Y(n15665) );
  AOI222XL U52094 ( .A0(net265967), .A1(n51118), .B0(n40193), .B1(n51117),
        .C0(n40352), .C1(n51116), .Y(n15641) );
  AOI222XL U52095 ( .A0(net265967), .A1(n51117), .B0(n40194), .B1(n51116),
        .C0(n40352), .C1(n51115), .Y(n15617) );
  AOI222XL U52096 ( .A0(net265948), .A1(n51116), .B0(n40194), .B1(n51115),
        .C0(n40353), .C1(n51114), .Y(n15593) );
  AOI222XL U52097 ( .A0(net265948), .A1(n51115), .B0(n40194), .B1(n51114),
        .C0(n40353), .C1(n51113), .Y(n15569) );
  AOI222XL U52098 ( .A0(net265948), .A1(n51114), .B0(n40195), .B1(n51113),
        .C0(n40354), .C1(n51112), .Y(n15545) );
  AOI222XL U52099 ( .A0(net265929), .A1(n51113), .B0(n40195), .B1(n51112),
        .C0(n40354), .C1(n51111), .Y(n15521) );
  AOI222XL U52100 ( .A0(net265929), .A1(n51112), .B0(n40196), .B1(n51111),
        .C0(n40354), .C1(n51110), .Y(n15497) );
  AOI222XL U52101 ( .A0(net265929), .A1(n51111), .B0(n40196), .B1(n51110),
        .C0(n40355), .C1(n51109), .Y(n15473) );
  AOI222XL U52102 ( .A0(net265910), .A1(n51110), .B0(n40196), .B1(n51109),
        .C0(n40355), .C1(n51108), .Y(n15449) );
  AOI222XL U52103 ( .A0(net265910), .A1(n51109), .B0(n40197), .B1(n51108),
        .C0(n40355), .C1(n51107), .Y(n15425) );
  AOI222XL U52104 ( .A0(net265910), .A1(n51108), .B0(n40197), .B1(n51107),
        .C0(n40356), .C1(n51106), .Y(n15401) );
  AOI222XL U52105 ( .A0(net265891), .A1(n51107), .B0(n40198), .B1(n51106),
        .C0(n40356), .C1(n51105), .Y(n15377) );
  AOI222XL U52106 ( .A0(net265891), .A1(n51106), .B0(n40198), .B1(n51105),
        .C0(n40356), .C1(n51104), .Y(n15353) );
  AOI222XL U52107 ( .A0(net265891), .A1(n51105), .B0(n40198), .B1(n51104),
        .C0(n40357), .C1(n51103), .Y(n15329) );
  AOI222XL U52108 ( .A0(net265872), .A1(n51104), .B0(n40199), .B1(n51103),
        .C0(n40357), .C1(n51102), .Y(n15305) );
  AOI222XL U52109 ( .A0(net265872), .A1(n51103), .B0(n40199), .B1(n51102),
        .C0(n40357), .C1(n51101), .Y(n15281) );
  AOI222XL U52110 ( .A0(net265872), .A1(n51102), .B0(n40200), .B1(n51101),
        .C0(n40358), .C1(n51100), .Y(n15257) );
  AOI222XL U52111 ( .A0(net265853), .A1(n51101), .B0(n40200), .B1(n51100),
        .C0(n40358), .C1(n51099), .Y(n15233) );
  AOI222XL U52112 ( .A0(net265853), .A1(n51100), .B0(n40200), .B1(n51099),
        .C0(n40358), .C1(n51098), .Y(n15209) );
  AOI222XL U52113 ( .A0(net265853), .A1(n51099), .B0(n40201), .B1(n51098),
        .C0(n40359), .C1(n51097), .Y(n15185) );
  AOI222XL U52114 ( .A0(net265834), .A1(n51098), .B0(n40201), .B1(n51097),
        .C0(n40359), .C1(n51096), .Y(n15161) );
  AOI222XL U52115 ( .A0(net265834), .A1(n51097), .B0(n40202), .B1(n51096),
        .C0(n40360), .C1(n51095), .Y(n15137) );
  AOI222XL U52116 ( .A0(net265834), .A1(n51096), .B0(n40202), .B1(n51095),
        .C0(n40360), .C1(n51094), .Y(n15113) );
  AOI222XL U52117 ( .A0(net265815), .A1(n51095), .B0(n40202), .B1(n51094),
        .C0(n40360), .C1(n51093), .Y(n15089) );
  AOI222XL U52118 ( .A0(net265815), .A1(n51094), .B0(n40203), .B1(n51093),
        .C0(n40377), .C1(n51092), .Y(n15065) );
  AOI222XL U52119 ( .A0(net265815), .A1(n51093), .B0(n40203), .B1(n51092),
        .C0(n40377), .C1(n51091), .Y(n15041) );
  AOI222XL U52120 ( .A0(net221892), .A1(n51091), .B0(n40184), .B1(n51090),
        .C0(n40361), .C1(n51089), .Y(n14993) );
  AOI222XL U52121 ( .A0(net221892), .A1(n51090), .B0(n40184), .B1(n51089),
        .C0(n40361), .C1(n51088), .Y(n14969) );
  AOI222XL U52122 ( .A0(net266119), .A1(n51089), .B0(n40184), .B1(n51088),
        .C0(n40361), .C1(n51087), .Y(n14945) );
  AOI222XL U52123 ( .A0(net266119), .A1(n51088), .B0(n40185), .B1(n51087),
        .C0(n40362), .C1(n51086), .Y(n14921) );
  OAI211X1 U52124 ( .A0(n32989), .A1(n42986), .B0(n14896), .C0(n14897), .Y(
        n35138) );
  OA22X1 U52125 ( .A0(net263748), .A1(n32973), .B0(n32981), .B1(n40053), .Y(
        n14896) );
  AOI222XL U52126 ( .A0(net266119), .A1(n51087), .B0(n40185), .B1(n51086),
        .C0(n40362), .C1(n51085), .Y(n14897) );
  OAI211X1 U52127 ( .A0(n32981), .A1(n42987), .B0(n14872), .C0(n14873), .Y(
        n35130) );
  AOI222XL U52128 ( .A0(net266100), .A1(n51086), .B0(n40194), .B1(n51085),
        .C0(n40362), .C1(n51084), .Y(n14873) );
  OAI211X1 U52129 ( .A0(n32973), .A1(n42988), .B0(n14848), .C0(n14849), .Y(
        n35122) );
  OA22X1 U52130 ( .A0(net263767), .A1(n32957), .B0(n32965), .B1(n40052), .Y(
        n14848) );
  AOI222XL U52131 ( .A0(net266100), .A1(n51085), .B0(n40195), .B1(n51084),
        .C0(n40363), .C1(n51083), .Y(n14849) );
  OAI211X1 U52132 ( .A0(n32965), .A1(n42989), .B0(n14824), .C0(n14825), .Y(
        n35114) );
  OA22X1 U52133 ( .A0(net262665), .A1(n32949), .B0(n32957), .B1(n40052), .Y(
        n14824) );
  AOI222XL U52134 ( .A0(net266100), .A1(n51084), .B0(n40195), .B1(n51083),
        .C0(n40363), .C1(n51082), .Y(n14825) );
  OAI211X1 U52135 ( .A0(n32957), .A1(n42990), .B0(n14800), .C0(n14801), .Y(
        n35106) );
  OA22X1 U52136 ( .A0(net263064), .A1(n32941), .B0(n32949), .B1(n40051), .Y(
        n14800) );
  AOI222XL U52137 ( .A0(net266081), .A1(n51083), .B0(n40186), .B1(n51082),
        .C0(n40363), .C1(n51081), .Y(n14801) );
  OAI211X1 U52138 ( .A0(n32949), .A1(n42963), .B0(n14776), .C0(n14777), .Y(
        n35098) );
  OA22X1 U52139 ( .A0(net263805), .A1(n32933), .B0(n32941), .B1(n40051), .Y(
        n14776) );
  AOI222XL U52140 ( .A0(net266081), .A1(n51082), .B0(n40186), .B1(n51081),
        .C0(n40364), .C1(n51080), .Y(n14777) );
  OAI211X1 U52141 ( .A0(n32941), .A1(n42960), .B0(n14752), .C0(n14753), .Y(
        n35090) );
  OA22X1 U52142 ( .A0(net263805), .A1(n32925), .B0(n32933), .B1(n40050), .Y(
        n14752) );
  AOI222XL U52143 ( .A0(net266081), .A1(n51081), .B0(n40187), .B1(n51080),
        .C0(n40367), .C1(n51079), .Y(n14753) );
  OAI211X1 U52144 ( .A0(n32933), .A1(n42961), .B0(n14728), .C0(n14729), .Y(
        n35082) );
  OA22X1 U52145 ( .A0(net263824), .A1(n32917), .B0(n32925), .B1(n40049), .Y(
        n14728) );
  AOI222XL U52146 ( .A0(net266062), .A1(n51080), .B0(n40187), .B1(n51079),
        .C0(n40364), .C1(n51078), .Y(n14729) );
  OAI211X1 U52147 ( .A0(n32925), .A1(n42962), .B0(n14704), .C0(n14705), .Y(
        n35074) );
  OA22X1 U52148 ( .A0(net263824), .A1(n32909), .B0(n32917), .B1(n40049), .Y(
        n14704) );
  AOI222XL U52149 ( .A0(net266062), .A1(n51079), .B0(n40188), .B1(n51078),
        .C0(n40364), .C1(n51077), .Y(n14705) );
  OAI211X1 U52150 ( .A0(n32917), .A1(n42964), .B0(n14680), .C0(n14681), .Y(
        n35066) );
  OA22X1 U52151 ( .A0(net263843), .A1(n32901), .B0(n32909), .B1(n40048), .Y(
        n14680) );
  AOI222XL U52152 ( .A0(net266062), .A1(n51078), .B0(n40188), .B1(n51077),
        .C0(n40364), .C1(n51076), .Y(n14681) );
  OAI211X1 U52153 ( .A0(n32909), .A1(n42965), .B0(n14656), .C0(n14657), .Y(
        n35058) );
  OA22X1 U52154 ( .A0(net263843), .A1(n32893), .B0(n32901), .B1(n40048), .Y(
        n14656) );
  AOI222XL U52155 ( .A0(net266043), .A1(n51077), .B0(n40188), .B1(n51076),
        .C0(n40365), .C1(n51075), .Y(n14657) );
  OAI211X1 U52156 ( .A0(n32901), .A1(n42966), .B0(n14632), .C0(n14633), .Y(
        n35050) );
  OA22X1 U52157 ( .A0(net263843), .A1(n32885), .B0(n32893), .B1(n40047), .Y(
        n14632) );
  AOI222XL U52158 ( .A0(net266043), .A1(n51076), .B0(n40189), .B1(n51075),
        .C0(n40365), .C1(n51074), .Y(n14633) );
  OAI211X1 U52159 ( .A0(n32893), .A1(n42967), .B0(n14608), .C0(n14609), .Y(
        n35042) );
  OA22X1 U52160 ( .A0(net263862), .A1(n32877), .B0(n32885), .B1(n40047), .Y(
        n14608) );
  AOI222XL U52161 ( .A0(net266043), .A1(n51075), .B0(n40189), .B1(n51074),
        .C0(n40365), .C1(n51073), .Y(n14609) );
  OAI211X1 U52162 ( .A0(n32885), .A1(n42968), .B0(n14584), .C0(n14585), .Y(
        n35034) );
  OA22X1 U52163 ( .A0(net263862), .A1(n32869), .B0(n32877), .B1(n40046), .Y(
        n14584) );
  AOI222XL U52164 ( .A0(net266024), .A1(n51074), .B0(n40190), .B1(n51073),
        .C0(n40366), .C1(n51072), .Y(n14585) );
  OAI211X1 U52165 ( .A0(n32877), .A1(n42969), .B0(n14560), .C0(n14561), .Y(
        n35026) );
  OA22X1 U52166 ( .A0(net263064), .A1(n32861), .B0(n32869), .B1(n40092), .Y(
        n14560) );
  AOI222XL U52167 ( .A0(net266024), .A1(n51073), .B0(n40190), .B1(n51072),
        .C0(n40366), .C1(n51071), .Y(n14561) );
  OAI211X1 U52168 ( .A0(n32869), .A1(n42971), .B0(n14536), .C0(n14537), .Y(
        n35018) );
  OA22X1 U52169 ( .A0(net263064), .A1(n32853), .B0(n32861), .B1(n40092), .Y(
        n14536) );
  AOI222XL U52170 ( .A0(net266024), .A1(n51072), .B0(n40190), .B1(n51071),
        .C0(n40366), .C1(n51070), .Y(n14537) );
  OAI211X1 U52171 ( .A0(n32861), .A1(n42972), .B0(n14512), .C0(n14513), .Y(
        n35010) );
  OA22X1 U52172 ( .A0(net263083), .A1(n32845), .B0(n32853), .B1(n40091), .Y(
        n14512) );
  AOI222XL U52173 ( .A0(net266005), .A1(n51071), .B0(n40191), .B1(n51070),
        .C0(n40367), .C1(n51069), .Y(n14513) );
  OAI211X1 U52174 ( .A0(n32853), .A1(n42973), .B0(n14488), .C0(n14489), .Y(
        n35002) );
  OA22X1 U52175 ( .A0(net263083), .A1(n32837), .B0(n32845), .B1(n40091), .Y(
        n14488) );
  AOI222XL U52176 ( .A0(net266005), .A1(n51070), .B0(n40191), .B1(n51069),
        .C0(n40367), .C1(n51068), .Y(n14489) );
  OAI211X1 U52177 ( .A0(n32845), .A1(n42974), .B0(n14464), .C0(n14465), .Y(
        n34994) );
  OA22X1 U52178 ( .A0(net263102), .A1(n32829), .B0(n32837), .B1(n40090), .Y(
        n14464) );
  AOI222XL U52179 ( .A0(net266005), .A1(n51069), .B0(n40192), .B1(n51068),
        .C0(n40367), .C1(n51067), .Y(n14465) );
  OAI211X1 U52180 ( .A0(n32837), .A1(n42975), .B0(n14440), .C0(n14441), .Y(
        n34986) );
  OA22X1 U52181 ( .A0(net263102), .A1(n32821), .B0(n32829), .B1(n40090), .Y(
        n14440) );
  AOI222XL U52182 ( .A0(net265416), .A1(n51068), .B0(n40192), .B1(n51067),
        .C0(n40368), .C1(n51066), .Y(n14441) );
  OAI211X1 U52183 ( .A0(n32829), .A1(n42879), .B0(n14416), .C0(n14417), .Y(
        n34978) );
  OA22X1 U52184 ( .A0(net263121), .A1(n32813), .B0(n32821), .B1(n40089), .Y(
        n14416) );
  AOI222XL U52185 ( .A0(net265264), .A1(n51067), .B0(n40192), .B1(n51066),
        .C0(n40368), .C1(n51065), .Y(n14417) );
  OAI211X1 U52186 ( .A0(n32821), .A1(n42880), .B0(n14392), .C0(n14393), .Y(
        n34970) );
  OA22X1 U52187 ( .A0(net263121), .A1(n32805), .B0(n32813), .B1(n40089), .Y(
        n14392) );
  AOI222XL U52188 ( .A0(net265530), .A1(n51066), .B0(n40187), .B1(n51065),
        .C0(n40368), .C1(n51064), .Y(n14393) );
  OAI211X1 U52189 ( .A0(n32813), .A1(n42881), .B0(n14368), .C0(n14369), .Y(
        n34962) );
  OA22X1 U52190 ( .A0(net263140), .A1(n32797), .B0(n32805), .B1(n40088), .Y(
        n14368) );
  AOI222XL U52191 ( .A0(net265625), .A1(n51065), .B0(n40214), .B1(n51064),
        .C0(n40369), .C1(n51063), .Y(n14369) );
  OAI211X1 U52192 ( .A0(n32805), .A1(n42883), .B0(n14344), .C0(n14345), .Y(
        n34954) );
  OA22X1 U52193 ( .A0(net263140), .A1(n32789), .B0(n32797), .B1(n40088), .Y(
        n14344) );
  AOI222XL U52194 ( .A0(net265625), .A1(n51064), .B0(n40215), .B1(n51063),
        .C0(n40369), .C1(n51062), .Y(n14345) );
  OAI211X1 U52195 ( .A0(n32797), .A1(n42884), .B0(n14320), .C0(n14321), .Y(
        n34946) );
  OA22X1 U52196 ( .A0(net263140), .A1(n32781), .B0(n32789), .B1(n40087), .Y(
        n14320) );
  AOI222XL U52197 ( .A0(net265625), .A1(n51063), .B0(n40215), .B1(n51062),
        .C0(n40370), .C1(n51061), .Y(n14321) );
  OAI211X1 U52198 ( .A0(n32789), .A1(n42885), .B0(n14296), .C0(n14297), .Y(
        n34938) );
  OA22X1 U52199 ( .A0(net263159), .A1(n32773), .B0(n32781), .B1(n40087), .Y(
        n14296) );
  AOI222XL U52200 ( .A0(net265606), .A1(n51062), .B0(n40216), .B1(n51061),
        .C0(n40370), .C1(n51060), .Y(n14297) );
  OAI211X1 U52201 ( .A0(n32781), .A1(n42886), .B0(n14272), .C0(n14273), .Y(
        n34930) );
  OA22X1 U52202 ( .A0(net263159), .A1(n32765), .B0(n32773), .B1(n40086), .Y(
        n14272) );
  AOI222XL U52203 ( .A0(net265606), .A1(n51061), .B0(n40216), .B1(n51060),
        .C0(n40370), .C1(n51059), .Y(n14273) );
  OAI211X1 U52204 ( .A0(n32773), .A1(n42887), .B0(n14248), .C0(n14249), .Y(
        n34922) );
  OA22X1 U52205 ( .A0(net263178), .A1(n32757), .B0(n32765), .B1(n40086), .Y(
        n14248) );
  AOI222XL U52206 ( .A0(net265606), .A1(n51060), .B0(n40216), .B1(n51059),
        .C0(n40371), .C1(n51058), .Y(n14249) );
  OAI211X1 U52207 ( .A0(n32765), .A1(n42888), .B0(n14224), .C0(n14225), .Y(
        n34914) );
  OA22X1 U52208 ( .A0(net263178), .A1(n32749), .B0(n32757), .B1(n40085), .Y(
        n14224) );
  AOI222XL U52209 ( .A0(net265587), .A1(n51059), .B0(n40217), .B1(n51058),
        .C0(n40371), .C1(n51057), .Y(n14225) );
  OAI211X1 U52210 ( .A0(n32757), .A1(n42890), .B0(n14200), .C0(n14201), .Y(
        n34906) );
  OA22X1 U52211 ( .A0(net218434), .A1(n32741), .B0(n32749), .B1(n40085), .Y(
        n14200) );
  AOI222XL U52212 ( .A0(net265587), .A1(n51058), .B0(n40217), .B1(n51057),
        .C0(n40371), .C1(n51056), .Y(n14201) );
  OAI211X1 U52213 ( .A0(n32749), .A1(n42891), .B0(n14176), .C0(n14177), .Y(
        n34898) );
  OA22X1 U52214 ( .A0(net262931), .A1(n32733), .B0(n32741), .B1(n40100), .Y(
        n14176) );
  AOI222XL U52215 ( .A0(net265587), .A1(n51057), .B0(n40218), .B1(n51056),
        .C0(n40372), .C1(n51055), .Y(n14177) );
  OAI211X1 U52216 ( .A0(n32741), .A1(n42892), .B0(n14152), .C0(n14153), .Y(
        n34890) );
  OA22X1 U52217 ( .A0(net262931), .A1(n32725), .B0(n32733), .B1(n40100), .Y(
        n14152) );
  AOI222XL U52218 ( .A0(net265568), .A1(n51056), .B0(n40218), .B1(n51055),
        .C0(n40372), .C1(n51054), .Y(n14153) );
  OAI211X1 U52219 ( .A0(n32733), .A1(n42893), .B0(n14128), .C0(n14129), .Y(
        n34882) );
  OA22X1 U52220 ( .A0(net262950), .A1(n32717), .B0(n32725), .B1(n40099), .Y(
        n14128) );
  AOI222XL U52221 ( .A0(net265568), .A1(n51055), .B0(n40218), .B1(n51054),
        .C0(n40372), .C1(n51053), .Y(n14129) );
  OAI211X1 U52222 ( .A0(n32725), .A1(n42894), .B0(n14104), .C0(n14105), .Y(
        n34874) );
  OA22X1 U52223 ( .A0(net262950), .A1(n32709), .B0(n32717), .B1(n40099), .Y(
        n14104) );
  AOI222XL U52224 ( .A0(net265568), .A1(n51054), .B0(n40219), .B1(n51053),
        .C0(n40373), .C1(n51052), .Y(n14105) );
  OAI211X1 U52225 ( .A0(n32717), .A1(n42863), .B0(n14080), .C0(n14081), .Y(
        n34866) );
  OA22X1 U52226 ( .A0(net262969), .A1(n32701), .B0(n32709), .B1(n40098), .Y(
        n14080) );
  AOI222XL U52227 ( .A0(net265549), .A1(n51053), .B0(n40219), .B1(n51052),
        .C0(n40373), .C1(n51051), .Y(n14081) );
  OAI211X1 U52228 ( .A0(n32709), .A1(n42864), .B0(n14056), .C0(n14057), .Y(
        n34858) );
  OA22X1 U52229 ( .A0(net262969), .A1(n32693), .B0(n32701), .B1(n40098), .Y(
        n14056) );
  AOI222XL U52230 ( .A0(net265549), .A1(n51052), .B0(n40220), .B1(n51051),
        .C0(n40373), .C1(n51050), .Y(n14057) );
  OAI211X1 U52231 ( .A0(n32701), .A1(n42865), .B0(n14032), .C0(n14033), .Y(
        n34850) );
  OA22X1 U52232 ( .A0(net262988), .A1(n32685), .B0(n32693), .B1(n40097), .Y(
        n14032) );
  AOI222XL U52233 ( .A0(net265549), .A1(n51051), .B0(n40220), .B1(n51050),
        .C0(n40374), .C1(n51049), .Y(n14033) );
  OAI211X1 U52234 ( .A0(n32693), .A1(n42867), .B0(n14008), .C0(n14009), .Y(
        n34842) );
  OA22X1 U52235 ( .A0(net262988), .A1(n32677), .B0(n32685), .B1(n40097), .Y(
        n14008) );
  AOI222XL U52236 ( .A0(net265530), .A1(n51050), .B0(n40220), .B1(n51049),
        .C0(n40374), .C1(n51048), .Y(n14009) );
  OAI211X1 U52237 ( .A0(n32685), .A1(n42868), .B0(n13984), .C0(n13985), .Y(
        n34834) );
  OA22X1 U52238 ( .A0(net263007), .A1(n32669), .B0(n32677), .B1(n40096), .Y(
        n13984) );
  AOI222XL U52239 ( .A0(net265530), .A1(n51049), .B0(n40221), .B1(n51048),
        .C0(n40374), .C1(n51047), .Y(n13985) );
  OAI211X1 U52240 ( .A0(n32677), .A1(n42869), .B0(n13960), .C0(n13961), .Y(
        n34826) );
  OA22X1 U52241 ( .A0(net263007), .A1(n32661), .B0(n32669), .B1(n40095), .Y(
        n13960) );
  AOI222XL U52242 ( .A0(net265530), .A1(n51048), .B0(n40221), .B1(n51047),
        .C0(n40375), .C1(n51046), .Y(n13961) );
  OAI211X1 U52243 ( .A0(n32669), .A1(n42870), .B0(n13936), .C0(n13937), .Y(
        n34818) );
  OA22X1 U52244 ( .A0(net263007), .A1(n32653), .B0(n32661), .B1(n40095), .Y(
        n13936) );
  AOI222XL U52245 ( .A0(net265511), .A1(n51047), .B0(n40222), .B1(n51046),
        .C0(n40375), .C1(n51045), .Y(n13937) );
  OAI211X1 U52246 ( .A0(n32661), .A1(n42871), .B0(n13912), .C0(n13913), .Y(
        n34810) );
  OA22X1 U52247 ( .A0(net263026), .A1(n32645), .B0(n32653), .B1(n40094), .Y(
        n13912) );
  AOI222XL U52248 ( .A0(net265511), .A1(n51046), .B0(n40222), .B1(n51045),
        .C0(n40376), .C1(n51044), .Y(n13913) );
  OAI211X1 U52249 ( .A0(n32653), .A1(n42872), .B0(n13888), .C0(n13889), .Y(
        n34802) );
  OA22X1 U52250 ( .A0(net263026), .A1(n32637), .B0(n32645), .B1(n40094), .Y(
        n13888) );
  AOI222XL U52251 ( .A0(net265511), .A1(n51045), .B0(n40222), .B1(n51044),
        .C0(n40376), .C1(n51043), .Y(n13889) );
  OAI211X1 U52252 ( .A0(n32645), .A1(n42874), .B0(n13864), .C0(n13865), .Y(
        n34794) );
  OA22X1 U52253 ( .A0(net263045), .A1(n32629), .B0(n32637), .B1(n40093), .Y(
        n13864) );
  AOI222XL U52254 ( .A0(net265492), .A1(n51044), .B0(n40223), .B1(n51043),
        .C0(n40376), .C1(n51042), .Y(n13865) );
  OAI211X1 U52255 ( .A0(n32637), .A1(n42875), .B0(n13840), .C0(n13841), .Y(
        n34786) );
  OA22X1 U52256 ( .A0(net263045), .A1(n32621), .B0(n32629), .B1(n40093), .Y(
        n13840) );
  AOI222XL U52257 ( .A0(net265492), .A1(n51043), .B0(n40223), .B1(n51042),
        .C0(n40377), .C1(n51041), .Y(n13841) );
  OAI211X1 U52258 ( .A0(n32629), .A1(n42876), .B0(n13816), .C0(n13817), .Y(
        n34778) );
  OA22X1 U52259 ( .A0(net263064), .A1(n32613), .B0(n32621), .B1(n40092), .Y(
        n13816) );
  AOI222XL U52260 ( .A0(net265492), .A1(n51042), .B0(n40224), .B1(n51041),
        .C0(n40377), .C1(n51040), .Y(n13817) );
  OAI211X1 U52261 ( .A0(n32621), .A1(n42877), .B0(n13792), .C0(n13793), .Y(
        n34770) );
  OA22X1 U52262 ( .A0(net263330), .A1(n32605), .B0(n32613), .B1(n40077), .Y(
        n13792) );
  AOI222XL U52263 ( .A0(net265473), .A1(n51041), .B0(n40224), .B1(n51040),
        .C0(n40377), .C1(n51039), .Y(n13793) );
  OAI211X1 U52264 ( .A0(n32613), .A1(n42878), .B0(n13768), .C0(n13769), .Y(
        n34762) );
  OA22X1 U52265 ( .A0(net263349), .A1(n32597), .B0(n32605), .B1(n40077), .Y(
        n13768) );
  AOI222XL U52266 ( .A0(net265473), .A1(n51040), .B0(n40224), .B1(n51039),
        .C0(n40378), .C1(n51038), .Y(n13769) );
  OAI211X1 U52267 ( .A0(n32605), .A1(n42919), .B0(n13744), .C0(n13745), .Y(
        n34754) );
  OA22X1 U52268 ( .A0(net263349), .A1(n32589), .B0(n32597), .B1(n40076), .Y(
        n13744) );
  AOI222XL U52269 ( .A0(net265815), .A1(n51039), .B0(n40204), .B1(n51038),
        .C0(n40378), .C1(n51037), .Y(n13745) );
  OAI211X1 U52270 ( .A0(n32597), .A1(n42912), .B0(n13720), .C0(n13721), .Y(
        n34746) );
  OA22X1 U52271 ( .A0(net263368), .A1(n32581), .B0(n32589), .B1(n40076), .Y(
        n13720) );
  AOI222XL U52272 ( .A0(net265796), .A1(n51038), .B0(n40204), .B1(n51037),
        .C0(n40378), .C1(n51036), .Y(n13721) );
  OAI211X1 U52273 ( .A0(n32589), .A1(n42914), .B0(n13696), .C0(n13697), .Y(
        n34738) );
  OA22X1 U52274 ( .A0(net263368), .A1(n32573), .B0(n32581), .B1(n40075), .Y(
        n13696) );
  AOI222XL U52275 ( .A0(net265796), .A1(n51037), .B0(n40204), .B1(n51036),
        .C0(n40379), .C1(n51035), .Y(n13697) );
  OAI211X1 U52276 ( .A0(n32581), .A1(n42915), .B0(n13672), .C0(n13673), .Y(
        n34730) );
  OA22X1 U52277 ( .A0(net263368), .A1(n32565), .B0(n32573), .B1(n40075), .Y(
        n13672) );
  AOI222XL U52278 ( .A0(net265796), .A1(n51036), .B0(n40205), .B1(n51035),
        .C0(n40379), .C1(n51034), .Y(n13673) );
  OAI211X1 U52279 ( .A0(n32573), .A1(n42916), .B0(n13648), .C0(n13649), .Y(
        n34722) );
  OA22X1 U52280 ( .A0(net263387), .A1(n32557), .B0(n32565), .B1(n40074), .Y(
        n13648) );
  AOI222XL U52281 ( .A0(net265777), .A1(n51035), .B0(n40205), .B1(n51034),
        .C0(n40379), .C1(n51033), .Y(n13649) );
  OAI211X1 U52282 ( .A0(n32565), .A1(n42917), .B0(n13624), .C0(n13625), .Y(
        n34714) );
  OA22X1 U52283 ( .A0(net263387), .A1(n32549), .B0(n32557), .B1(n40074), .Y(
        n13624) );
  AOI222XL U52284 ( .A0(net265777), .A1(n51034), .B0(n40206), .B1(n51033),
        .C0(n40380), .C1(n51032), .Y(n13625) );
  OAI211X1 U52285 ( .A0(n32557), .A1(n42918), .B0(n13600), .C0(n13601), .Y(
        n34706) );
  OA22X1 U52286 ( .A0(net263406), .A1(n32541), .B0(n32549), .B1(n40073), .Y(
        n13600) );
  AOI222XL U52287 ( .A0(net265777), .A1(n51033), .B0(n40206), .B1(n51032),
        .C0(n40380), .C1(n51031), .Y(n13601) );
  OAI211X1 U52288 ( .A0(n32549), .A1(n42919), .B0(n13576), .C0(n13577), .Y(
        n34698) );
  OA22X1 U52289 ( .A0(net263406), .A1(n32533), .B0(n32541), .B1(n40072), .Y(
        n13576) );
  AOI222XL U52290 ( .A0(net265758), .A1(n51032), .B0(n40206), .B1(n51031),
        .C0(n40380), .C1(n51030), .Y(n13577) );
  OAI211X1 U52291 ( .A0(n32541), .A1(n42921), .B0(n13552), .C0(n13553), .Y(
        n34690) );
  OA22X1 U52292 ( .A0(net218378), .A1(n32525), .B0(n32533), .B1(n40072), .Y(
        n13552) );
  AOI222XL U52293 ( .A0(net265758), .A1(n51031), .B0(n40207), .B1(n51030),
        .C0(n40381), .C1(n51029), .Y(n13553) );
  OAI211X1 U52294 ( .A0(n32533), .A1(n42922), .B0(n13528), .C0(n13529), .Y(
        n34682) );
  OA22X1 U52295 ( .A0(net218380), .A1(n32517), .B0(n32525), .B1(n40071), .Y(
        n13528) );
  AOI222XL U52296 ( .A0(net265758), .A1(n51030), .B0(n40207), .B1(n51029),
        .C0(n40381), .C1(n51028), .Y(n13529) );
  OAI211X1 U52297 ( .A0(n32525), .A1(n42923), .B0(n13504), .C0(n13505), .Y(
        n34674) );
  OA22X1 U52298 ( .A0(net263444), .A1(n32509), .B0(n32517), .B1(n40071), .Y(
        n13504) );
  AOI222XL U52299 ( .A0(net265739), .A1(n51029), .B0(n40208), .B1(n51028),
        .C0(n40382), .C1(n51027), .Y(n13505) );
  OAI211X1 U52300 ( .A0(n32517), .A1(n42924), .B0(n13480), .C0(n13481), .Y(
        n34666) );
  OA22X1 U52301 ( .A0(net263444), .A1(n32501), .B0(n32509), .B1(n40070), .Y(
        n13480) );
  AOI222XL U52302 ( .A0(net265739), .A1(n51028), .B0(n40208), .B1(n51027),
        .C0(n40382), .C1(n51026), .Y(n13481) );
  OAI211X1 U52303 ( .A0(n32509), .A1(n42925), .B0(n13456), .C0(n13457), .Y(
        n34658) );
  OA22X1 U52304 ( .A0(net263463), .A1(n32493), .B0(n32501), .B1(n40070), .Y(
        n13456) );
  AOI222XL U52305 ( .A0(net265739), .A1(n51027), .B0(n40208), .B1(n51026),
        .C0(n40382), .C1(n51025), .Y(n13457) );
  OAI211X1 U52306 ( .A0(n32501), .A1(n42926), .B0(n13432), .C0(n13433), .Y(
        n34650) );
  OA22X1 U52307 ( .A0(net263463), .A1(n32485), .B0(n32493), .B1(n40069), .Y(
        n13432) );
  AOI222XL U52308 ( .A0(net265720), .A1(n51026), .B0(n40209), .B1(n51025),
        .C0(n40383), .C1(n51024), .Y(n13433) );
  OAI211X1 U52309 ( .A0(n32493), .A1(n42903), .B0(n13408), .C0(n13409), .Y(
        n34642) );
  OA22X1 U52310 ( .A0(net261943), .A1(n32477), .B0(n32485), .B1(n40084), .Y(
        n13408) );
  AOI222XL U52311 ( .A0(net265720), .A1(n51025), .B0(n40209), .B1(n51024),
        .C0(n40383), .C1(n51023), .Y(n13409) );
  OAI211X1 U52312 ( .A0(n32485), .A1(n42896), .B0(n13384), .C0(n13385), .Y(
        n34634) );
  OA22X1 U52313 ( .A0(net263216), .A1(n32469), .B0(n32477), .B1(n40083), .Y(
        n13384) );
  AOI222XL U52314 ( .A0(net265720), .A1(n51024), .B0(n40210), .B1(n51023),
        .C0(n40383), .C1(n51022), .Y(n13385) );
  OAI211X1 U52315 ( .A0(n32477), .A1(n42897), .B0(n13360), .C0(n13361), .Y(
        n34626) );
  OA22X1 U52316 ( .A0(net263216), .A1(n32461), .B0(n32469), .B1(n40083), .Y(
        n13360) );
  AOI222XL U52317 ( .A0(net265701), .A1(n51023), .B0(n40210), .B1(n51022),
        .C0(n40384), .C1(n51021), .Y(n13361) );
  OAI211X1 U52318 ( .A0(n32469), .A1(n42899), .B0(n13336), .C0(n13337), .Y(
        n34618) );
  OA22X1 U52319 ( .A0(net263235), .A1(n32453), .B0(n32461), .B1(n40082), .Y(
        n13336) );
  AOI222XL U52320 ( .A0(net265701), .A1(n51022), .B0(n40210), .B1(n51021),
        .C0(n40384), .C1(n51020), .Y(n13337) );
  OAI211X1 U52321 ( .A0(n32461), .A1(n42900), .B0(n13312), .C0(n13313), .Y(
        n34610) );
  OA22X1 U52322 ( .A0(net263235), .A1(n32445), .B0(n32453), .B1(n40082), .Y(
        n13312) );
  AOI222XL U52323 ( .A0(net265701), .A1(n51021), .B0(n40211), .B1(n51020),
        .C0(n40384), .C1(n51019), .Y(n13313) );
  OAI211X1 U52324 ( .A0(n32453), .A1(n42901), .B0(n13288), .C0(n13289), .Y(
        n34602) );
  OA22X1 U52325 ( .A0(net263235), .A1(n32437), .B0(n32445), .B1(n40081), .Y(
        n13288) );
  AOI222XL U52326 ( .A0(net265682), .A1(n51020), .B0(n40211), .B1(n51019),
        .C0(n40385), .C1(n51018), .Y(n13289) );
  OAI211X1 U52327 ( .A0(n32445), .A1(n42902), .B0(n13264), .C0(n13265), .Y(
        n34594) );
  OA22X1 U52328 ( .A0(net263254), .A1(n32429), .B0(n32437), .B1(n40081), .Y(
        n13264) );
  AOI222XL U52329 ( .A0(net265682), .A1(n51019), .B0(n40212), .B1(n51018),
        .C0(n40385), .C1(n51017), .Y(n13265) );
  OAI211X1 U52330 ( .A0(n32437), .A1(n42903), .B0(n13240), .C0(n13241), .Y(
        n34586) );
  OA22X1 U52331 ( .A0(net263254), .A1(n32421), .B0(n32429), .B1(n40080), .Y(
        n13240) );
  AOI222XL U52332 ( .A0(net265682), .A1(n51018), .B0(n40212), .B1(n51017),
        .C0(n40385), .C1(n51016), .Y(n13241) );
  OAI211X1 U52333 ( .A0(n32429), .A1(n42904), .B0(n13216), .C0(n13217), .Y(
        n34578) );
  OA22X1 U52334 ( .A0(net218426), .A1(n32413), .B0(n32421), .B1(n40080), .Y(
        n13216) );
  AOI222XL U52335 ( .A0(net265112), .A1(n51017), .B0(n40212), .B1(n51016),
        .C0(net217030), .C1(n51015), .Y(n13217) );
  OAI211X1 U52336 ( .A0(n32421), .A1(n42906), .B0(n13192), .C0(n13193), .Y(
        n34570) );
  OA22X1 U52337 ( .A0(net218332), .A1(n32405), .B0(n32413), .B1(n40079), .Y(
        n13192) );
  AOI222XL U52338 ( .A0(net221812), .A1(n51016), .B0(n40213), .B1(n51015),
        .C0(net217048), .C1(n51014), .Y(n13193) );
  OAI211X1 U52339 ( .A0(n32413), .A1(n42907), .B0(n13168), .C0(n13169), .Y(
        n34562) );
  AOI222XL U52340 ( .A0(net265492), .A1(n51015), .B0(n40213), .B1(n51014),
        .C0(net217028), .C1(n51013), .Y(n13169) );
  OAI211X1 U52341 ( .A0(n32405), .A1(n42908), .B0(n13144), .C0(n13145), .Y(
        n34554) );
  AOI222XL U52342 ( .A0(net265644), .A1(n51014), .B0(n40214), .B1(n51013),
        .C0(n40381), .C1(n51012), .Y(n13145) );
  OAI211X1 U52343 ( .A0(n34422), .A1(n42911), .B0(n13034), .C0(n50079), .Y(
        n34520) );
  OAI222XL U52344 ( .A0(net266654), .A1(n9666), .B0(n40159), .B1(n9665), .C0(
        n40292), .C1(n34430), .Y(n13036) );
  CLKINVX1 U52345 ( .A(n19173), .Y(n49560) );
  OAI222XL U52346 ( .A0(net266381), .A1(n9665), .B0(n40171), .B1(n34430), .C0(
        n40298), .C1(n34422), .Y(n19173) );
  OAI211X1 U52347 ( .A0(n34102), .A1(n42826), .B0(n18235), .C0(n18236), .Y(
        n36251) );
  OA22X1 U52348 ( .A0(net262855), .A1(n34086), .B0(n34094), .B1(n40104), .Y(
        n18235) );
  AOI222XL U52349 ( .A0(net264960), .A1(n49515), .B0(n40225), .B1(n49514),
        .C0(n40368), .C1(n51010), .Y(n18236) );
  AOI222XL U52350 ( .A0(net265302), .A1(n49514), .B0(n40189), .B1(n51010),
        .C0(net217108), .C1(n51009), .Y(n18212) );
  AOI222XL U52351 ( .A0(net265283), .A1(n51010), .B0(n40190), .B1(n51009),
        .C0(n40318), .C1(n51008), .Y(n18188) );
  AOI222XL U52352 ( .A0(net265283), .A1(n51009), .B0(n40198), .B1(n51008),
        .C0(n40318), .C1(n51007), .Y(n18164) );
  AOI222XL U52353 ( .A0(net265283), .A1(n51008), .B0(n40236), .B1(n51007),
        .C0(n40318), .C1(n51006), .Y(n18140) );
  AOI222XL U52354 ( .A0(net265264), .A1(n51007), .B0(n40236), .B1(n51006),
        .C0(n40319), .C1(n51005), .Y(n18116) );
  AOI222XL U52355 ( .A0(net265264), .A1(n51006), .B0(n40237), .B1(n51005),
        .C0(n40319), .C1(n51004), .Y(n18092) );
  AOI222XL U52356 ( .A0(net265264), .A1(n51005), .B0(n40237), .B1(n51004),
        .C0(n40319), .C1(n51003), .Y(n18068) );
  AOI222XL U52357 ( .A0(net265245), .A1(n51004), .B0(n40237), .B1(n51003),
        .C0(n40320), .C1(n51002), .Y(n18044) );
  AOI222XL U52358 ( .A0(net265245), .A1(n51003), .B0(n40238), .B1(n51002),
        .C0(n40320), .C1(n51001), .Y(n18020) );
  AOI222XL U52359 ( .A0(net265245), .A1(n51002), .B0(n40238), .B1(n51001),
        .C0(n40320), .C1(n51000), .Y(n17996) );
  AOI222XL U52360 ( .A0(net265226), .A1(n51001), .B0(n40239), .B1(n51000),
        .C0(n40321), .C1(n50999), .Y(n17972) );
  AOI222XL U52361 ( .A0(net265226), .A1(n51000), .B0(n40239), .B1(n50999),
        .C0(n40321), .C1(n50998), .Y(n17948) );
  AOI222XL U52362 ( .A0(net265226), .A1(n50999), .B0(n40239), .B1(n50998),
        .C0(n40322), .C1(n50997), .Y(n17924) );
  AOI222XL U52363 ( .A0(net265207), .A1(n50998), .B0(n40240), .B1(n50997),
        .C0(n40322), .C1(n50996), .Y(n17900) );
  AOI222XL U52364 ( .A0(net265207), .A1(n50997), .B0(n40240), .B1(n50996),
        .C0(n40322), .C1(n50995), .Y(n17876) );
  AOI222XL U52365 ( .A0(net265207), .A1(n50996), .B0(n40241), .B1(n50995),
        .C0(n40323), .C1(n50994), .Y(n17852) );
  AOI222XL U52366 ( .A0(net265188), .A1(n50995), .B0(n40241), .B1(n50994),
        .C0(n40323), .C1(n50993), .Y(n17828) );
  AOI222XL U52367 ( .A0(net265188), .A1(n50994), .B0(n40241), .B1(n50993),
        .C0(n40323), .C1(n50992), .Y(n17804) );
  AOI222XL U52368 ( .A0(net265188), .A1(n50993), .B0(n40242), .B1(n50992),
        .C0(n40324), .C1(n50991), .Y(n17780) );
  AOI222XL U52369 ( .A0(net265169), .A1(n50992), .B0(n40242), .B1(n50991),
        .C0(n40324), .C1(n50990), .Y(n17756) );
  AOI222XL U52370 ( .A0(net265169), .A1(n50991), .B0(n40243), .B1(n50990),
        .C0(n40324), .C1(n50989), .Y(n17732) );
  AOI222XL U52371 ( .A0(net265169), .A1(n50990), .B0(n40243), .B1(n50989),
        .C0(n40325), .C1(n50988), .Y(n17708) );
  AOI222XL U52372 ( .A0(net265150), .A1(n50989), .B0(n40243), .B1(n50988),
        .C0(n40325), .C1(n50987), .Y(n17684) );
  AOI222XL U52373 ( .A0(net265150), .A1(n50988), .B0(n40244), .B1(n50987),
        .C0(n40325), .C1(n50986), .Y(n17660) );
  AOI222XL U52374 ( .A0(net265150), .A1(n50987), .B0(n40244), .B1(n50986),
        .C0(net217096), .C1(n50985), .Y(n17636) );
  AOI222XL U52375 ( .A0(net265131), .A1(n50986), .B0(n40245), .B1(n50985),
        .C0(n40350), .C1(n50984), .Y(n17612) );
  AOI222XL U52376 ( .A0(net265207), .A1(n50985), .B0(n40240), .B1(n50984),
        .C0(n40318), .C1(n50983), .Y(n17588) );
  AOI222XL U52377 ( .A0(net265454), .A1(n50984), .B0(n40225), .B1(n50983),
        .C0(n40326), .C1(n50982), .Y(n17564) );
  AOI222XL U52378 ( .A0(net265454), .A1(n50983), .B0(n40226), .B1(n50982),
        .C0(n40326), .C1(n50981), .Y(n17540) );
  AOI222XL U52379 ( .A0(net265454), .A1(n50982), .B0(n40226), .B1(n50981),
        .C0(n40327), .C1(n50980), .Y(n17516) );
  AOI222XL U52380 ( .A0(net265435), .A1(n50981), .B0(n40226), .B1(n50980),
        .C0(n40327), .C1(n50979), .Y(n17492) );
  AOI222XL U52381 ( .A0(net265435), .A1(n50980), .B0(n40227), .B1(n50979),
        .C0(n40327), .C1(n50978), .Y(n17468) );
  AOI222XL U52382 ( .A0(net265435), .A1(n50979), .B0(n40227), .B1(n50978),
        .C0(n40328), .C1(n50977), .Y(n17444) );
  AOI222XL U52383 ( .A0(net265416), .A1(n50978), .B0(n40228), .B1(n50977),
        .C0(n40328), .C1(n50976), .Y(n17420) );
  AOI222XL U52384 ( .A0(net265416), .A1(n50977), .B0(n40228), .B1(n50976),
        .C0(n40328), .C1(n50975), .Y(n17396) );
  AOI222XL U52385 ( .A0(net265416), .A1(n50976), .B0(n40228), .B1(n50975),
        .C0(n40329), .C1(n50974), .Y(n17372) );
  AOI222XL U52386 ( .A0(net265397), .A1(n50975), .B0(n40229), .B1(n50974),
        .C0(n40329), .C1(n50973), .Y(n17348) );
  AOI222XL U52387 ( .A0(net265397), .A1(n50974), .B0(n40229), .B1(n50973),
        .C0(n40329), .C1(n50972), .Y(n17324) );
  AOI222XL U52388 ( .A0(net265397), .A1(n50973), .B0(n40230), .B1(n50972),
        .C0(n40330), .C1(n50971), .Y(n17300) );
  AOI222XL U52389 ( .A0(net265378), .A1(n50972), .B0(n40230), .B1(n50971),
        .C0(n40330), .C1(n50970), .Y(n17276) );
  AOI222XL U52390 ( .A0(net265378), .A1(n50971), .B0(n40230), .B1(n50970),
        .C0(n40330), .C1(n50969), .Y(n17252) );
  AOI222XL U52391 ( .A0(net265378), .A1(n50970), .B0(n40231), .B1(n50969),
        .C0(n40331), .C1(n50968), .Y(n17228) );
  AOI222XL U52392 ( .A0(net265359), .A1(n50969), .B0(n40231), .B1(n50968),
        .C0(n40331), .C1(n50967), .Y(n17204) );
  AOI222XL U52393 ( .A0(net265359), .A1(n50968), .B0(n40232), .B1(n50967),
        .C0(n40331), .C1(n50966), .Y(n17180) );
  AOI222XL U52394 ( .A0(net265359), .A1(n50967), .B0(n40232), .B1(n50966),
        .C0(n40332), .C1(n50965), .Y(n17156) );
  AOI222XL U52395 ( .A0(net265340), .A1(n50966), .B0(n40232), .B1(n50965),
        .C0(n40332), .C1(n50964), .Y(n17132) );
  AOI222XL U52396 ( .A0(net265340), .A1(n50965), .B0(n40233), .B1(n50964),
        .C0(n40333), .C1(n50963), .Y(n17108) );
  AOI222XL U52397 ( .A0(net265340), .A1(n50964), .B0(n40233), .B1(n50963),
        .C0(n40333), .C1(n50962), .Y(n17084) );
  AOI222XL U52398 ( .A0(net265321), .A1(n50963), .B0(n40234), .B1(n50962),
        .C0(n40333), .C1(n50961), .Y(n17060) );
  AOI222XL U52399 ( .A0(net265321), .A1(n50962), .B0(n40234), .B1(n50961),
        .C0(n40334), .C1(n50960), .Y(n17036) );
  AOI222XL U52400 ( .A0(net265321), .A1(n50961), .B0(n40234), .B1(n50960),
        .C0(n40334), .C1(n50959), .Y(n17012) );
  AOI222XL U52401 ( .A0(net265302), .A1(n50960), .B0(n40235), .B1(n50959),
        .C0(n40334), .C1(n50958), .Y(n16988) );
  AOI222XL U52402 ( .A0(net265302), .A1(n50959), .B0(n40235), .B1(n50958),
        .C0(n40335), .C1(n50957), .Y(n16964) );
  AOI222XL U52403 ( .A0(net264960), .A1(n50958), .B0(n40256), .B1(n50957),
        .C0(n40335), .C1(n50956), .Y(n16940) );
  AOI222XL U52404 ( .A0(net264960), .A1(n50957), .B0(n40256), .B1(n50956),
        .C0(n40335), .C1(n50955), .Y(n16916) );
  AOI222XL U52405 ( .A0(net264941), .A1(n50956), .B0(n40257), .B1(n50955),
        .C0(n40336), .C1(n50954), .Y(n16892) );
  AOI222XL U52406 ( .A0(net264941), .A1(n50955), .B0(n40257), .B1(n50954),
        .C0(n40336), .C1(n50953), .Y(n16868) );
  AOI222XL U52407 ( .A0(net264941), .A1(n50954), .B0(n40257), .B1(n50953),
        .C0(n40336), .C1(n50952), .Y(n16844) );
  AOI222XL U52408 ( .A0(net264922), .A1(n50953), .B0(n40258), .B1(n50952),
        .C0(n40337), .C1(n50951), .Y(n16820) );
  AOI222XL U52409 ( .A0(net264922), .A1(n50952), .B0(n40258), .B1(n50951),
        .C0(n40337), .C1(n50950), .Y(n16796) );
  AOI222XL U52410 ( .A0(net264922), .A1(n50951), .B0(n40259), .B1(n50950),
        .C0(n40337), .C1(n50949), .Y(n16772) );
  AOI222XL U52411 ( .A0(net264903), .A1(n50950), .B0(n40259), .B1(n50949),
        .C0(n40338), .C1(n50948), .Y(n16748) );
  AOI222XL U52412 ( .A0(net264903), .A1(n50949), .B0(n40259), .B1(n50948),
        .C0(n40338), .C1(n50947), .Y(n16724) );
  AOI222XL U52413 ( .A0(net264903), .A1(n50948), .B0(n40260), .B1(n50947),
        .C0(n40339), .C1(n50946), .Y(n16700) );
  AOI222XL U52414 ( .A0(net264884), .A1(n50947), .B0(n40260), .B1(n50946),
        .C0(n40339), .C1(n50945), .Y(n16676) );
  AOI222XL U52415 ( .A0(net264884), .A1(n50946), .B0(n40261), .B1(n50945),
        .C0(n40339), .C1(n50944), .Y(n16652) );
  AOI222XL U52416 ( .A0(net264884), .A1(n50945), .B0(n40264), .B1(n50944),
        .C0(n40340), .C1(n50943), .Y(n16628) );
  AOI222XL U52417 ( .A0(net264808), .A1(n50944), .B0(n40266), .B1(n50943),
        .C0(n40340), .C1(n50942), .Y(n16604) );
  AOI222XL U52418 ( .A0(net264808), .A1(n50943), .B0(n40266), .B1(n50942),
        .C0(n40340), .C1(n50941), .Y(n16580) );
  AOI222XL U52419 ( .A0(net264808), .A1(n50942), .B0(n40265), .B1(n50941),
        .C0(n40341), .C1(n50940), .Y(n16556) );
  AOI222XL U52420 ( .A0(net264808), .A1(n50941), .B0(n40265), .B1(n50940),
        .C0(n40341), .C1(n50939), .Y(n16532) );
  AOI222XL U52421 ( .A0(net264827), .A1(n50940), .B0(n40264), .B1(n50939),
        .C0(n40341), .C1(n50938), .Y(n16508) );
  AOI222XL U52422 ( .A0(net264827), .A1(n50939), .B0(n40264), .B1(n50938),
        .C0(n40342), .C1(n50937), .Y(n16484) );
  AOI222XL U52423 ( .A0(net264846), .A1(n50938), .B0(n40264), .B1(n50937),
        .C0(n40342), .C1(n50936), .Y(n16460) );
  AOI222XL U52424 ( .A0(net264846), .A1(n50937), .B0(n40263), .B1(n50936),
        .C0(n40342), .C1(n50935), .Y(n16436) );
  AOI222XL U52425 ( .A0(net264846), .A1(n50936), .B0(n40263), .B1(n50935),
        .C0(n40343), .C1(n50934), .Y(n16412) );
  AOI222XL U52426 ( .A0(net264865), .A1(n50935), .B0(n40262), .B1(n50934),
        .C0(n40343), .C1(n50933), .Y(n16388) );
  AOI222XL U52427 ( .A0(net264865), .A1(n50934), .B0(n40262), .B1(n50933),
        .C0(n40343), .C1(n50932), .Y(n16364) );
  AOI222XL U52428 ( .A0(net264865), .A1(n50933), .B0(n40262), .B1(n50932),
        .C0(n40344), .C1(n50931), .Y(n16340) );
  AOI222XL U52429 ( .A0(net264884), .A1(n50932), .B0(n40261), .B1(n50931),
        .C0(n40344), .C1(n50930), .Y(n16316) );
  AOI222XL U52430 ( .A0(net265131), .A1(n50931), .B0(n40245), .B1(n50930),
        .C0(n40345), .C1(n50929), .Y(n16292) );
  AOI222XL U52431 ( .A0(net265112), .A1(n50930), .B0(n40246), .B1(n50929),
        .C0(n40345), .C1(n50928), .Y(n16268) );
  AOI222XL U52432 ( .A0(net265112), .A1(n50929), .B0(n40246), .B1(n50928),
        .C0(n40345), .C1(n50927), .Y(n16244) );
  AOI222XL U52433 ( .A0(net265112), .A1(n50928), .B0(n40247), .B1(n50927),
        .C0(n40346), .C1(n50926), .Y(n16220) );
  AOI222XL U52434 ( .A0(net221822), .A1(n50927), .B0(n40247), .B1(n50926),
        .C0(n40346), .C1(n50925), .Y(n16196) );
  AOI222XL U52435 ( .A0(net221812), .A1(n50926), .B0(n40247), .B1(n50925),
        .C0(n40346), .C1(n50924), .Y(n16172) );
  AOI222XL U52436 ( .A0(net221810), .A1(n50925), .B0(n40248), .B1(n50924),
        .C0(n40347), .C1(n50923), .Y(n16148) );
  AOI222XL U52437 ( .A0(net265074), .A1(n50924), .B0(n40248), .B1(n50923),
        .C0(n40347), .C1(n50922), .Y(n16124) );
  AOI222XL U52438 ( .A0(net265074), .A1(n50923), .B0(n40249), .B1(n50922),
        .C0(n40347), .C1(n50921), .Y(n16100) );
  AOI222XL U52439 ( .A0(net265074), .A1(n50922), .B0(n40249), .B1(n50921),
        .C0(n40348), .C1(n50920), .Y(n16076) );
  AOI222XL U52440 ( .A0(net265055), .A1(n50921), .B0(n40249), .B1(n50920),
        .C0(n40348), .C1(n50919), .Y(n16052) );
  AOI222XL U52441 ( .A0(net265055), .A1(n50920), .B0(n40250), .B1(n50919),
        .C0(n40348), .C1(n50918), .Y(n16028) );
  AOI222XL U52442 ( .A0(net265055), .A1(n50919), .B0(n40250), .B1(n50918),
        .C0(n40349), .C1(n50917), .Y(n16004) );
  AOI222XL U52443 ( .A0(net265036), .A1(n50918), .B0(n40251), .B1(n50917),
        .C0(n40349), .C1(n50916), .Y(n15980) );
  AOI222XL U52444 ( .A0(net265036), .A1(n50917), .B0(n40251), .B1(n50916),
        .C0(n40349), .C1(n50915), .Y(n15956) );
  AOI222XL U52445 ( .A0(net265036), .A1(n50916), .B0(n40251), .B1(n50915),
        .C0(n40382), .C1(n50914), .Y(n15932) );
  AOI222XL U52446 ( .A0(net265017), .A1(n50915), .B0(n40252), .B1(n50914),
        .C0(n40382), .C1(n50913), .Y(n15908) );
  AOI222XL U52447 ( .A0(net265017), .A1(n50914), .B0(n40252), .B1(n50913),
        .C0(n40350), .C1(n50912), .Y(n15884) );
  AOI222XL U52448 ( .A0(net265017), .A1(n50913), .B0(n40253), .B1(n50912),
        .C0(n40350), .C1(n50911), .Y(n15860) );
  AOI222XL U52449 ( .A0(net264998), .A1(n50912), .B0(n40253), .B1(n50911),
        .C0(n40350), .C1(n50910), .Y(n15836) );
  AOI222XL U52450 ( .A0(net264998), .A1(n50911), .B0(n40253), .B1(n50910),
        .C0(n40343), .C1(n50909), .Y(n15812) );
  AOI222XL U52451 ( .A0(net264998), .A1(n50910), .B0(n40254), .B1(n50909),
        .C0(net217036), .C1(n50908), .Y(n15788) );
  AOI222XL U52452 ( .A0(net264979), .A1(n50909), .B0(n40254), .B1(n50908),
        .C0(net217036), .C1(n50907), .Y(n15764) );
  AOI222XL U52453 ( .A0(net264979), .A1(n50908), .B0(n40255), .B1(n50907),
        .C0(n40351), .C1(n50906), .Y(n15740) );
  AOI222XL U52454 ( .A0(net264979), .A1(n50907), .B0(n40255), .B1(n50906),
        .C0(n40351), .C1(n50905), .Y(n15716) );
  AOI222XL U52455 ( .A0(net264960), .A1(n50906), .B0(n40255), .B1(n50905),
        .C0(n40351), .C1(n50904), .Y(n15692) );
  AOI222XL U52456 ( .A0(net265131), .A1(n50905), .B0(n40193), .B1(n50904),
        .C0(n40352), .C1(n50903), .Y(n15668) );
  AOI222XL U52457 ( .A0(net265967), .A1(n50904), .B0(n40193), .B1(n50903),
        .C0(n40352), .C1(n50902), .Y(n15644) );
  AOI222XL U52458 ( .A0(net265967), .A1(n50903), .B0(n40194), .B1(n50902),
        .C0(n40352), .C1(n50901), .Y(n15620) );
  AOI222XL U52459 ( .A0(net265967), .A1(n50902), .B0(n40194), .B1(n50901),
        .C0(n40353), .C1(n50900), .Y(n15596) );
  AOI222XL U52460 ( .A0(net265948), .A1(n50901), .B0(n40194), .B1(n50900),
        .C0(n40353), .C1(n50899), .Y(n15572) );
  AOI222XL U52461 ( .A0(net265948), .A1(n50900), .B0(n40195), .B1(n50899),
        .C0(n40353), .C1(n50898), .Y(n15548) );
  AOI222XL U52462 ( .A0(net265948), .A1(n50899), .B0(n40195), .B1(n50898),
        .C0(n40354), .C1(n50897), .Y(n15524) );
  AOI222XL U52463 ( .A0(net265929), .A1(n50898), .B0(n40196), .B1(n50897),
        .C0(n40354), .C1(n50896), .Y(n15500) );
  AOI222XL U52464 ( .A0(net265929), .A1(n50897), .B0(n40196), .B1(n50896),
        .C0(n40355), .C1(n50895), .Y(n15476) );
  AOI222XL U52465 ( .A0(net265929), .A1(n50896), .B0(n40196), .B1(n50895),
        .C0(n40355), .C1(n50894), .Y(n15452) );
  AOI222XL U52466 ( .A0(net265910), .A1(n50895), .B0(n40197), .B1(n50894),
        .C0(n40355), .C1(n50893), .Y(n15428) );
  AOI222XL U52467 ( .A0(net265910), .A1(n50894), .B0(n40197), .B1(n50893),
        .C0(n40356), .C1(n50892), .Y(n15404) );
  AOI222XL U52468 ( .A0(net265910), .A1(n50893), .B0(n40198), .B1(n50892),
        .C0(n40356), .C1(n50891), .Y(n15380) );
  AOI222XL U52469 ( .A0(net265891), .A1(n50892), .B0(n40198), .B1(n50891),
        .C0(n40356), .C1(n50890), .Y(n15356) );
  AOI222XL U52470 ( .A0(net265891), .A1(n50891), .B0(n40198), .B1(n50890),
        .C0(n40357), .C1(n50889), .Y(n15332) );
  AOI222XL U52471 ( .A0(net265872), .A1(n50890), .B0(n40199), .B1(n50889),
        .C0(n40357), .C1(n50888), .Y(n15308) );
  AOI222XL U52472 ( .A0(net265872), .A1(n50889), .B0(n40199), .B1(n50888),
        .C0(n40357), .C1(n50887), .Y(n15284) );
  AOI222XL U52473 ( .A0(net265872), .A1(n50888), .B0(n40200), .B1(n50887),
        .C0(n40358), .C1(n50886), .Y(n15260) );
  AOI222XL U52474 ( .A0(net265853), .A1(n50887), .B0(n40200), .B1(n50886),
        .C0(n40358), .C1(n50885), .Y(n15236) );
  AOI222XL U52475 ( .A0(net265853), .A1(n50886), .B0(n40200), .B1(n50885),
        .C0(n40358), .C1(n50884), .Y(n15212) );
  AOI222XL U52476 ( .A0(net265853), .A1(n50885), .B0(n40201), .B1(n50884),
        .C0(n40359), .C1(n50883), .Y(n15188) );
  AOI222XL U52477 ( .A0(net265834), .A1(n50884), .B0(n40201), .B1(n50883),
        .C0(n40359), .C1(n50882), .Y(n15164) );
  AOI222XL U52478 ( .A0(net265834), .A1(n50883), .B0(n40202), .B1(n50882),
        .C0(n40359), .C1(n50881), .Y(n15140) );
  AOI222XL U52479 ( .A0(net265834), .A1(n50882), .B0(n40202), .B1(n50881),
        .C0(n40360), .C1(n50880), .Y(n15116) );
  AOI222XL U52480 ( .A0(net265815), .A1(n50881), .B0(n40202), .B1(n50880),
        .C0(n40360), .C1(n50879), .Y(n15092) );
  AOI222XL U52481 ( .A0(net265815), .A1(n50880), .B0(n40203), .B1(n50879),
        .C0(n40377), .C1(n50878), .Y(n15068) );
  AOI222XL U52482 ( .A0(net265815), .A1(n50879), .B0(n40203), .B1(n50878),
        .C0(n40356), .C1(n50877), .Y(n15044) );
  AOI222XL U52483 ( .A0(net221892), .A1(n50877), .B0(n40184), .B1(n50876),
        .C0(n40361), .C1(n50875), .Y(n14996) );
  AOI222XL U52484 ( .A0(net221892), .A1(n50876), .B0(n40184), .B1(n50875),
        .C0(n40361), .C1(n50874), .Y(n14972) );
  AOI222XL U52485 ( .A0(net266119), .A1(n50875), .B0(n40184), .B1(n50874),
        .C0(n40361), .C1(n50873), .Y(n14948) );
  AOI222XL U52486 ( .A0(net266119), .A1(n50874), .B0(n40185), .B1(n50873),
        .C0(n40362), .C1(n50872), .Y(n14924) );
  OAI211X1 U52487 ( .A0(n32990), .A1(n42985), .B0(n14899), .C0(n14900), .Y(
        n35139) );
  AOI222XL U52488 ( .A0(net266119), .A1(n50873), .B0(n40185), .B1(n50872),
        .C0(n40362), .C1(n50871), .Y(n14900) );
  OAI211X1 U52489 ( .A0(n32982), .A1(n42987), .B0(n14875), .C0(n14876), .Y(
        n35131) );
  AOI222XL U52490 ( .A0(net266100), .A1(n50872), .B0(n40194), .B1(n50871),
        .C0(n40362), .C1(n50870), .Y(n14876) );
  OAI211X1 U52491 ( .A0(n32974), .A1(n42988), .B0(n14851), .C0(n14852), .Y(
        n35123) );
  OA22X1 U52492 ( .A0(net263767), .A1(n32958), .B0(n32966), .B1(n40052), .Y(
        n14851) );
  AOI222XL U52493 ( .A0(net266100), .A1(n50871), .B0(n40196), .B1(n50870),
        .C0(n40363), .C1(n50869), .Y(n14852) );
  OAI211X1 U52494 ( .A0(n32966), .A1(n42989), .B0(n14827), .C0(n14828), .Y(
        n35115) );
  OA22X1 U52495 ( .A0(net263501), .A1(n32950), .B0(n32958), .B1(n40052), .Y(
        n14827) );
  AOI222XL U52496 ( .A0(net266100), .A1(n50870), .B0(n40197), .B1(n50869),
        .C0(n40363), .C1(n50868), .Y(n14828) );
  OAI211X1 U52497 ( .A0(n32958), .A1(n42990), .B0(n14803), .C0(n14804), .Y(
        n35107) );
  OA22X1 U52498 ( .A0(net262969), .A1(n32942), .B0(n32950), .B1(n40051), .Y(
        n14803) );
  AOI222XL U52499 ( .A0(net266081), .A1(n50869), .B0(n40186), .B1(n50868),
        .C0(n40363), .C1(n50867), .Y(n14804) );
  OAI211X1 U52500 ( .A0(n32950), .A1(n42960), .B0(n14779), .C0(n14780), .Y(
        n35099) );
  OA22X1 U52501 ( .A0(net263805), .A1(n32934), .B0(n32942), .B1(n40051), .Y(
        n14779) );
  AOI222XL U52502 ( .A0(net266081), .A1(n50868), .B0(n40186), .B1(n50867),
        .C0(n40374), .C1(n50866), .Y(n14780) );
  OAI211X1 U52503 ( .A0(n32942), .A1(n42960), .B0(n14755), .C0(n14756), .Y(
        n35091) );
  OA22X1 U52504 ( .A0(net263805), .A1(n32926), .B0(n32934), .B1(n40050), .Y(
        n14755) );
  AOI222XL U52505 ( .A0(net266081), .A1(n50867), .B0(n40187), .B1(n50866),
        .C0(n40374), .C1(n50865), .Y(n14756) );
  OAI211X1 U52506 ( .A0(n32934), .A1(n42961), .B0(n14731), .C0(n14732), .Y(
        n35083) );
  OA22X1 U52507 ( .A0(net263824), .A1(n32918), .B0(n32926), .B1(n40050), .Y(
        n14731) );
  AOI222XL U52508 ( .A0(net266062), .A1(n50866), .B0(n40187), .B1(n50865),
        .C0(n40364), .C1(n50864), .Y(n14732) );
  OAI211X1 U52509 ( .A0(n32926), .A1(n42962), .B0(n14707), .C0(n14708), .Y(
        n35075) );
  OA22X1 U52510 ( .A0(net263824), .A1(n32910), .B0(n32918), .B1(n40049), .Y(
        n14707) );
  AOI222XL U52511 ( .A0(net266062), .A1(n50865), .B0(n40187), .B1(n50864),
        .C0(n40364), .C1(n50863), .Y(n14708) );
  OAI211X1 U52512 ( .A0(n32918), .A1(n42963), .B0(n14683), .C0(n14684), .Y(
        n35067) );
  OA22X1 U52513 ( .A0(net263824), .A1(n32902), .B0(n32910), .B1(n40049), .Y(
        n14683) );
  AOI222XL U52514 ( .A0(net266062), .A1(n50864), .B0(n40188), .B1(n50863),
        .C0(n40364), .C1(n50862), .Y(n14684) );
  OAI211X1 U52515 ( .A0(n32910), .A1(n42965), .B0(n14659), .C0(n14660), .Y(
        n35059) );
  OA22X1 U52516 ( .A0(net263843), .A1(n32894), .B0(n32902), .B1(n40048), .Y(
        n14659) );
  AOI222XL U52517 ( .A0(net266043), .A1(n50863), .B0(n40188), .B1(n50862),
        .C0(n40365), .C1(n50861), .Y(n14660) );
  OAI211X1 U52518 ( .A0(n32902), .A1(n42966), .B0(n14635), .C0(n14636), .Y(
        n35051) );
  OA22X1 U52519 ( .A0(net263843), .A1(n32886), .B0(n32894), .B1(n40048), .Y(
        n14635) );
  AOI222XL U52520 ( .A0(net266043), .A1(n50862), .B0(n40189), .B1(n50861),
        .C0(n40365), .C1(n50860), .Y(n14636) );
  OAI211X1 U52521 ( .A0(n32894), .A1(n42967), .B0(n14611), .C0(n14612), .Y(
        n35043) );
  OA22X1 U52522 ( .A0(net263862), .A1(n32878), .B0(n32886), .B1(n40047), .Y(
        n14611) );
  AOI222XL U52523 ( .A0(net266043), .A1(n50861), .B0(n40189), .B1(n50860),
        .C0(n40365), .C1(n50859), .Y(n14612) );
  OAI211X1 U52524 ( .A0(n32886), .A1(n42968), .B0(n14587), .C0(n14588), .Y(
        n35035) );
  OA22X1 U52525 ( .A0(net263862), .A1(n32870), .B0(n32878), .B1(n40047), .Y(
        n14587) );
  AOI222XL U52526 ( .A0(net266024), .A1(n50860), .B0(n40189), .B1(n50859),
        .C0(n40366), .C1(n50858), .Y(n14588) );
  OAI211X1 U52527 ( .A0(n32878), .A1(n42969), .B0(n14563), .C0(n14564), .Y(
        n35027) );
  OA22X1 U52528 ( .A0(net263064), .A1(n32862), .B0(n32870), .B1(n40092), .Y(
        n14563) );
  AOI222XL U52529 ( .A0(net266024), .A1(n50859), .B0(n40190), .B1(n50858),
        .C0(n40366), .C1(n50857), .Y(n14564) );
  OAI211X1 U52530 ( .A0(n32870), .A1(n42970), .B0(n14539), .C0(n14540), .Y(
        n35019) );
  OA22X1 U52531 ( .A0(net263064), .A1(n32854), .B0(n32862), .B1(n40092), .Y(
        n14539) );
  AOI222XL U52532 ( .A0(net266024), .A1(n50858), .B0(n40190), .B1(n50857),
        .C0(n40366), .C1(n50856), .Y(n14540) );
  OAI211X1 U52533 ( .A0(n32862), .A1(n42972), .B0(n14515), .C0(n14516), .Y(
        n35011) );
  OA22X1 U52534 ( .A0(net263083), .A1(n32846), .B0(n32854), .B1(n40091), .Y(
        n14515) );
  AOI222XL U52535 ( .A0(net266005), .A1(n50857), .B0(n40191), .B1(n50856),
        .C0(n40367), .C1(n50855), .Y(n14516) );
  OAI211X1 U52536 ( .A0(n32854), .A1(n42973), .B0(n14491), .C0(n14492), .Y(
        n35003) );
  OA22X1 U52537 ( .A0(net263083), .A1(n32838), .B0(n32846), .B1(n40091), .Y(
        n14491) );
  AOI222XL U52538 ( .A0(net266005), .A1(n50856), .B0(n40191), .B1(n50855),
        .C0(n40367), .C1(n50854), .Y(n14492) );
  OAI211X1 U52539 ( .A0(n32846), .A1(n42974), .B0(n14467), .C0(n14468), .Y(
        n34995) );
  OA22X1 U52540 ( .A0(net263102), .A1(n32830), .B0(n32838), .B1(n40090), .Y(
        n14467) );
  AOI222XL U52541 ( .A0(net266005), .A1(n50855), .B0(n40191), .B1(n50854),
        .C0(n40367), .C1(n50853), .Y(n14468) );
  OAI211X1 U52542 ( .A0(n32838), .A1(n42975), .B0(n14443), .C0(n14444), .Y(
        n34987) );
  OA22X1 U52543 ( .A0(net263102), .A1(n32822), .B0(n32830), .B1(n40090), .Y(
        n14443) );
  AOI222XL U52544 ( .A0(net265321), .A1(n50854), .B0(n40192), .B1(n50853),
        .C0(n40368), .C1(n50852), .Y(n14444) );
  OAI211X1 U52545 ( .A0(n32830), .A1(n42887), .B0(n14419), .C0(n14420), .Y(
        n34979) );
  OA22X1 U52546 ( .A0(net263121), .A1(n32814), .B0(n32822), .B1(n40089), .Y(
        n14419) );
  AOI222XL U52547 ( .A0(net265644), .A1(n50853), .B0(n40192), .B1(n50852),
        .C0(n40368), .C1(n50851), .Y(n14420) );
  OAI211X1 U52548 ( .A0(n32822), .A1(n42880), .B0(n14395), .C0(n14396), .Y(
        n34971) );
  OA22X1 U52549 ( .A0(net263121), .A1(n32806), .B0(n32814), .B1(n40089), .Y(
        n14395) );
  AOI222XL U52550 ( .A0(net265682), .A1(n50852), .B0(n40193), .B1(n50851),
        .C0(n40368), .C1(n50850), .Y(n14396) );
  OAI211X1 U52551 ( .A0(n32814), .A1(n42881), .B0(n14371), .C0(n14372), .Y(
        n34963) );
  OA22X1 U52552 ( .A0(net263140), .A1(n32798), .B0(n32806), .B1(n40088), .Y(
        n14371) );
  AOI222XL U52553 ( .A0(net265644), .A1(n50851), .B0(n40214), .B1(n50850),
        .C0(n40369), .C1(n50849), .Y(n14372) );
  OAI211X1 U52554 ( .A0(n32806), .A1(n42882), .B0(n14347), .C0(n14348), .Y(
        n34955) );
  OA22X1 U52555 ( .A0(net263140), .A1(n32790), .B0(n32798), .B1(n40088), .Y(
        n14347) );
  AOI222XL U52556 ( .A0(net265625), .A1(n50850), .B0(n40215), .B1(n50849),
        .C0(n40369), .C1(n50848), .Y(n14348) );
  OAI211X1 U52557 ( .A0(n32798), .A1(n42884), .B0(n14323), .C0(n14324), .Y(
        n34947) );
  OA22X1 U52558 ( .A0(net263140), .A1(n32782), .B0(n32790), .B1(n40087), .Y(
        n14323) );
  AOI222XL U52559 ( .A0(net265625), .A1(n50849), .B0(n40215), .B1(n50848),
        .C0(n40369), .C1(n50847), .Y(n14324) );
  OAI211X1 U52560 ( .A0(n32790), .A1(n42885), .B0(n14299), .C0(n14300), .Y(
        n34939) );
  OA22X1 U52561 ( .A0(net263159), .A1(n32774), .B0(n32782), .B1(n40087), .Y(
        n14299) );
  AOI222XL U52562 ( .A0(net265625), .A1(n50848), .B0(n40216), .B1(n50847),
        .C0(n40370), .C1(n50846), .Y(n14300) );
  OAI211X1 U52563 ( .A0(n32782), .A1(n42886), .B0(n14275), .C0(n14276), .Y(
        n34931) );
  OA22X1 U52564 ( .A0(net263159), .A1(n32766), .B0(n32774), .B1(n40086), .Y(
        n14275) );
  AOI222XL U52565 ( .A0(net265606), .A1(n50847), .B0(n40216), .B1(n50846),
        .C0(n40370), .C1(n50845), .Y(n14276) );
  OAI211X1 U52566 ( .A0(n32774), .A1(n42887), .B0(n14251), .C0(n14252), .Y(
        n34923) );
  OA22X1 U52567 ( .A0(net263178), .A1(n32758), .B0(n32766), .B1(n40086), .Y(
        n14251) );
  AOI222XL U52568 ( .A0(net265606), .A1(n50846), .B0(n40216), .B1(n50845),
        .C0(n40371), .C1(n50844), .Y(n14252) );
  OAI211X1 U52569 ( .A0(n32766), .A1(n42888), .B0(n14227), .C0(n14228), .Y(
        n34915) );
  OA22X1 U52570 ( .A0(net263178), .A1(n32750), .B0(n32758), .B1(n40085), .Y(
        n14227) );
  AOI222XL U52571 ( .A0(net265606), .A1(n50845), .B0(n40217), .B1(n50844),
        .C0(n40371), .C1(n50843), .Y(n14228) );
  OAI211X1 U52572 ( .A0(n32758), .A1(n42889), .B0(n14203), .C0(n14204), .Y(
        n34907) );
  OA22X1 U52573 ( .A0(net218420), .A1(n32742), .B0(n32750), .B1(n40085), .Y(
        n14203) );
  AOI222XL U52574 ( .A0(net265587), .A1(n50844), .B0(n40217), .B1(n50843),
        .C0(n40371), .C1(n50842), .Y(n14204) );
  OAI211X1 U52575 ( .A0(n32750), .A1(n42891), .B0(n14179), .C0(n14180), .Y(
        n34899) );
  OA22X1 U52576 ( .A0(net262931), .A1(n32734), .B0(n32742), .B1(n40100), .Y(
        n14179) );
  AOI222XL U52577 ( .A0(net265587), .A1(n50843), .B0(n40218), .B1(n50842),
        .C0(n40372), .C1(n50841), .Y(n14180) );
  OAI211X1 U52578 ( .A0(n32742), .A1(n42892), .B0(n14155), .C0(n14156), .Y(
        n34891) );
  OA22X1 U52579 ( .A0(net262931), .A1(n32726), .B0(n32734), .B1(n40100), .Y(
        n14155) );
  AOI222XL U52580 ( .A0(net265587), .A1(n50842), .B0(n40218), .B1(n50841),
        .C0(n40372), .C1(n50840), .Y(n14156) );
  OAI211X1 U52581 ( .A0(n32734), .A1(n42893), .B0(n14131), .C0(n14132), .Y(
        n34883) );
  OA22X1 U52582 ( .A0(net262950), .A1(n32718), .B0(n32726), .B1(n40099), .Y(
        n14131) );
  AOI222XL U52583 ( .A0(net265568), .A1(n50841), .B0(n40218), .B1(n50840),
        .C0(n40372), .C1(n50839), .Y(n14132) );
  OAI211X1 U52584 ( .A0(n32726), .A1(n42894), .B0(n14107), .C0(n14108), .Y(
        n34875) );
  OA22X1 U52585 ( .A0(net262950), .A1(n32710), .B0(n32718), .B1(n40099), .Y(
        n14107) );
  AOI222XL U52586 ( .A0(net265568), .A1(n50840), .B0(n40219), .B1(n50839),
        .C0(n40373), .C1(n50838), .Y(n14108) );
  OAI211X1 U52587 ( .A0(n32718), .A1(n42871), .B0(n14083), .C0(n14084), .Y(
        n34867) );
  OA22X1 U52588 ( .A0(net262969), .A1(n32702), .B0(n32710), .B1(n40098), .Y(
        n14083) );
  AOI222XL U52589 ( .A0(net265568), .A1(n50839), .B0(n40219), .B1(n50838),
        .C0(n40373), .C1(n50837), .Y(n14084) );
  OAI211X1 U52590 ( .A0(n32710), .A1(n42864), .B0(n14059), .C0(n14060), .Y(
        n34859) );
  OA22X1 U52591 ( .A0(net262969), .A1(n32694), .B0(n32702), .B1(n40098), .Y(
        n14059) );
  AOI222XL U52592 ( .A0(net265549), .A1(n50838), .B0(n40220), .B1(n50837),
        .C0(n40373), .C1(n50836), .Y(n14060) );
  OAI211X1 U52593 ( .A0(n32702), .A1(n42865), .B0(n14035), .C0(n14036), .Y(
        n34851) );
  OA22X1 U52594 ( .A0(net262988), .A1(n32686), .B0(n32694), .B1(n40097), .Y(
        n14035) );
  AOI222XL U52595 ( .A0(net265549), .A1(n50837), .B0(n40220), .B1(n50836),
        .C0(n40374), .C1(n50835), .Y(n14036) );
  OAI211X1 U52596 ( .A0(n32694), .A1(n42866), .B0(n14011), .C0(n14012), .Y(
        n34843) );
  OA22X1 U52597 ( .A0(net262988), .A1(n32678), .B0(n32686), .B1(n40097), .Y(
        n14011) );
  AOI222XL U52598 ( .A0(net265530), .A1(n50836), .B0(n40220), .B1(n50835),
        .C0(n40374), .C1(n50834), .Y(n14012) );
  OAI211X1 U52599 ( .A0(n32686), .A1(n42868), .B0(n13987), .C0(n13988), .Y(
        n34835) );
  OA22X1 U52600 ( .A0(net262988), .A1(n32670), .B0(n32678), .B1(n40096), .Y(
        n13987) );
  AOI222XL U52601 ( .A0(net265530), .A1(n50835), .B0(n40221), .B1(n50834),
        .C0(n40374), .C1(n50833), .Y(n13988) );
  OAI211X1 U52602 ( .A0(n32678), .A1(n42869), .B0(n13963), .C0(n13964), .Y(
        n34827) );
  OA22X1 U52603 ( .A0(net263007), .A1(n32662), .B0(n32670), .B1(n40096), .Y(
        n13963) );
  AOI222XL U52604 ( .A0(net265530), .A1(n50834), .B0(n40221), .B1(n50833),
        .C0(n40375), .C1(n50832), .Y(n13964) );
  OAI211X1 U52605 ( .A0(n32670), .A1(n42870), .B0(n13939), .C0(n13940), .Y(
        n34819) );
  OA22X1 U52606 ( .A0(net263007), .A1(n32654), .B0(n32662), .B1(n40095), .Y(
        n13939) );
  AOI222XL U52607 ( .A0(net265511), .A1(n50833), .B0(n40222), .B1(n50832),
        .C0(n40375), .C1(n50831), .Y(n13940) );
  OAI211X1 U52608 ( .A0(n32662), .A1(n42871), .B0(n13915), .C0(n13916), .Y(
        n34811) );
  OA22X1 U52609 ( .A0(net263026), .A1(n32646), .B0(n32654), .B1(n40095), .Y(
        n13915) );
  AOI222XL U52610 ( .A0(net265511), .A1(n50832), .B0(n40222), .B1(n50831),
        .C0(n40375), .C1(n50830), .Y(n13916) );
  OAI211X1 U52611 ( .A0(n32654), .A1(n42872), .B0(n13891), .C0(n13892), .Y(
        n34803) );
  OA22X1 U52612 ( .A0(net263026), .A1(n32638), .B0(n32646), .B1(n40094), .Y(
        n13891) );
  AOI222XL U52613 ( .A0(net265511), .A1(n50831), .B0(n40222), .B1(n50830),
        .C0(n40376), .C1(n50829), .Y(n13892) );
  OAI211X1 U52614 ( .A0(n32646), .A1(n42873), .B0(n13867), .C0(n13868), .Y(
        n34795) );
  OA22X1 U52615 ( .A0(net263045), .A1(n32630), .B0(n32638), .B1(n40094), .Y(
        n13867) );
  AOI222XL U52616 ( .A0(net265492), .A1(n50830), .B0(n40223), .B1(n50829),
        .C0(n40376), .C1(n50828), .Y(n13868) );
  OAI211X1 U52617 ( .A0(n32638), .A1(n42875), .B0(n13843), .C0(n13844), .Y(
        n34787) );
  OA22X1 U52618 ( .A0(net263045), .A1(n32622), .B0(n32630), .B1(n40093), .Y(
        n13843) );
  AOI222XL U52619 ( .A0(net265492), .A1(n50829), .B0(n40223), .B1(n50828),
        .C0(n40377), .C1(n50827), .Y(n13844) );
  OAI211X1 U52620 ( .A0(n32630), .A1(n42876), .B0(n13819), .C0(n13820), .Y(
        n34779) );
  OA22X1 U52621 ( .A0(net263064), .A1(n32614), .B0(n32622), .B1(n40093), .Y(
        n13819) );
  AOI222XL U52622 ( .A0(net265492), .A1(n50828), .B0(n40224), .B1(n50827),
        .C0(n40377), .C1(n50826), .Y(n13820) );
  OAI211X1 U52623 ( .A0(n32622), .A1(n42877), .B0(n13795), .C0(n13796), .Y(
        n34771) );
  OA22X1 U52624 ( .A0(net263330), .A1(n32606), .B0(n32614), .B1(n40077), .Y(
        n13795) );
  AOI222XL U52625 ( .A0(net265473), .A1(n50827), .B0(n40224), .B1(n50826),
        .C0(n40377), .C1(n50825), .Y(n13796) );
  OAI211X1 U52626 ( .A0(n32614), .A1(n42878), .B0(n13771), .C0(n13772), .Y(
        n34763) );
  OA22X1 U52627 ( .A0(net263349), .A1(n32598), .B0(n32606), .B1(n40077), .Y(
        n13771) );
  AOI222XL U52628 ( .A0(net265473), .A1(n50826), .B0(n40224), .B1(n50825),
        .C0(n40378), .C1(n50824), .Y(n13772) );
  OAI211X1 U52629 ( .A0(n32606), .A1(n42927), .B0(n13747), .C0(n13748), .Y(
        n34755) );
  OA22X1 U52630 ( .A0(net263349), .A1(n32590), .B0(n32598), .B1(n40076), .Y(
        n13747) );
  AOI222XL U52631 ( .A0(net265549), .A1(n50825), .B0(n40203), .B1(n50824),
        .C0(n40378), .C1(n50823), .Y(n13748) );
  OAI211X1 U52632 ( .A0(n32598), .A1(n42912), .B0(n13723), .C0(n13724), .Y(
        n34747) );
  OA22X1 U52633 ( .A0(net263368), .A1(n32582), .B0(n32590), .B1(n40076), .Y(
        n13723) );
  AOI222XL U52634 ( .A0(net265796), .A1(n50824), .B0(n40204), .B1(n50823),
        .C0(n40378), .C1(n50822), .Y(n13724) );
  OAI211X1 U52635 ( .A0(n32590), .A1(n42913), .B0(n13699), .C0(n13700), .Y(
        n34739) );
  OA22X1 U52636 ( .A0(net263368), .A1(n32574), .B0(n32582), .B1(n40075), .Y(
        n13699) );
  AOI222XL U52637 ( .A0(net265796), .A1(n50823), .B0(n40204), .B1(n50822),
        .C0(n40379), .C1(n50821), .Y(n13700) );
  OAI211X1 U52638 ( .A0(n32582), .A1(n42915), .B0(n13675), .C0(n13676), .Y(
        n34731) );
  OA22X1 U52639 ( .A0(net263368), .A1(n32566), .B0(n32574), .B1(n40075), .Y(
        n13675) );
  AOI222XL U52640 ( .A0(net265796), .A1(n50822), .B0(n40205), .B1(n50821),
        .C0(n40379), .C1(n50820), .Y(n13676) );
  OAI211X1 U52641 ( .A0(n32574), .A1(n42916), .B0(n13651), .C0(n13652), .Y(
        n34723) );
  OA22X1 U52642 ( .A0(net263387), .A1(n32558), .B0(n32566), .B1(n40074), .Y(
        n13651) );
  AOI222XL U52643 ( .A0(net265777), .A1(n50821), .B0(n40205), .B1(n50820),
        .C0(n40379), .C1(n50819), .Y(n13652) );
  OAI211X1 U52644 ( .A0(n32566), .A1(n42917), .B0(n13627), .C0(n13628), .Y(
        n34715) );
  OA22X1 U52645 ( .A0(net263387), .A1(n32550), .B0(n32558), .B1(n40074), .Y(
        n13627) );
  AOI222XL U52646 ( .A0(net265777), .A1(n50820), .B0(n40205), .B1(n50819),
        .C0(n40380), .C1(n50818), .Y(n13628) );
  OAI211X1 U52647 ( .A0(n32558), .A1(n42918), .B0(n13603), .C0(n13604), .Y(
        n34707) );
  OA22X1 U52648 ( .A0(net263406), .A1(n32542), .B0(n32550), .B1(n40073), .Y(
        n13603) );
  AOI222XL U52649 ( .A0(net265777), .A1(n50819), .B0(n40206), .B1(n50818),
        .C0(n40380), .C1(n50817), .Y(n13604) );
  OAI211X1 U52650 ( .A0(n32550), .A1(n42919), .B0(n13579), .C0(n13580), .Y(
        n34699) );
  OA22X1 U52651 ( .A0(net263406), .A1(n32534), .B0(n32542), .B1(n40073), .Y(
        n13579) );
  AOI222XL U52652 ( .A0(net265758), .A1(n50818), .B0(n40206), .B1(n50817),
        .C0(n40380), .C1(n50816), .Y(n13580) );
  OAI211X1 U52653 ( .A0(n32542), .A1(n42920), .B0(n13555), .C0(n13556), .Y(
        n34691) );
  OA22X1 U52654 ( .A0(net218422), .A1(n32526), .B0(n32534), .B1(n40072), .Y(
        n13555) );
  AOI222XL U52655 ( .A0(net265758), .A1(n50817), .B0(n40207), .B1(n50816),
        .C0(n40381), .C1(n50815), .Y(n13556) );
  OAI211X1 U52656 ( .A0(n32534), .A1(n42922), .B0(n13531), .C0(n13532), .Y(
        n34683) );
  OA22X1 U52657 ( .A0(net218410), .A1(n32518), .B0(n32526), .B1(n40072), .Y(
        n13531) );
  AOI222XL U52658 ( .A0(net265758), .A1(n50816), .B0(n40207), .B1(n50815),
        .C0(n40381), .C1(n50814), .Y(n13532) );
  OAI211X1 U52659 ( .A0(n32526), .A1(n42923), .B0(n13507), .C0(n13508), .Y(
        n34675) );
  OA22X1 U52660 ( .A0(net263444), .A1(n32510), .B0(n32518), .B1(n40071), .Y(
        n13507) );
  AOI222XL U52661 ( .A0(net265739), .A1(n50815), .B0(n40207), .B1(n50814),
        .C0(n40381), .C1(n50813), .Y(n13508) );
  OAI211X1 U52662 ( .A0(n32518), .A1(n42924), .B0(n13483), .C0(n13484), .Y(
        n34667) );
  OA22X1 U52663 ( .A0(net263444), .A1(n32502), .B0(n32510), .B1(n40071), .Y(
        n13483) );
  AOI222XL U52664 ( .A0(net265739), .A1(n50814), .B0(n40208), .B1(n50813),
        .C0(n40382), .C1(n50812), .Y(n13484) );
  OAI211X1 U52665 ( .A0(n32510), .A1(n42925), .B0(n13459), .C0(n13460), .Y(
        n34659) );
  OA22X1 U52666 ( .A0(net263444), .A1(n32494), .B0(n32502), .B1(n40070), .Y(
        n13459) );
  AOI222XL U52667 ( .A0(net265739), .A1(n50813), .B0(n40208), .B1(n50812),
        .C0(n40382), .C1(n50811), .Y(n13460) );
  OAI211X1 U52668 ( .A0(n32502), .A1(n42926), .B0(n13435), .C0(n13436), .Y(
        n34651) );
  OA22X1 U52669 ( .A0(net263463), .A1(n32486), .B0(n32494), .B1(n40070), .Y(
        n13435) );
  AOI222XL U52670 ( .A0(net265720), .A1(n50812), .B0(n40209), .B1(n50811),
        .C0(n40383), .C1(n50810), .Y(n13436) );
  OAI211X1 U52671 ( .A0(n32494), .A1(n42927), .B0(n13411), .C0(n13412), .Y(
        n34643) );
  OA22X1 U52672 ( .A0(net261943), .A1(n32478), .B0(n32486), .B1(n40084), .Y(
        n13411) );
  AOI222XL U52673 ( .A0(net265720), .A1(n50811), .B0(n40209), .B1(n50810),
        .C0(n40383), .C1(n50809), .Y(n13412) );
  OAI211X1 U52674 ( .A0(n32486), .A1(n42896), .B0(n13387), .C0(n13388), .Y(
        n34635) );
  OA22X1 U52675 ( .A0(net263216), .A1(n32470), .B0(n32478), .B1(n40084), .Y(
        n13387) );
  AOI222XL U52676 ( .A0(net265720), .A1(n50810), .B0(n40210), .B1(n50809),
        .C0(n40383), .C1(n50808), .Y(n13388) );
  OAI211X1 U52677 ( .A0(n32478), .A1(n42897), .B0(n13363), .C0(n13364), .Y(
        n34627) );
  OA22X1 U52678 ( .A0(net263216), .A1(n32462), .B0(n32470), .B1(n40083), .Y(
        n13363) );
  AOI222XL U52679 ( .A0(net265701), .A1(n50809), .B0(n40210), .B1(n50808),
        .C0(n40384), .C1(n50807), .Y(n13364) );
  OAI211X1 U52680 ( .A0(n32470), .A1(n42898), .B0(n13339), .C0(n13340), .Y(
        n34619) );
  OA22X1 U52681 ( .A0(net263216), .A1(n32454), .B0(n32462), .B1(n40083), .Y(
        n13339) );
  AOI222XL U52682 ( .A0(net265701), .A1(n50808), .B0(n40210), .B1(n50807),
        .C0(n40384), .C1(n50806), .Y(n13340) );
  OAI211X1 U52683 ( .A0(n32462), .A1(n42900), .B0(n13315), .C0(n13316), .Y(
        n34611) );
  OA22X1 U52684 ( .A0(net263235), .A1(n32446), .B0(n32454), .B1(n40082), .Y(
        n13315) );
  AOI222XL U52685 ( .A0(net265701), .A1(n50807), .B0(n40211), .B1(n50806),
        .C0(n40384), .C1(n50805), .Y(n13316) );
  OAI211X1 U52686 ( .A0(n32454), .A1(n42901), .B0(n13291), .C0(n13292), .Y(
        n34603) );
  OA22X1 U52687 ( .A0(net263235), .A1(n32438), .B0(n32446), .B1(n40082), .Y(
        n13291) );
  AOI222XL U52688 ( .A0(net265682), .A1(n50806), .B0(n40211), .B1(n50805),
        .C0(n40385), .C1(n50804), .Y(n13292) );
  OAI211X1 U52689 ( .A0(n32446), .A1(n42902), .B0(n13267), .C0(n13268), .Y(
        n34595) );
  OA22X1 U52690 ( .A0(net263254), .A1(n32430), .B0(n32438), .B1(n40081), .Y(
        n13267) );
  AOI222XL U52691 ( .A0(net265682), .A1(n50805), .B0(n40212), .B1(n50804),
        .C0(n40385), .C1(n50803), .Y(n13268) );
  OAI211X1 U52692 ( .A0(n32438), .A1(n42903), .B0(n13243), .C0(n13244), .Y(
        n34587) );
  OA22X1 U52693 ( .A0(net263254), .A1(n32422), .B0(n32430), .B1(n40081), .Y(
        n13243) );
  AOI222XL U52694 ( .A0(net265682), .A1(n50804), .B0(n40212), .B1(n50803),
        .C0(n40385), .C1(n50802), .Y(n13244) );
  OAI211X1 U52695 ( .A0(n32430), .A1(n42904), .B0(n13219), .C0(n13220), .Y(
        n34579) );
  OA22X1 U52696 ( .A0(net218404), .A1(n32414), .B0(n32422), .B1(n40080), .Y(
        n13219) );
  AOI222XL U52697 ( .A0(net265226), .A1(n50803), .B0(n40212), .B1(n50802),
        .C0(net217058), .C1(n50801), .Y(n13220) );
  OAI211X1 U52698 ( .A0(n32422), .A1(n42905), .B0(n13195), .C0(n13196), .Y(
        n34571) );
  OA22X1 U52699 ( .A0(net218316), .A1(n32406), .B0(n32414), .B1(n40079), .Y(
        n13195) );
  AOI222XL U52700 ( .A0(net265169), .A1(n50802), .B0(n40213), .B1(n50801),
        .C0(net217032), .C1(n50800), .Y(n13196) );
  OAI211X1 U52701 ( .A0(n32414), .A1(n42907), .B0(n13171), .C0(n13172), .Y(
        n34563) );
  AOI222XL U52702 ( .A0(net265188), .A1(n50801), .B0(n40213), .B1(n50800),
        .C0(net217054), .C1(n50799), .Y(n13172) );
  OAI211X1 U52703 ( .A0(n32406), .A1(n42908), .B0(n13147), .C0(n13148), .Y(
        n34555) );
  AOI222XL U52704 ( .A0(net265644), .A1(n50800), .B0(n40214), .B1(n50799),
        .C0(n40381), .C1(n50798), .Y(n13148) );
  OAI211X1 U52705 ( .A0(n34423), .A1(n42911), .B0(n13031), .C0(n50080), .Y(
        n34519) );
  OAI222XL U52706 ( .A0(net266654), .A1(n9664), .B0(n40159), .B1(n9663), .C0(
        n40292), .C1(n34431), .Y(n13033) );
  CLKINVX1 U52707 ( .A(n19152), .Y(n49566) );
  OAI222XL U52708 ( .A0(net266402), .A1(n34431), .B0(n40174), .B1(n34423),
        .C0(n40303), .C1(n41806), .Y(n19152) );
  OAI222XL U52709 ( .A0(net266402), .A1(n34423), .B0(n40174), .B1(n41806),
        .C0(n40303), .C1(n41807), .Y(n19128) );
  OAI211X1 U52710 ( .A0(n34424), .A1(n42911), .B0(n13028), .C0(n50081), .Y(
        n34518) );
  OAI222XL U52711 ( .A0(net266654), .A1(n9662), .B0(n40159), .B1(n9661), .C0(
        n40292), .C1(n34432), .Y(n13030) );
  CLKINVX1 U52712 ( .A(n19179), .Y(n49558) );
  OAI222XL U52713 ( .A0(net266255), .A1(n9661), .B0(n40167), .B1(n34432), .C0(
        n40286), .C1(n34424), .Y(n19179) );
  AOI222XL U52714 ( .A0(net265302), .A1(n49513), .B0(net218130), .B1(n50796),
        .C0(net217108), .C1(n50795), .Y(n18218) );
  AOI222XL U52715 ( .A0(net265283), .A1(n50796), .B0(n40189), .B1(n50795),
        .C0(n40318), .C1(n50794), .Y(n18194) );
  AOI222XL U52716 ( .A0(net265283), .A1(n50795), .B0(n40216), .B1(n50794),
        .C0(n40318), .C1(n50793), .Y(n18170) );
  AOI222XL U52717 ( .A0(net265283), .A1(n50794), .B0(n40236), .B1(n50793),
        .C0(n40318), .C1(n50792), .Y(n18146) );
  AOI222XL U52718 ( .A0(net265264), .A1(n50793), .B0(n40236), .B1(n50792),
        .C0(n40319), .C1(n50791), .Y(n18122) );
  AOI222XL U52719 ( .A0(net265264), .A1(n50792), .B0(n40237), .B1(n50791),
        .C0(n40319), .C1(n50790), .Y(n18098) );
  AOI222XL U52720 ( .A0(net265264), .A1(n50791), .B0(n40237), .B1(n50790),
        .C0(n40319), .C1(n50789), .Y(n18074) );
  AOI222XL U52721 ( .A0(net265245), .A1(n50790), .B0(n40237), .B1(n50789),
        .C0(n40320), .C1(n50788), .Y(n18050) );
  AOI222XL U52722 ( .A0(net265245), .A1(n50789), .B0(n40238), .B1(n50788),
        .C0(n40320), .C1(n50787), .Y(n18026) );
  AOI222XL U52723 ( .A0(net265245), .A1(n50788), .B0(n40238), .B1(n50787),
        .C0(n40320), .C1(n50786), .Y(n18002) );
  AOI222XL U52724 ( .A0(net265226), .A1(n50787), .B0(n40239), .B1(n50786),
        .C0(n40321), .C1(n50785), .Y(n17978) );
  AOI222XL U52725 ( .A0(net265226), .A1(n50786), .B0(n40239), .B1(n50785),
        .C0(n40321), .C1(n50784), .Y(n17954) );
  AOI222XL U52726 ( .A0(net265226), .A1(n50785), .B0(n40239), .B1(n50784),
        .C0(n40321), .C1(n50783), .Y(n17930) );
  AOI222XL U52727 ( .A0(net265207), .A1(n50784), .B0(n40240), .B1(n50783),
        .C0(n40322), .C1(n50782), .Y(n17906) );
  AOI222XL U52728 ( .A0(net265207), .A1(n50783), .B0(n40240), .B1(n50782),
        .C0(n40322), .C1(n50781), .Y(n17882) );
  AOI222XL U52729 ( .A0(net265207), .A1(n50782), .B0(n40241), .B1(n50781),
        .C0(n40323), .C1(n50780), .Y(n17858) );
  AOI222XL U52730 ( .A0(net265188), .A1(n50781), .B0(n40241), .B1(n50780),
        .C0(n40323), .C1(n50779), .Y(n17834) );
  AOI222XL U52731 ( .A0(net265188), .A1(n50780), .B0(n40241), .B1(n50779),
        .C0(n40323), .C1(n50778), .Y(n17810) );
  AOI222XL U52732 ( .A0(net265188), .A1(n50779), .B0(n40242), .B1(n50778),
        .C0(n40324), .C1(n50777), .Y(n17786) );
  AOI222XL U52733 ( .A0(net265169), .A1(n50778), .B0(n40242), .B1(n50777),
        .C0(n40324), .C1(n50776), .Y(n17762) );
  AOI222XL U52734 ( .A0(net265169), .A1(n50777), .B0(n40243), .B1(n50776),
        .C0(n40324), .C1(n50775), .Y(n17738) );
  AOI222XL U52735 ( .A0(net265169), .A1(n50776), .B0(n40243), .B1(n50775),
        .C0(n40325), .C1(n50774), .Y(n17714) );
  AOI222XL U52736 ( .A0(net265150), .A1(n50775), .B0(n40243), .B1(n50774),
        .C0(n40325), .C1(n50773), .Y(n17690) );
  AOI222XL U52737 ( .A0(net265150), .A1(n50774), .B0(n40244), .B1(n50773),
        .C0(n40325), .C1(n50772), .Y(n17666) );
  AOI222XL U52738 ( .A0(net265150), .A1(n50773), .B0(n40244), .B1(n50772),
        .C0(n40348), .C1(n50771), .Y(n17642) );
  AOI222XL U52739 ( .A0(net265131), .A1(n50772), .B0(n40245), .B1(n50771),
        .C0(n40319), .C1(n50770), .Y(n17618) );
  AOI222XL U52740 ( .A0(net265131), .A1(n50771), .B0(n40245), .B1(n50770),
        .C0(n40350), .C1(n50769), .Y(n17594) );
  AOI222XL U52741 ( .A0(net265473), .A1(n50770), .B0(n40225), .B1(n50769),
        .C0(n40326), .C1(n50768), .Y(n17570) );
  AOI222XL U52742 ( .A0(net265454), .A1(n50769), .B0(n40225), .B1(n50768),
        .C0(n40326), .C1(n50767), .Y(n17546) );
  AOI222XL U52743 ( .A0(net265454), .A1(n50768), .B0(n40226), .B1(n50767),
        .C0(n40326), .C1(n50766), .Y(n17522) );
  AOI222XL U52744 ( .A0(net265454), .A1(n50767), .B0(n40226), .B1(n50766),
        .C0(n40327), .C1(n50765), .Y(n17498) );
  AOI222XL U52745 ( .A0(net265435), .A1(n50766), .B0(n40227), .B1(n50765),
        .C0(n40327), .C1(n50764), .Y(n17474) );
  AOI222XL U52746 ( .A0(net265435), .A1(n50765), .B0(n40227), .B1(n50764),
        .C0(n40328), .C1(n50763), .Y(n17450) );
  AOI222XL U52747 ( .A0(net265435), .A1(n50764), .B0(n40227), .B1(n50763),
        .C0(n40328), .C1(n50762), .Y(n17426) );
  AOI222XL U52748 ( .A0(net265416), .A1(n50763), .B0(n40228), .B1(n50762),
        .C0(n40328), .C1(n50761), .Y(n17402) );
  AOI222XL U52749 ( .A0(net265416), .A1(n50762), .B0(n40228), .B1(n50761),
        .C0(n40329), .C1(n50760), .Y(n17378) );
  AOI222XL U52750 ( .A0(net265416), .A1(n50761), .B0(n40229), .B1(n50760),
        .C0(n40329), .C1(n50759), .Y(n17354) );
  AOI222XL U52751 ( .A0(net265397), .A1(n50760), .B0(n40229), .B1(n50759),
        .C0(n40329), .C1(n50758), .Y(n17330) );
  AOI222XL U52752 ( .A0(net265397), .A1(n50759), .B0(n40229), .B1(n50758),
        .C0(n40330), .C1(n50757), .Y(n17306) );
  AOI222XL U52753 ( .A0(net265397), .A1(n50758), .B0(n40230), .B1(n50757),
        .C0(n40330), .C1(n50756), .Y(n17282) );
  AOI222XL U52754 ( .A0(net265378), .A1(n50757), .B0(n40230), .B1(n50756),
        .C0(n40330), .C1(n50755), .Y(n17258) );
  AOI222XL U52755 ( .A0(net265378), .A1(n50756), .B0(n40231), .B1(n50755),
        .C0(n40331), .C1(n50754), .Y(n17234) );
  AOI222XL U52756 ( .A0(net265359), .A1(n50755), .B0(n40231), .B1(n50754),
        .C0(n40331), .C1(n50753), .Y(n17210) );
  AOI222XL U52757 ( .A0(net265359), .A1(n50754), .B0(n40232), .B1(n50753),
        .C0(n40331), .C1(n50752), .Y(n17186) );
  AOI222XL U52758 ( .A0(net265359), .A1(n50753), .B0(n40232), .B1(n50752),
        .C0(n40332), .C1(n50751), .Y(n17162) );
  AOI222XL U52759 ( .A0(net265340), .A1(n50752), .B0(n40232), .B1(n50751),
        .C0(n40332), .C1(n50750), .Y(n17138) );
  AOI222XL U52760 ( .A0(net265340), .A1(n50751), .B0(n40233), .B1(n50750),
        .C0(n40332), .C1(n50749), .Y(n17114) );
  AOI222XL U52761 ( .A0(net265340), .A1(n50750), .B0(n40233), .B1(n50749),
        .C0(n40333), .C1(n50748), .Y(n17090) );
  AOI222XL U52762 ( .A0(net265321), .A1(n50749), .B0(n40234), .B1(n50748),
        .C0(n40333), .C1(n50747), .Y(n17066) );
  AOI222XL U52763 ( .A0(net265321), .A1(n50748), .B0(n40234), .B1(n50747),
        .C0(n40334), .C1(n50746), .Y(n17042) );
  AOI222XL U52764 ( .A0(net265321), .A1(n50747), .B0(n40234), .B1(n50746),
        .C0(n40334), .C1(n50745), .Y(n17018) );
  AOI222XL U52765 ( .A0(net265302), .A1(n50746), .B0(n40235), .B1(n50745),
        .C0(n40334), .C1(n50744), .Y(n16994) );
  AOI222XL U52766 ( .A0(net265302), .A1(n50745), .B0(n40235), .B1(n50744),
        .C0(n40335), .C1(n50743), .Y(n16970) );
  AOI222XL U52767 ( .A0(net264960), .A1(n50744), .B0(n40256), .B1(n50743),
        .C0(n40335), .C1(n50742), .Y(n16946) );
  AOI222XL U52768 ( .A0(net264960), .A1(n50743), .B0(n40256), .B1(n50742),
        .C0(n40335), .C1(n50741), .Y(n16922) );
  AOI222XL U52769 ( .A0(net264941), .A1(n50742), .B0(n40257), .B1(n50741),
        .C0(n40336), .C1(n50740), .Y(n16898) );
  AOI222XL U52770 ( .A0(net264941), .A1(n50741), .B0(n40257), .B1(n50740),
        .C0(n40336), .C1(n50739), .Y(n16874) );
  AOI222XL U52771 ( .A0(net264941), .A1(n50740), .B0(n40257), .B1(n50739),
        .C0(n40336), .C1(n50738), .Y(n16850) );
  AOI222XL U52772 ( .A0(net264922), .A1(n50739), .B0(n40258), .B1(n50738),
        .C0(n40337), .C1(n50737), .Y(n16826) );
  AOI222XL U52773 ( .A0(net264922), .A1(n50738), .B0(n40258), .B1(n50737),
        .C0(n40337), .C1(n50736), .Y(n16802) );
  AOI222XL U52774 ( .A0(net264922), .A1(n50737), .B0(n40259), .B1(n50736),
        .C0(n40337), .C1(n50735), .Y(n16778) );
  AOI222XL U52775 ( .A0(net264903), .A1(n50736), .B0(n40259), .B1(n50735),
        .C0(n40338), .C1(n50734), .Y(n16754) );
  AOI222XL U52776 ( .A0(net264903), .A1(n50735), .B0(n40259), .B1(n50734),
        .C0(n40338), .C1(n50733), .Y(n16730) );
  AOI222XL U52777 ( .A0(net265473), .A1(n50734), .B0(n40260), .B1(n50733),
        .C0(n40338), .C1(n50732), .Y(n16706) );
  AOI222XL U52778 ( .A0(net264884), .A1(n50733), .B0(n40260), .B1(n50732),
        .C0(n40339), .C1(n50731), .Y(n16682) );
  AOI222XL U52779 ( .A0(net264884), .A1(n50732), .B0(n40261), .B1(n50731),
        .C0(n40339), .C1(n50730), .Y(n16658) );
  AOI222XL U52780 ( .A0(net264884), .A1(n50731), .B0(n40261), .B1(n50730),
        .C0(n40340), .C1(n50729), .Y(n16634) );
  AOI222XL U52781 ( .A0(net265207), .A1(n50730), .B0(n40266), .B1(n50729),
        .C0(n40340), .C1(n50728), .Y(n16610) );
  AOI222XL U52782 ( .A0(net264808), .A1(n50729), .B0(n40266), .B1(n50728),
        .C0(n40340), .C1(n50727), .Y(n16586) );
  AOI222XL U52783 ( .A0(net264808), .A1(n50728), .B0(n40265), .B1(n50727),
        .C0(n40341), .C1(n50726), .Y(n16562) );
  AOI222XL U52784 ( .A0(net264808), .A1(n50727), .B0(n40265), .B1(n50726),
        .C0(n40341), .C1(n50725), .Y(n16538) );
  AOI222XL U52785 ( .A0(net264827), .A1(n50726), .B0(n40264), .B1(n50725),
        .C0(n40341), .C1(n50724), .Y(n16514) );
  AOI222XL U52786 ( .A0(net264827), .A1(n50725), .B0(n40264), .B1(n50724),
        .C0(n40342), .C1(n50723), .Y(n16490) );
  AOI222XL U52787 ( .A0(net264827), .A1(n50724), .B0(n40264), .B1(n50723),
        .C0(n40342), .C1(n50722), .Y(n16466) );
  AOI222XL U52788 ( .A0(net264846), .A1(n50723), .B0(n40263), .B1(n50722),
        .C0(n40342), .C1(n50721), .Y(n16442) );
  AOI222XL U52789 ( .A0(net264846), .A1(n50722), .B0(n40263), .B1(n50721),
        .C0(n40343), .C1(n50720), .Y(n16418) );
  AOI222XL U52790 ( .A0(net264846), .A1(n50721), .B0(n40262), .B1(n50720),
        .C0(n40343), .C1(n50719), .Y(n16394) );
  AOI222XL U52791 ( .A0(net264865), .A1(n50720), .B0(n40262), .B1(n50719),
        .C0(n40343), .C1(n50718), .Y(n16370) );
  AOI222XL U52792 ( .A0(net264865), .A1(n50719), .B0(n40262), .B1(n50718),
        .C0(n40344), .C1(n50717), .Y(n16346) );
  AOI222XL U52793 ( .A0(net264865), .A1(n50718), .B0(n40261), .B1(n50717),
        .C0(n40344), .C1(n50716), .Y(n16322) );
  AOI222XL U52794 ( .A0(net265131), .A1(n50717), .B0(n40245), .B1(n50716),
        .C0(n40344), .C1(n50715), .Y(n16298) );
  AOI222XL U52795 ( .A0(net265112), .A1(n50716), .B0(n40246), .B1(n50715),
        .C0(n40345), .C1(n50714), .Y(n16274) );
  AOI222XL U52796 ( .A0(net265112), .A1(n50715), .B0(n40246), .B1(n50714),
        .C0(n40345), .C1(n50713), .Y(n16250) );
  AOI222XL U52797 ( .A0(net265112), .A1(n50714), .B0(n40247), .B1(n50713),
        .C0(n40346), .C1(n50712), .Y(n16226) );
  AOI222XL U52798 ( .A0(net221810), .A1(n50713), .B0(n40247), .B1(n50712),
        .C0(n40346), .C1(n50711), .Y(n16202) );
  AOI222XL U52799 ( .A0(net221814), .A1(n50712), .B0(n40247), .B1(n50711),
        .C0(n40346), .C1(n50710), .Y(n16178) );
  AOI222XL U52800 ( .A0(net221802), .A1(n50711), .B0(n40248), .B1(n50710),
        .C0(n40347), .C1(n50709), .Y(n16154) );
  AOI222XL U52801 ( .A0(net265074), .A1(n50710), .B0(n40248), .B1(n50709),
        .C0(n40347), .C1(n50708), .Y(n16130) );
  AOI222XL U52802 ( .A0(net265074), .A1(n50709), .B0(n40249), .B1(n50708),
        .C0(n40347), .C1(n50707), .Y(n16106) );
  AOI222XL U52803 ( .A0(net265074), .A1(n50708), .B0(n40249), .B1(n50707),
        .C0(n40348), .C1(n50706), .Y(n16082) );
  AOI222XL U52804 ( .A0(net265055), .A1(n50707), .B0(n40249), .B1(n50706),
        .C0(n40348), .C1(n50705), .Y(n16058) );
  AOI222XL U52805 ( .A0(net265055), .A1(n50706), .B0(n40250), .B1(n50705),
        .C0(n40348), .C1(n50704), .Y(n16034) );
  AOI222XL U52806 ( .A0(net265055), .A1(n50705), .B0(n40250), .B1(n50704),
        .C0(n40349), .C1(n50703), .Y(n16010) );
  AOI222XL U52807 ( .A0(net265036), .A1(n50704), .B0(n40251), .B1(n50703),
        .C0(n40349), .C1(n50702), .Y(n15986) );
  AOI222XL U52808 ( .A0(net265036), .A1(n50703), .B0(n40251), .B1(n50702),
        .C0(n40349), .C1(n50701), .Y(n15962) );
  AOI222XL U52809 ( .A0(net265036), .A1(n50702), .B0(n40251), .B1(n50701),
        .C0(n40383), .C1(n50700), .Y(n15938) );
  AOI222XL U52810 ( .A0(net265017), .A1(n50701), .B0(n40252), .B1(n50700),
        .C0(n40383), .C1(n50699), .Y(n15914) );
  AOI222XL U52811 ( .A0(net265017), .A1(n50700), .B0(n40252), .B1(n50699),
        .C0(n40382), .C1(n50698), .Y(n15890) );
  AOI222XL U52812 ( .A0(net265017), .A1(n50699), .B0(n40253), .B1(n50698),
        .C0(n40350), .C1(n50697), .Y(n15866) );
  AOI222XL U52813 ( .A0(net264998), .A1(n50698), .B0(n40253), .B1(n50697),
        .C0(n40350), .C1(n50696), .Y(n15842) );
  AOI222XL U52814 ( .A0(net264998), .A1(n50697), .B0(n40253), .B1(n50696),
        .C0(n40341), .C1(n50695), .Y(n15818) );
  AOI222XL U52815 ( .A0(net264998), .A1(n50696), .B0(n40254), .B1(n50695),
        .C0(net217036), .C1(n50694), .Y(n15794) );
  AOI222XL U52816 ( .A0(net264979), .A1(n50695), .B0(n40254), .B1(n50694),
        .C0(net217036), .C1(n50693), .Y(n15770) );
  AOI222XL U52817 ( .A0(net264979), .A1(n50694), .B0(n40255), .B1(n50693),
        .C0(n40351), .C1(n50692), .Y(n15746) );
  AOI222XL U52818 ( .A0(net264979), .A1(n50693), .B0(n40255), .B1(n50692),
        .C0(n40351), .C1(n50691), .Y(n15722) );
  AOI222XL U52819 ( .A0(net264960), .A1(n50692), .B0(n40255), .B1(n50691),
        .C0(n40351), .C1(n50690), .Y(n15698) );
  AOI222XL U52820 ( .A0(net265055), .A1(n50691), .B0(n40245), .B1(n50690),
        .C0(n40352), .C1(n50689), .Y(n15674) );
  AOI222XL U52821 ( .A0(net265967), .A1(n50690), .B0(n40193), .B1(n50689),
        .C0(n40352), .C1(n50688), .Y(n15650) );
  AOI222XL U52822 ( .A0(net265967), .A1(n50689), .B0(n40193), .B1(n50688),
        .C0(n40352), .C1(n50687), .Y(n15626) );
  AOI222XL U52823 ( .A0(net265967), .A1(n50688), .B0(n40194), .B1(n50687),
        .C0(n40353), .C1(n50686), .Y(n15602) );
  AOI222XL U52824 ( .A0(net265948), .A1(n50687), .B0(n40194), .B1(n50686),
        .C0(n40353), .C1(n50685), .Y(n15578) );
  AOI222XL U52825 ( .A0(net265948), .A1(n50686), .B0(n40195), .B1(n50685),
        .C0(n40353), .C1(n50684), .Y(n15554) );
  AOI222XL U52826 ( .A0(net265948), .A1(n50685), .B0(n40195), .B1(n50684),
        .C0(n40354), .C1(n50683), .Y(n15530) );
  AOI222XL U52827 ( .A0(net265929), .A1(n50684), .B0(n40195), .B1(n50683),
        .C0(n40354), .C1(n50682), .Y(n15506) );
  AOI222XL U52828 ( .A0(net265929), .A1(n50683), .B0(n40196), .B1(n50682),
        .C0(n40354), .C1(n50681), .Y(n15482) );
  AOI222XL U52829 ( .A0(net265929), .A1(n50682), .B0(n40196), .B1(n50681),
        .C0(n40355), .C1(n50680), .Y(n15458) );
  AOI222XL U52830 ( .A0(net265910), .A1(n50681), .B0(n40197), .B1(n50680),
        .C0(n40355), .C1(n50679), .Y(n15434) );
  AOI222XL U52831 ( .A0(net265910), .A1(n50680), .B0(n40197), .B1(n50679),
        .C0(n40356), .C1(n50678), .Y(n15410) );
  AOI222XL U52832 ( .A0(net265910), .A1(n50679), .B0(n40197), .B1(n50678),
        .C0(n40356), .C1(n50677), .Y(n15386) );
  AOI222XL U52833 ( .A0(net265891), .A1(n50678), .B0(n40198), .B1(n50677),
        .C0(n40356), .C1(n50676), .Y(n15362) );
  AOI222XL U52834 ( .A0(net265891), .A1(n50677), .B0(n40198), .B1(n50676),
        .C0(n40357), .C1(n50675), .Y(n15338) );
  AOI222XL U52835 ( .A0(net265891), .A1(n50676), .B0(n40199), .B1(n50675),
        .C0(n40357), .C1(n50674), .Y(n15314) );
  AOI222XL U52836 ( .A0(net265872), .A1(n50675), .B0(n40199), .B1(n50674),
        .C0(n40357), .C1(n50673), .Y(n15290) );
  AOI222XL U52837 ( .A0(net265872), .A1(n50674), .B0(n40200), .B1(n50673),
        .C0(n40358), .C1(n50672), .Y(n15266) );
  AOI222XL U52838 ( .A0(net265872), .A1(n50673), .B0(n40200), .B1(n50672),
        .C0(n40358), .C1(n50671), .Y(n15242) );
  AOI222XL U52839 ( .A0(net265853), .A1(n50672), .B0(n40200), .B1(n50671),
        .C0(n40358), .C1(n50670), .Y(n15218) );
  AOI222XL U52840 ( .A0(net265853), .A1(n50671), .B0(n40201), .B1(n50670),
        .C0(n40359), .C1(n50669), .Y(n15194) );
  AOI222XL U52841 ( .A0(net265853), .A1(n50670), .B0(n40201), .B1(n50669),
        .C0(n40359), .C1(n50668), .Y(n15170) );
  AOI222XL U52842 ( .A0(net265834), .A1(n50669), .B0(n40202), .B1(n50668),
        .C0(n40359), .C1(n50667), .Y(n15146) );
  AOI222XL U52843 ( .A0(net265834), .A1(n50668), .B0(n40202), .B1(n50667),
        .C0(n40360), .C1(n50666), .Y(n15122) );
  AOI222XL U52844 ( .A0(net265834), .A1(n50667), .B0(n40202), .B1(n50666),
        .C0(n40360), .C1(n50665), .Y(n15098) );
  AOI222XL U52845 ( .A0(net265815), .A1(n50666), .B0(n40203), .B1(n50665),
        .C0(n40360), .C1(n50664), .Y(n15074) );
  AOI222XL U52846 ( .A0(net265815), .A1(n50665), .B0(n40203), .B1(n50664),
        .C0(n40377), .C1(n50663), .Y(n15050) );
  AOI222XL U52847 ( .A0(net221892), .A1(n50663), .B0(n40184), .B1(n50662),
        .C0(n40361), .C1(n50661), .Y(n15002) );
  AOI222XL U52848 ( .A0(net221892), .A1(n50662), .B0(n40184), .B1(n50661),
        .C0(n40361), .C1(n50660), .Y(n14978) );
  AOI222XL U52849 ( .A0(net266119), .A1(n50661), .B0(n40184), .B1(n50660),
        .C0(n40361), .C1(n50659), .Y(n14954) );
  AOI222XL U52850 ( .A0(net266119), .A1(n50660), .B0(n40185), .B1(n50659),
        .C0(n40362), .C1(n50658), .Y(n14930) );
  OAI211X1 U52851 ( .A0(n32992), .A1(n42985), .B0(n14905), .C0(n14906), .Y(
        n35141) );
  OA22X1 U52852 ( .A0(net263748), .A1(n32976), .B0(n32984), .B1(n40053), .Y(
        n14905) );
  AOI222XL U52853 ( .A0(net266119), .A1(n50659), .B0(n40185), .B1(n50658),
        .C0(n40362), .C1(n50657), .Y(n14906) );
  OAI211X1 U52854 ( .A0(n32984), .A1(n42986), .B0(n14881), .C0(n14882), .Y(
        n35133) );
  AOI222XL U52855 ( .A0(net266100), .A1(n50658), .B0(n40197), .B1(n50657),
        .C0(n40362), .C1(n50656), .Y(n14882) );
  OAI211X1 U52856 ( .A0(n32976), .A1(n42987), .B0(n14857), .C0(n14858), .Y(
        n35125) );
  OA22X1 U52857 ( .A0(net263767), .A1(n32960), .B0(n32968), .B1(n40052), .Y(
        n14857) );
  AOI222XL U52858 ( .A0(net266100), .A1(n50657), .B0(n40195), .B1(n50656),
        .C0(n40363), .C1(n50655), .Y(n14858) );
  OAI211X1 U52859 ( .A0(n32968), .A1(n42989), .B0(n14833), .C0(n14834), .Y(
        n35117) );
  OA22X1 U52860 ( .A0(net263539), .A1(n32952), .B0(n32960), .B1(n40052), .Y(
        n14833) );
  AOI222XL U52861 ( .A0(net266100), .A1(n50656), .B0(n40194), .B1(n50655),
        .C0(n40363), .C1(n50654), .Y(n14834) );
  OAI211X1 U52862 ( .A0(n32960), .A1(n42990), .B0(n14809), .C0(n14810), .Y(
        n35109) );
  OA22X1 U52863 ( .A0(net263026), .A1(n32944), .B0(n32952), .B1(n40051), .Y(
        n14809) );
  AOI222XL U52864 ( .A0(net266081), .A1(n50655), .B0(n40186), .B1(n50654),
        .C0(n40363), .C1(n50653), .Y(n14810) );
  OAI211X1 U52865 ( .A0(n32952), .A1(n42975), .B0(n14785), .C0(n14786), .Y(
        n35101) );
  OA22X1 U52866 ( .A0(net263805), .A1(n32936), .B0(n32944), .B1(n40051), .Y(
        n14785) );
  AOI222XL U52867 ( .A0(net266081), .A1(n50654), .B0(n40186), .B1(n50653),
        .C0(n40364), .C1(n50652), .Y(n14786) );
  OAI211X1 U52868 ( .A0(n32944), .A1(n42968), .B0(n14761), .C0(n14762), .Y(
        n35093) );
  OA22X1 U52869 ( .A0(net263805), .A1(n32928), .B0(n32936), .B1(n40050), .Y(
        n14761) );
  AOI222XL U52870 ( .A0(net266081), .A1(n50653), .B0(n40187), .B1(n50652),
        .C0(n40374), .C1(n50651), .Y(n14762) );
  OAI211X1 U52871 ( .A0(n32936), .A1(n42961), .B0(n14737), .C0(n14738), .Y(
        n35085) );
  OA22X1 U52872 ( .A0(net263805), .A1(n32920), .B0(n32928), .B1(n40050), .Y(
        n14737) );
  AOI222XL U52873 ( .A0(net266062), .A1(n50652), .B0(n40187), .B1(n50651),
        .C0(n40374), .C1(n50650), .Y(n14738) );
  OAI211X1 U52874 ( .A0(n32928), .A1(n42962), .B0(n14713), .C0(n14714), .Y(
        n35077) );
  OA22X1 U52875 ( .A0(net263824), .A1(n32912), .B0(n32920), .B1(n40049), .Y(
        n14713) );
  AOI222XL U52876 ( .A0(net266062), .A1(n50651), .B0(n40187), .B1(n50650),
        .C0(n40364), .C1(n50649), .Y(n14714) );
  OAI211X1 U52877 ( .A0(n32920), .A1(n42963), .B0(n14689), .C0(n14690), .Y(
        n35069) );
  OA22X1 U52878 ( .A0(net263824), .A1(n32904), .B0(n32912), .B1(n40049), .Y(
        n14689) );
  AOI222XL U52879 ( .A0(net266062), .A1(n50650), .B0(n40188), .B1(n50649),
        .C0(n40364), .C1(n50648), .Y(n14690) );
  OAI211X1 U52880 ( .A0(n32912), .A1(n42964), .B0(n14665), .C0(n14666), .Y(
        n35061) );
  OA22X1 U52881 ( .A0(net263843), .A1(n32896), .B0(n32904), .B1(n40048), .Y(
        n14665) );
  AOI222XL U52882 ( .A0(net266043), .A1(n50649), .B0(n40188), .B1(n50648),
        .C0(n40364), .C1(n50647), .Y(n14666) );
  OAI211X1 U52883 ( .A0(n32904), .A1(n42965), .B0(n14641), .C0(n14642), .Y(
        n35053) );
  OA22X1 U52884 ( .A0(net263843), .A1(n32888), .B0(n32896), .B1(n40048), .Y(
        n14641) );
  AOI222XL U52885 ( .A0(net266043), .A1(n50648), .B0(n40189), .B1(n50647),
        .C0(n40365), .C1(n50646), .Y(n14642) );
  OAI211X1 U52886 ( .A0(n32896), .A1(n42967), .B0(n14617), .C0(n14618), .Y(
        n35045) );
  OA22X1 U52887 ( .A0(net263862), .A1(n32880), .B0(n32888), .B1(n40047), .Y(
        n14617) );
  AOI222XL U52888 ( .A0(net266043), .A1(n50647), .B0(n40189), .B1(n50646),
        .C0(n40365), .C1(n50645), .Y(n14618) );
  OAI211X1 U52889 ( .A0(n32888), .A1(n42968), .B0(n14593), .C0(n14594), .Y(
        n35037) );
  OA22X1 U52890 ( .A0(net263862), .A1(n32872), .B0(n32880), .B1(n40047), .Y(
        n14593) );
  AOI222XL U52891 ( .A0(net266024), .A1(n50646), .B0(n40189), .B1(n50645),
        .C0(n40366), .C1(n50644), .Y(n14594) );
  OAI211X1 U52892 ( .A0(n32880), .A1(n42969), .B0(n14569), .C0(n14570), .Y(
        n35029) );
  OA22X1 U52893 ( .A0(net263121), .A1(n32864), .B0(n32872), .B1(n40088), .Y(
        n14569) );
  AOI222XL U52894 ( .A0(net266024), .A1(n50645), .B0(n40190), .B1(n50644),
        .C0(n40366), .C1(n50643), .Y(n14570) );
  OAI211X1 U52895 ( .A0(n32872), .A1(n42970), .B0(n14545), .C0(n14546), .Y(
        n35021) );
  OA22X1 U52896 ( .A0(net263064), .A1(n32856), .B0(n32864), .B1(n40092), .Y(
        n14545) );
  AOI222XL U52897 ( .A0(net266024), .A1(n50644), .B0(n40190), .B1(n50643),
        .C0(n40366), .C1(n50642), .Y(n14546) );
  OAI211X1 U52898 ( .A0(n32864), .A1(n42971), .B0(n14521), .C0(n14522), .Y(
        n35013) );
  OA22X1 U52899 ( .A0(net263083), .A1(n32848), .B0(n32856), .B1(n40091), .Y(
        n14521) );
  AOI222XL U52900 ( .A0(net266005), .A1(n50643), .B0(n40191), .B1(n50642),
        .C0(n40367), .C1(n50641), .Y(n14522) );
  OAI211X1 U52901 ( .A0(n32856), .A1(n42972), .B0(n14497), .C0(n14498), .Y(
        n35005) );
  OA22X1 U52902 ( .A0(net263083), .A1(n32840), .B0(n32848), .B1(n40091), .Y(
        n14497) );
  AOI222XL U52903 ( .A0(net266005), .A1(n50642), .B0(n40191), .B1(n50641),
        .C0(n40367), .C1(n50640), .Y(n14498) );
  OAI211X1 U52904 ( .A0(n32848), .A1(n42974), .B0(n14473), .C0(n14474), .Y(
        n34997) );
  OA22X1 U52905 ( .A0(net263102), .A1(n32832), .B0(n32840), .B1(n40090), .Y(
        n14473) );
  AOI222XL U52906 ( .A0(net266005), .A1(n50641), .B0(n40191), .B1(n50640),
        .C0(n40367), .C1(n50639), .Y(n14474) );
  OAI211X1 U52907 ( .A0(n32840), .A1(n42975), .B0(n14449), .C0(n14450), .Y(
        n34989) );
  OA22X1 U52908 ( .A0(net263102), .A1(n32824), .B0(n32832), .B1(n40090), .Y(
        n14449) );
  AOI222XL U52909 ( .A0(net265796), .A1(n50640), .B0(n40192), .B1(n50639),
        .C0(n40368), .C1(n50638), .Y(n14450) );
  OAI211X1 U52910 ( .A0(n32832), .A1(n42976), .B0(n14425), .C0(n14426), .Y(
        n34981) );
  OA22X1 U52911 ( .A0(net263102), .A1(n32816), .B0(n32824), .B1(n40089), .Y(
        n14425) );
  AOI222XL U52912 ( .A0(net265777), .A1(n50639), .B0(n40192), .B1(n50638),
        .C0(n40368), .C1(n50637), .Y(n14426) );
  OAI211X1 U52913 ( .A0(n32824), .A1(n42880), .B0(n14401), .C0(n14402), .Y(
        n34973) );
  OA22X1 U52914 ( .A0(net263121), .A1(n32808), .B0(n32816), .B1(n40089), .Y(
        n14401) );
  AOI222XL U52915 ( .A0(net265739), .A1(n50638), .B0(n40193), .B1(n50637),
        .C0(n40368), .C1(n50636), .Y(n14402) );
  OAI211X1 U52916 ( .A0(n32816), .A1(n42881), .B0(n14377), .C0(n14378), .Y(
        n34965) );
  OA22X1 U52917 ( .A0(net263121), .A1(n32800), .B0(n32808), .B1(n40088), .Y(
        n14377) );
  AOI222XL U52918 ( .A0(net265644), .A1(n50637), .B0(n40214), .B1(n50636),
        .C0(n40369), .C1(n50635), .Y(n14378) );
  OAI211X1 U52919 ( .A0(n32808), .A1(n42882), .B0(n14353), .C0(n14354), .Y(
        n34957) );
  OA22X1 U52920 ( .A0(net263140), .A1(n32792), .B0(n32800), .B1(n40088), .Y(
        n14353) );
  AOI222XL U52921 ( .A0(net265625), .A1(n50636), .B0(n40215), .B1(n50635),
        .C0(n40369), .C1(n50634), .Y(n14354) );
  OAI211X1 U52922 ( .A0(n32800), .A1(n42883), .B0(n14329), .C0(n14330), .Y(
        n34949) );
  OA22X1 U52923 ( .A0(net263140), .A1(n32784), .B0(n32792), .B1(n40087), .Y(
        n14329) );
  AOI222XL U52924 ( .A0(net265625), .A1(n50635), .B0(n40215), .B1(n50634),
        .C0(n40369), .C1(n50633), .Y(n14330) );
  OAI211X1 U52925 ( .A0(n32792), .A1(n42884), .B0(n14305), .C0(n14306), .Y(
        n34941) );
  OA22X1 U52926 ( .A0(net263159), .A1(n32776), .B0(n32784), .B1(n40087), .Y(
        n14305) );
  AOI222XL U52927 ( .A0(net265625), .A1(n50634), .B0(n40215), .B1(n50633),
        .C0(n40370), .C1(n50632), .Y(n14306) );
  OAI211X1 U52928 ( .A0(n32784), .A1(n42886), .B0(n14281), .C0(n14282), .Y(
        n34933) );
  OA22X1 U52929 ( .A0(net263159), .A1(n32768), .B0(n32776), .B1(n40086), .Y(
        n14281) );
  AOI222XL U52930 ( .A0(net265606), .A1(n50633), .B0(n40216), .B1(n50632),
        .C0(n40370), .C1(n50631), .Y(n14282) );
  OAI211X1 U52931 ( .A0(n32776), .A1(n42887), .B0(n14257), .C0(n14258), .Y(
        n34925) );
  OA22X1 U52932 ( .A0(net263178), .A1(n32760), .B0(n32768), .B1(n40086), .Y(
        n14257) );
  AOI222XL U52933 ( .A0(net265606), .A1(n50632), .B0(n40216), .B1(n50631),
        .C0(n40370), .C1(n50630), .Y(n14258) );
  OAI211X1 U52934 ( .A0(n32768), .A1(n42888), .B0(n14233), .C0(n14234), .Y(
        n34917) );
  OA22X1 U52935 ( .A0(net263178), .A1(n32752), .B0(n32760), .B1(n40085), .Y(
        n14233) );
  AOI222XL U52936 ( .A0(net265606), .A1(n50631), .B0(n40217), .B1(n50630),
        .C0(n40371), .C1(n50629), .Y(n14234) );
  OAI211X1 U52937 ( .A0(n32760), .A1(n42889), .B0(n14209), .C0(n14210), .Y(
        n34909) );
  OA22X1 U52938 ( .A0(net218352), .A1(n32744), .B0(n32752), .B1(n40085), .Y(
        n14209) );
  AOI222XL U52939 ( .A0(net265587), .A1(n50630), .B0(n40217), .B1(n50629),
        .C0(n40371), .C1(n50628), .Y(n14210) );
  OAI211X1 U52940 ( .A0(n32752), .A1(n42890), .B0(n14185), .C0(n14186), .Y(
        n34901) );
  OA22X1 U52941 ( .A0(net262931), .A1(n32736), .B0(n32744), .B1(n40100), .Y(
        n14185) );
  AOI222XL U52942 ( .A0(net265587), .A1(n50629), .B0(n40217), .B1(n50628),
        .C0(n40372), .C1(n50627), .Y(n14186) );
  OAI211X1 U52943 ( .A0(n32744), .A1(n42891), .B0(n14161), .C0(n14162), .Y(
        n34893) );
  OA22X1 U52944 ( .A0(net262931), .A1(n32728), .B0(n32736), .B1(n40100), .Y(
        n14161) );
  AOI222XL U52945 ( .A0(net265587), .A1(n50628), .B0(n40218), .B1(n50627),
        .C0(n40372), .C1(n50626), .Y(n14162) );
  OAI211X1 U52946 ( .A0(n32736), .A1(n42893), .B0(n14137), .C0(n14138), .Y(
        n34885) );
  OA22X1 U52947 ( .A0(net262950), .A1(n32720), .B0(n32728), .B1(n40099), .Y(
        n14137) );
  AOI222XL U52948 ( .A0(net265568), .A1(n50627), .B0(n40218), .B1(n50626),
        .C0(n40372), .C1(n50625), .Y(n14138) );
  OAI211X1 U52949 ( .A0(n32728), .A1(n42894), .B0(n14113), .C0(n14114), .Y(
        n34877) );
  OA22X1 U52950 ( .A0(net262950), .A1(n32712), .B0(n32720), .B1(n40099), .Y(
        n14113) );
  AOI222XL U52951 ( .A0(net265568), .A1(n50626), .B0(n40219), .B1(n50625),
        .C0(n40373), .C1(n50624), .Y(n14114) );
  OAI211X1 U52952 ( .A0(n32720), .A1(n42895), .B0(n14089), .C0(n14090), .Y(
        n34869) );
  OA22X1 U52953 ( .A0(net262969), .A1(n32704), .B0(n32712), .B1(n40098), .Y(
        n14089) );
  AOI222XL U52954 ( .A0(net265568), .A1(n50625), .B0(n40219), .B1(n50624),
        .C0(n40373), .C1(n50623), .Y(n14090) );
  OAI211X1 U52955 ( .A0(n32712), .A1(n42864), .B0(n14065), .C0(n14066), .Y(
        n34861) );
  OA22X1 U52956 ( .A0(net262969), .A1(n32696), .B0(n32704), .B1(n40098), .Y(
        n14065) );
  AOI222XL U52957 ( .A0(net265549), .A1(n50624), .B0(n40220), .B1(n50623),
        .C0(n40373), .C1(n50622), .Y(n14066) );
  OAI211X1 U52958 ( .A0(n32704), .A1(n42865), .B0(n14041), .C0(n14042), .Y(
        n34853) );
  OA22X1 U52959 ( .A0(net262969), .A1(n32688), .B0(n32696), .B1(n40097), .Y(
        n14041) );
  AOI222XL U52960 ( .A0(net265549), .A1(n50623), .B0(n40220), .B1(n50622),
        .C0(n40374), .C1(n50621), .Y(n14042) );
  OAI211X1 U52961 ( .A0(n32696), .A1(n42866), .B0(n14017), .C0(n14018), .Y(
        n34845) );
  OA22X1 U52962 ( .A0(net262988), .A1(n32680), .B0(n32688), .B1(n40097), .Y(
        n14017) );
  AOI222XL U52963 ( .A0(net265549), .A1(n50622), .B0(n40220), .B1(n50621),
        .C0(n40374), .C1(n50620), .Y(n14018) );
  OAI211X1 U52964 ( .A0(n32688), .A1(n42867), .B0(n13993), .C0(n13994), .Y(
        n34837) );
  OA22X1 U52965 ( .A0(net262988), .A1(n32672), .B0(n32680), .B1(n40096), .Y(
        n13993) );
  AOI222XL U52966 ( .A0(net265530), .A1(n50621), .B0(n40221), .B1(n50620),
        .C0(n40374), .C1(n50619), .Y(n13994) );
  OAI211X1 U52967 ( .A0(n32680), .A1(n42868), .B0(n13969), .C0(n13970), .Y(
        n34829) );
  OA22X1 U52968 ( .A0(net263007), .A1(n32664), .B0(n32672), .B1(n40096), .Y(
        n13969) );
  AOI222XL U52969 ( .A0(net265530), .A1(n50620), .B0(n40221), .B1(n50619),
        .C0(n40375), .C1(n50618), .Y(n13970) );
  OAI211X1 U52970 ( .A0(n32672), .A1(n42870), .B0(n13945), .C0(n13946), .Y(
        n34821) );
  OA22X1 U52971 ( .A0(net263007), .A1(n32656), .B0(n32664), .B1(n40095), .Y(
        n13945) );
  AOI222XL U52972 ( .A0(net265530), .A1(n50619), .B0(n40222), .B1(n50618),
        .C0(n40375), .C1(n50617), .Y(n13946) );
  OAI211X1 U52973 ( .A0(n32664), .A1(n42871), .B0(n13921), .C0(n13922), .Y(
        n34813) );
  OA22X1 U52974 ( .A0(net263026), .A1(n32648), .B0(n32656), .B1(n40095), .Y(
        n13921) );
  AOI222XL U52975 ( .A0(net265511), .A1(n50618), .B0(n40222), .B1(n50617),
        .C0(n40375), .C1(n50616), .Y(n13922) );
  OAI211X1 U52976 ( .A0(n32656), .A1(n42872), .B0(n13897), .C0(n13898), .Y(
        n34805) );
  OA22X1 U52977 ( .A0(net263026), .A1(n32640), .B0(n32648), .B1(n40094), .Y(
        n13897) );
  AOI222XL U52978 ( .A0(net265511), .A1(n50617), .B0(n40222), .B1(n50616),
        .C0(n40376), .C1(n50615), .Y(n13898) );
  OAI211X1 U52979 ( .A0(n32648), .A1(n42873), .B0(n13873), .C0(n13874), .Y(
        n34797) );
  OA22X1 U52980 ( .A0(net263045), .A1(n32632), .B0(n32640), .B1(n40094), .Y(
        n13873) );
  AOI222XL U52981 ( .A0(net265511), .A1(n50616), .B0(n40223), .B1(n50615),
        .C0(n40376), .C1(n50614), .Y(n13874) );
  OAI211X1 U52982 ( .A0(n32640), .A1(n42874), .B0(n13849), .C0(n13850), .Y(
        n34789) );
  OA22X1 U52983 ( .A0(net263045), .A1(n32624), .B0(n32632), .B1(n40093), .Y(
        n13849) );
  AOI222XL U52984 ( .A0(net265492), .A1(n50615), .B0(n40223), .B1(n50614),
        .C0(n40376), .C1(n50613), .Y(n13850) );
  OAI211X1 U52985 ( .A0(n32632), .A1(n42875), .B0(n13825), .C0(n13826), .Y(
        n34781) );
  OA22X1 U52986 ( .A0(net263045), .A1(n32616), .B0(n32624), .B1(n40093), .Y(
        n13825) );
  AOI222XL U52987 ( .A0(net265492), .A1(n50614), .B0(n40224), .B1(n50613),
        .C0(n40377), .C1(n50612), .Y(n13826) );
  OAI211X1 U52988 ( .A0(n32624), .A1(n42877), .B0(n13801), .C0(n13802), .Y(
        n34773) );
  OA22X1 U52989 ( .A0(net263330), .A1(n32608), .B0(n32616), .B1(n40077), .Y(
        n13801) );
  AOI222XL U52990 ( .A0(net265492), .A1(n50613), .B0(n40224), .B1(n50612),
        .C0(n40377), .C1(n50611), .Y(n13802) );
  OAI211X1 U52991 ( .A0(n32616), .A1(n42878), .B0(n13777), .C0(n13778), .Y(
        n34765) );
  OA22X1 U52992 ( .A0(net263349), .A1(n32600), .B0(n32608), .B1(n40077), .Y(
        n13777) );
  AOI222XL U52993 ( .A0(net265473), .A1(n50612), .B0(n40224), .B1(n50611),
        .C0(n40378), .C1(n50610), .Y(n13778) );
  OAI211X1 U52994 ( .A0(n32608), .A1(n42879), .B0(n13753), .C0(n13754), .Y(
        n34757) );
  OA22X1 U52995 ( .A0(net263349), .A1(n32592), .B0(n32600), .B1(n40076), .Y(
        n13753) );
  AOI222XL U52996 ( .A0(net265473), .A1(n50611), .B0(n40219), .B1(n50610),
        .C0(n40378), .C1(n50609), .Y(n13754) );
  OAI211X1 U52997 ( .A0(n32600), .A1(n42912), .B0(n13729), .C0(n13730), .Y(
        n34749) );
  OA22X1 U52998 ( .A0(net263349), .A1(n32584), .B0(n32592), .B1(n40076), .Y(
        n13729) );
  AOI222XL U52999 ( .A0(net265796), .A1(n50610), .B0(n40204), .B1(n50609),
        .C0(n40378), .C1(n50608), .Y(n13730) );
  OAI211X1 U53000 ( .A0(n32592), .A1(n42913), .B0(n13705), .C0(n13706), .Y(
        n34741) );
  OA22X1 U53001 ( .A0(net263368), .A1(n32576), .B0(n32584), .B1(n40075), .Y(
        n13705) );
  AOI222XL U53002 ( .A0(net265796), .A1(n50609), .B0(n40204), .B1(n50608),
        .C0(n40379), .C1(n50607), .Y(n13706) );
  OAI211X1 U53003 ( .A0(n32584), .A1(n42914), .B0(n13681), .C0(n13682), .Y(
        n34733) );
  OA22X1 U53004 ( .A0(net263368), .A1(n32568), .B0(n32576), .B1(n40075), .Y(
        n13681) );
  AOI222XL U53005 ( .A0(net265796), .A1(n50608), .B0(n40205), .B1(n50607),
        .C0(n40379), .C1(n50606), .Y(n13682) );
  OAI211X1 U53006 ( .A0(n32576), .A1(n42915), .B0(n13657), .C0(n13658), .Y(
        n34725) );
  OA22X1 U53007 ( .A0(net263387), .A1(n32560), .B0(n32568), .B1(n40074), .Y(
        n13657) );
  AOI222XL U53008 ( .A0(net265777), .A1(n50607), .B0(n40205), .B1(n50606),
        .C0(n40379), .C1(n50605), .Y(n13658) );
  OAI211X1 U53009 ( .A0(n32568), .A1(n42917), .B0(n13633), .C0(n13634), .Y(
        n34717) );
  OA22X1 U53010 ( .A0(net263387), .A1(n32552), .B0(n32560), .B1(n40074), .Y(
        n13633) );
  AOI222XL U53011 ( .A0(net265777), .A1(n50606), .B0(n40205), .B1(n50605),
        .C0(n40380), .C1(n50604), .Y(n13634) );
  OAI211X1 U53012 ( .A0(n32560), .A1(n42918), .B0(n13609), .C0(n13610), .Y(
        n34709) );
  OA22X1 U53013 ( .A0(net263406), .A1(n32544), .B0(n32552), .B1(n40073), .Y(
        n13609) );
  AOI222XL U53014 ( .A0(net265777), .A1(n50605), .B0(n40206), .B1(n50604),
        .C0(n40380), .C1(n50603), .Y(n13610) );
  OAI211X1 U53015 ( .A0(n32552), .A1(n42919), .B0(n13585), .C0(n13586), .Y(
        n34701) );
  OA22X1 U53016 ( .A0(net263406), .A1(n32536), .B0(n32544), .B1(n40073), .Y(
        n13585) );
  AOI222XL U53017 ( .A0(net265758), .A1(n50604), .B0(n40206), .B1(n50603),
        .C0(n40380), .C1(n50602), .Y(n13586) );
  OAI211X1 U53018 ( .A0(n32544), .A1(n42920), .B0(n13561), .C0(n13562), .Y(
        n34693) );
  OA22X1 U53019 ( .A0(net218408), .A1(n32528), .B0(n32536), .B1(n40072), .Y(
        n13561) );
  AOI222XL U53020 ( .A0(net265758), .A1(n50603), .B0(n40207), .B1(n50602),
        .C0(n40381), .C1(n50601), .Y(n13562) );
  OAI211X1 U53021 ( .A0(n32536), .A1(n42921), .B0(n13537), .C0(n13538), .Y(
        n34685) );
  OA22X1 U53022 ( .A0(net218334), .A1(n32520), .B0(n32528), .B1(n40072), .Y(
        n13537) );
  AOI222XL U53023 ( .A0(net265758), .A1(n50602), .B0(n40207), .B1(n50601),
        .C0(n40381), .C1(n50600), .Y(n13538) );
  OAI211X1 U53024 ( .A0(n32528), .A1(n42922), .B0(n13513), .C0(n13514), .Y(
        n34677) );
  OA22X1 U53025 ( .A0(net218418), .A1(n32512), .B0(n32520), .B1(n40071), .Y(
        n13513) );
  AOI222XL U53026 ( .A0(net265739), .A1(n50601), .B0(n40207), .B1(n50600),
        .C0(n40381), .C1(n50599), .Y(n13514) );
  OAI211X1 U53027 ( .A0(n32520), .A1(n42924), .B0(n13489), .C0(n13490), .Y(
        n34669) );
  OA22X1 U53028 ( .A0(net263444), .A1(n32504), .B0(n32512), .B1(n40071), .Y(
        n13489) );
  AOI222XL U53029 ( .A0(net265739), .A1(n50600), .B0(n40208), .B1(n50599),
        .C0(n40382), .C1(n50598), .Y(n13490) );
  OAI211X1 U53030 ( .A0(n32512), .A1(n42925), .B0(n13465), .C0(n13466), .Y(
        n34661) );
  OA22X1 U53031 ( .A0(net263444), .A1(n32496), .B0(n32504), .B1(n40070), .Y(
        n13465) );
  AOI222XL U53032 ( .A0(net265739), .A1(n50599), .B0(n40208), .B1(n50598),
        .C0(n40382), .C1(n50597), .Y(n13466) );
  OAI211X1 U53033 ( .A0(n32504), .A1(n42926), .B0(n13441), .C0(n13442), .Y(
        n34653) );
  OA22X1 U53034 ( .A0(net263463), .A1(n32488), .B0(n32496), .B1(n40070), .Y(
        n13441) );
  AOI222XL U53035 ( .A0(net265720), .A1(n50598), .B0(n40209), .B1(n50597),
        .C0(n40382), .C1(n50596), .Y(n13442) );
  OAI211X1 U53036 ( .A0(n32496), .A1(n42927), .B0(n13417), .C0(n13418), .Y(
        n34645) );
  OA22X1 U53037 ( .A0(net261981), .A1(n32480), .B0(n32488), .B1(n40084), .Y(
        n13417) );
  AOI222XL U53038 ( .A0(net265720), .A1(n50597), .B0(n40209), .B1(n50596),
        .C0(n40383), .C1(n50595), .Y(n13418) );
  OAI211X1 U53039 ( .A0(n32488), .A1(n42896), .B0(n13393), .C0(n13394), .Y(
        n34637) );
  OA22X1 U53040 ( .A0(net218424), .A1(n32472), .B0(n32480), .B1(n40084), .Y(
        n13393) );
  AOI222XL U53041 ( .A0(net265720), .A1(n50596), .B0(n40209), .B1(n50595),
        .C0(n40383), .C1(n50594), .Y(n13394) );
  OAI211X1 U53042 ( .A0(n32480), .A1(n42897), .B0(n13369), .C0(n13370), .Y(
        n34629) );
  OA22X1 U53043 ( .A0(net263216), .A1(n32464), .B0(n32472), .B1(n40083), .Y(
        n13369) );
  AOI222XL U53044 ( .A0(net265701), .A1(n50595), .B0(n40210), .B1(n50594),
        .C0(n40384), .C1(n50593), .Y(n13370) );
  OAI211X1 U53045 ( .A0(n32472), .A1(n42898), .B0(n13345), .C0(n13346), .Y(
        n34621) );
  OA22X1 U53046 ( .A0(net263216), .A1(n32456), .B0(n32464), .B1(n40083), .Y(
        n13345) );
  AOI222XL U53047 ( .A0(net265701), .A1(n50594), .B0(n40210), .B1(n50593),
        .C0(n40384), .C1(n50592), .Y(n13346) );
  OAI211X1 U53048 ( .A0(n32464), .A1(n42899), .B0(n13321), .C0(n13322), .Y(
        n34613) );
  OA22X1 U53049 ( .A0(net263235), .A1(n32448), .B0(n32456), .B1(n40082), .Y(
        n13321) );
  AOI222XL U53050 ( .A0(net265701), .A1(n50593), .B0(n40211), .B1(n50592),
        .C0(n40384), .C1(n50591), .Y(n13322) );
  OAI211X1 U53051 ( .A0(n32456), .A1(n42900), .B0(n13297), .C0(n13298), .Y(
        n34605) );
  OA22X1 U53052 ( .A0(net263235), .A1(n32440), .B0(n32448), .B1(n40082), .Y(
        n13297) );
  AOI222XL U53053 ( .A0(net265682), .A1(n50592), .B0(n40211), .B1(n50591),
        .C0(n40385), .C1(n50590), .Y(n13298) );
  OAI211X1 U53054 ( .A0(n32448), .A1(n42902), .B0(n13273), .C0(n13274), .Y(
        n34597) );
  OA22X1 U53055 ( .A0(net263254), .A1(n32432), .B0(n32440), .B1(n40081), .Y(
        n13273) );
  AOI222XL U53056 ( .A0(net265682), .A1(n50591), .B0(n40211), .B1(n50590),
        .C0(n40385), .C1(n50589), .Y(n13274) );
  OAI211X1 U53057 ( .A0(n32440), .A1(n42903), .B0(n13249), .C0(n13250), .Y(
        n34589) );
  OA22X1 U53058 ( .A0(net263254), .A1(n32424), .B0(n32432), .B1(n40081), .Y(
        n13249) );
  AOI222XL U53059 ( .A0(net265682), .A1(n50590), .B0(n40212), .B1(n50589),
        .C0(n40385), .C1(n50588), .Y(n13250) );
  OAI211X1 U53060 ( .A0(n32432), .A1(n42904), .B0(n13225), .C0(n13226), .Y(
        n34581) );
  OA22X1 U53061 ( .A0(net218366), .A1(n32416), .B0(n32424), .B1(n40080), .Y(
        n13225) );
  AOI222XL U53062 ( .A0(net265245), .A1(n50589), .B0(n40212), .B1(n50588),
        .C0(net217056), .C1(n50587), .Y(n13226) );
  OAI211X1 U53063 ( .A0(n32424), .A1(n42905), .B0(n13201), .C0(n13202), .Y(
        n34573) );
  OA22X1 U53064 ( .A0(net218346), .A1(n32408), .B0(n32416), .B1(n40080), .Y(
        n13201) );
  AOI222XL U53065 ( .A0(net264979), .A1(n50588), .B0(n40213), .B1(n50587),
        .C0(net217036), .C1(n50586), .Y(n13202) );
  OAI211X1 U53066 ( .A0(n32416), .A1(n42906), .B0(n13177), .C0(n13178), .Y(
        n34565) );
  AOI222XL U53067 ( .A0(net265150), .A1(n50587), .B0(n40213), .B1(n50586),
        .C0(net217060), .C1(n50585), .Y(n13178) );
  OAI211X1 U53068 ( .A0(n32408), .A1(n42907), .B0(n13153), .C0(n13154), .Y(
        n34557) );
  AOI222XL U53069 ( .A0(net265644), .A1(n50586), .B0(n40213), .B1(n50585),
        .C0(n40381), .C1(n50584), .Y(n13154) );
  OAI211X1 U53070 ( .A0(n34417), .A1(n42910), .B0(n13049), .C0(n50074), .Y(
        n34525) );
  OAI222XL U53071 ( .A0(net266654), .A1(n9660), .B0(n40160), .B1(n9659), .C0(
        n40292), .C1(n34425), .Y(n13051) );
  CLKINVX1 U53072 ( .A(n19158), .Y(n49565) );
  OAI222XL U53073 ( .A0(net266381), .A1(n9659), .B0(n40174), .B1(n34425), .C0(
        n40303), .C1(n34417), .Y(n19158) );
  OA22X1 U53074 ( .A0(net262855), .A1(n34081), .B0(n34089), .B1(n40103), .Y(
        n18220) );
  AOI222XL U53075 ( .A0(net265302), .A1(n49512), .B0(n40235), .B1(n49511),
        .C0(net217108), .C1(n50582), .Y(n18221) );
  OAI211X1 U53076 ( .A0(n34089), .A1(n42828), .B0(n18196), .C0(n18197), .Y(
        n36238) );
  OA22X1 U53077 ( .A0(net262874), .A1(n34073), .B0(n34081), .B1(n40103), .Y(
        n18196) );
  AOI222XL U53078 ( .A0(net265283), .A1(n49511), .B0(n40189), .B1(n50582),
        .C0(n40318), .C1(n50581), .Y(n18197) );
  AOI222XL U53079 ( .A0(net265283), .A1(n50582), .B0(net218124), .B1(n50581),
        .C0(n40318), .C1(n50580), .Y(n18173) );
  AOI222XL U53080 ( .A0(net265283), .A1(n50581), .B0(n40236), .B1(n50580),
        .C0(n40318), .C1(n50579), .Y(n18149) );
  AOI222XL U53081 ( .A0(net265264), .A1(n50580), .B0(n40236), .B1(n50579),
        .C0(n40319), .C1(n50578), .Y(n18125) );
  AOI222XL U53082 ( .A0(net265264), .A1(n50579), .B0(n40236), .B1(n50578),
        .C0(n40319), .C1(n50577), .Y(n18101) );
  AOI222XL U53083 ( .A0(net265264), .A1(n50578), .B0(n40237), .B1(n50577),
        .C0(n40319), .C1(n50576), .Y(n18077) );
  AOI222XL U53084 ( .A0(net265245), .A1(n50577), .B0(n40237), .B1(n50576),
        .C0(n40320), .C1(n50575), .Y(n18053) );
  AOI222XL U53085 ( .A0(net265245), .A1(n50576), .B0(n40238), .B1(n50575),
        .C0(n40320), .C1(n50574), .Y(n18029) );
  AOI222XL U53086 ( .A0(net265245), .A1(n50575), .B0(n40238), .B1(n50574),
        .C0(n40320), .C1(n50573), .Y(n18005) );
  AOI222XL U53087 ( .A0(net265226), .A1(n50574), .B0(n40238), .B1(n50573),
        .C0(n40321), .C1(n50572), .Y(n17981) );
  AOI222XL U53088 ( .A0(net265226), .A1(n50573), .B0(n40239), .B1(n50572),
        .C0(n40321), .C1(n50571), .Y(n17957) );
  AOI222XL U53089 ( .A0(net265226), .A1(n50572), .B0(n40239), .B1(n50571),
        .C0(n40321), .C1(n50570), .Y(n17933) );
  AOI222XL U53090 ( .A0(net265207), .A1(n50571), .B0(n40240), .B1(n50570),
        .C0(n40322), .C1(n50569), .Y(n17909) );
  AOI222XL U53091 ( .A0(net265207), .A1(n50570), .B0(n40240), .B1(n50569),
        .C0(n40322), .C1(n50568), .Y(n17885) );
  AOI222XL U53092 ( .A0(net265207), .A1(n50569), .B0(n40241), .B1(n50568),
        .C0(n40322), .C1(n50567), .Y(n17861) );
  AOI222XL U53093 ( .A0(net265188), .A1(n50568), .B0(n40241), .B1(n50567),
        .C0(n40323), .C1(n50566), .Y(n17837) );
  AOI222XL U53094 ( .A0(net265188), .A1(n50567), .B0(n40241), .B1(n50566),
        .C0(n40323), .C1(n50565), .Y(n17813) );
  AOI222XL U53095 ( .A0(net265188), .A1(n50566), .B0(n40242), .B1(n50565),
        .C0(n40324), .C1(n50564), .Y(n17789) );
  AOI222XL U53096 ( .A0(net265169), .A1(n50565), .B0(n40242), .B1(n50564),
        .C0(n40324), .C1(n50563), .Y(n17765) );
  AOI222XL U53097 ( .A0(net265169), .A1(n50564), .B0(n40243), .B1(n50563),
        .C0(n40324), .C1(n50562), .Y(n17741) );
  AOI222XL U53098 ( .A0(net265169), .A1(n50563), .B0(n40243), .B1(n50562),
        .C0(n40325), .C1(n50561), .Y(n17717) );
  AOI222XL U53099 ( .A0(net265150), .A1(n50562), .B0(n40243), .B1(n50561),
        .C0(n40325), .C1(n50560), .Y(n17693) );
  AOI222XL U53100 ( .A0(net265150), .A1(n50561), .B0(n40244), .B1(n50560),
        .C0(n40325), .C1(n50559), .Y(n17669) );
  AOI222XL U53101 ( .A0(net265150), .A1(n50560), .B0(n40244), .B1(n50559),
        .C0(net217102), .C1(n50558), .Y(n17645) );
  AOI222XL U53102 ( .A0(net265131), .A1(n50559), .B0(n40245), .B1(n50558),
        .C0(net217094), .C1(n50557), .Y(n17621) );
  AOI222XL U53103 ( .A0(net265131), .A1(n50558), .B0(n40245), .B1(n50557),
        .C0(net217100), .C1(n50556), .Y(n17597) );
  AOI222XL U53104 ( .A0(net265473), .A1(n50557), .B0(n40225), .B1(n50556),
        .C0(n40326), .C1(n50555), .Y(n17573) );
  AOI222XL U53105 ( .A0(net265454), .A1(n50556), .B0(n40225), .B1(n50555),
        .C0(n40326), .C1(n50554), .Y(n17549) );
  AOI222XL U53106 ( .A0(net265454), .A1(n50555), .B0(n40226), .B1(n50554),
        .C0(n40326), .C1(n50553), .Y(n17525) );
  AOI222XL U53107 ( .A0(net265454), .A1(n50554), .B0(n40226), .B1(n50553),
        .C0(n40327), .C1(n50552), .Y(n17501) );
  AOI222XL U53108 ( .A0(net265435), .A1(n50553), .B0(n40227), .B1(n50552),
        .C0(n40327), .C1(n50551), .Y(n17477) );
  AOI222XL U53109 ( .A0(net265435), .A1(n50552), .B0(n40227), .B1(n50551),
        .C0(n40327), .C1(n50550), .Y(n17453) );
  AOI222XL U53110 ( .A0(net265435), .A1(n50551), .B0(n40227), .B1(n50550),
        .C0(n40328), .C1(n50549), .Y(n17429) );
  AOI222XL U53111 ( .A0(net265416), .A1(n50550), .B0(n40228), .B1(n50549),
        .C0(n40328), .C1(n50548), .Y(n17405) );
  AOI222XL U53112 ( .A0(net265416), .A1(n50549), .B0(n40228), .B1(n50548),
        .C0(n40329), .C1(n50547), .Y(n17381) );
  AOI222XL U53113 ( .A0(net265416), .A1(n50548), .B0(n40229), .B1(n50547),
        .C0(n40329), .C1(n50546), .Y(n17357) );
  AOI222XL U53114 ( .A0(net265397), .A1(n50547), .B0(n40229), .B1(n50546),
        .C0(n40329), .C1(n50545), .Y(n17333) );
  AOI222XL U53115 ( .A0(net265397), .A1(n50546), .B0(n40229), .B1(n50545),
        .C0(n40330), .C1(n50544), .Y(n17309) );
  AOI222XL U53116 ( .A0(net265397), .A1(n50545), .B0(n40230), .B1(n50544),
        .C0(n40330), .C1(n50543), .Y(n17285) );
  AOI222XL U53117 ( .A0(net265378), .A1(n50544), .B0(n40230), .B1(n50543),
        .C0(n40330), .C1(n50542), .Y(n17261) );
  AOI222XL U53118 ( .A0(net265378), .A1(n50543), .B0(n40231), .B1(n50542),
        .C0(n40331), .C1(n50541), .Y(n17237) );
  AOI222XL U53119 ( .A0(net265378), .A1(n50542), .B0(n40231), .B1(n50541),
        .C0(n40331), .C1(n50540), .Y(n17213) );
  AOI222XL U53120 ( .A0(net265359), .A1(n50541), .B0(n40231), .B1(n50540),
        .C0(n40331), .C1(n50539), .Y(n17189) );
  AOI222XL U53121 ( .A0(net265359), .A1(n50540), .B0(n40232), .B1(n50539),
        .C0(n40332), .C1(n50538), .Y(n17165) );
  AOI222XL U53122 ( .A0(net265359), .A1(n50539), .B0(n40232), .B1(n50538),
        .C0(n40332), .C1(n50537), .Y(n17141) );
  AOI222XL U53123 ( .A0(net265340), .A1(n50538), .B0(n40233), .B1(n50537),
        .C0(n40332), .C1(n50536), .Y(n17117) );
  AOI222XL U53124 ( .A0(net265340), .A1(n50537), .B0(n40233), .B1(n50536),
        .C0(n40333), .C1(n50535), .Y(n17093) );
  AOI222XL U53125 ( .A0(net265340), .A1(n50536), .B0(n40233), .B1(n50535),
        .C0(n40333), .C1(n50534), .Y(n17069) );
  AOI222XL U53126 ( .A0(net265321), .A1(n50535), .B0(n40234), .B1(n50534),
        .C0(n40333), .C1(n50533), .Y(n17045) );
  AOI222XL U53127 ( .A0(net265321), .A1(n50534), .B0(n40234), .B1(n50533),
        .C0(n40334), .C1(n50532), .Y(n17021) );
  AOI222XL U53128 ( .A0(net265321), .A1(n50533), .B0(n40235), .B1(n50532),
        .C0(n40334), .C1(n50531), .Y(n16997) );
  AOI222XL U53129 ( .A0(net265302), .A1(n50532), .B0(n40235), .B1(n50531),
        .C0(n40335), .C1(n50530), .Y(n16973) );
  AOI222XL U53130 ( .A0(net265378), .A1(n50531), .B0(n40256), .B1(n50530),
        .C0(n40335), .C1(n50529), .Y(n16949) );
  AOI222XL U53131 ( .A0(net264960), .A1(n50530), .B0(n40256), .B1(n50529),
        .C0(n40335), .C1(n50528), .Y(n16925) );
  AOI222XL U53132 ( .A0(net264941), .A1(n50529), .B0(n40257), .B1(n50528),
        .C0(n40336), .C1(n50527), .Y(n16901) );
  AOI222XL U53133 ( .A0(net264941), .A1(n50528), .B0(n40257), .B1(n50527),
        .C0(n40336), .C1(n50526), .Y(n16877) );
  AOI222XL U53134 ( .A0(net264941), .A1(n50527), .B0(n40257), .B1(n50526),
        .C0(n40336), .C1(n50525), .Y(n16853) );
  AOI222XL U53135 ( .A0(net264922), .A1(n50526), .B0(n40258), .B1(n50525),
        .C0(n40337), .C1(n50524), .Y(n16829) );
  AOI222XL U53136 ( .A0(net264922), .A1(n50525), .B0(n40258), .B1(n50524),
        .C0(n40337), .C1(n50523), .Y(n16805) );
  AOI222XL U53137 ( .A0(net264922), .A1(n50524), .B0(n40259), .B1(n50523),
        .C0(n40337), .C1(n50522), .Y(n16781) );
  AOI222XL U53138 ( .A0(net264903), .A1(n50523), .B0(n40259), .B1(n50522),
        .C0(n40338), .C1(n50521), .Y(n16757) );
  AOI222XL U53139 ( .A0(net264903), .A1(n50522), .B0(n40259), .B1(n50521),
        .C0(n40338), .C1(n50520), .Y(n16733) );
  AOI222XL U53140 ( .A0(net264903), .A1(n50521), .B0(n40260), .B1(n50520),
        .C0(n40338), .C1(n50519), .Y(n16709) );
  AOI222XL U53141 ( .A0(net264884), .A1(n50520), .B0(n40260), .B1(n50519),
        .C0(n40339), .C1(n50518), .Y(n16685) );
  AOI222XL U53142 ( .A0(net264884), .A1(n50519), .B0(n40261), .B1(n50518),
        .C0(n40339), .C1(n50517), .Y(n16661) );
  AOI222XL U53143 ( .A0(net264884), .A1(n50518), .B0(n40261), .B1(n50517),
        .C0(n40339), .C1(n50516), .Y(n16637) );
  AOI222XL U53144 ( .A0(net264808), .A1(n50517), .B0(n40266), .B1(n50516),
        .C0(n40340), .C1(n50515), .Y(n16613) );
  AOI222XL U53145 ( .A0(net264884), .A1(n50516), .B0(n40266), .B1(n50515),
        .C0(n40340), .C1(n50514), .Y(n16589) );
  AOI222XL U53146 ( .A0(net264808), .A1(n50515), .B0(n40265), .B1(n50514),
        .C0(n40341), .C1(n50513), .Y(n16565) );
  AOI222XL U53147 ( .A0(net264808), .A1(n50514), .B0(n40265), .B1(n50513),
        .C0(n40341), .C1(n50512), .Y(n16541) );
  AOI222XL U53148 ( .A0(net264827), .A1(n50513), .B0(n40265), .B1(n50512),
        .C0(n40341), .C1(n50511), .Y(n16517) );
  AOI222XL U53149 ( .A0(net264827), .A1(n50512), .B0(n40264), .B1(n50511),
        .C0(n40342), .C1(n50510), .Y(n16493) );
  AOI222XL U53150 ( .A0(net264827), .A1(n50511), .B0(n40264), .B1(n50510),
        .C0(n40342), .C1(n50509), .Y(n16469) );
  AOI222XL U53151 ( .A0(net264846), .A1(n50510), .B0(n40263), .B1(n50509),
        .C0(n40342), .C1(n50508), .Y(n16445) );
  AOI222XL U53152 ( .A0(net264846), .A1(n50509), .B0(n40263), .B1(n50508),
        .C0(n40343), .C1(n50507), .Y(n16421) );
  AOI222XL U53153 ( .A0(net264846), .A1(n50508), .B0(n40262), .B1(n50507),
        .C0(n40343), .C1(n50506), .Y(n16397) );
  AOI222XL U53154 ( .A0(net264865), .A1(n50507), .B0(n40262), .B1(n50506),
        .C0(n40343), .C1(n50505), .Y(n16373) );
  AOI222XL U53155 ( .A0(net264865), .A1(n50506), .B0(n40262), .B1(n50505),
        .C0(n40344), .C1(n50504), .Y(n16349) );
  AOI222XL U53156 ( .A0(net264865), .A1(n50505), .B0(n40261), .B1(n50504),
        .C0(n40344), .C1(n50503), .Y(n16325) );
  AOI222XL U53157 ( .A0(net265131), .A1(n50504), .B0(n40245), .B1(n50503),
        .C0(n40344), .C1(n50502), .Y(n16301) );
  AOI222XL U53158 ( .A0(net265131), .A1(n50503), .B0(n40246), .B1(n50502),
        .C0(n40345), .C1(n50501), .Y(n16277) );
  AOI222XL U53159 ( .A0(net265112), .A1(n50502), .B0(n40246), .B1(n50501),
        .C0(n40345), .C1(n50500), .Y(n16253) );
  AOI222XL U53160 ( .A0(net265112), .A1(n50501), .B0(n40246), .B1(n50500),
        .C0(n40345), .C1(n50499), .Y(n16229) );
  AOI222XL U53161 ( .A0(net265112), .A1(n50500), .B0(n40247), .B1(n50499),
        .C0(n40346), .C1(n50498), .Y(n16205) );
  AOI222XL U53162 ( .A0(net221818), .A1(n50499), .B0(n40247), .B1(n50498),
        .C0(n40346), .C1(n50497), .Y(n16181) );
  AOI222XL U53163 ( .A0(net221804), .A1(n50498), .B0(n40248), .B1(n50497),
        .C0(n40347), .C1(n50496), .Y(n16157) );
  AOI222XL U53164 ( .A0(net221820), .A1(n50497), .B0(n40248), .B1(n50496),
        .C0(n40347), .C1(n50495), .Y(n16133) );
  AOI222XL U53165 ( .A0(net265074), .A1(n50496), .B0(n40248), .B1(n50495),
        .C0(n40347), .C1(n37251), .Y(n16109) );
  AOI222XL U53166 ( .A0(net265074), .A1(n50495), .B0(n40249), .B1(n37251),
        .C0(n40348), .C1(n50494), .Y(n16085) );
  AOI222XL U53167 ( .A0(net265074), .A1(n37251), .B0(n40249), .B1(n50494),
        .C0(n40348), .C1(n50493), .Y(n16061) );
  AOI222XL U53168 ( .A0(net265055), .A1(n50494), .B0(n40250), .B1(n50493),
        .C0(n40348), .C1(n50492), .Y(n16037) );
  AOI222XL U53169 ( .A0(net265055), .A1(n50493), .B0(n40250), .B1(n50492),
        .C0(n40349), .C1(n50491), .Y(n16013) );
  AOI222XL U53170 ( .A0(net265036), .A1(n50492), .B0(n40251), .B1(n50491),
        .C0(n40349), .C1(n50490), .Y(n15989) );
  AOI222XL U53171 ( .A0(net265036), .A1(n50491), .B0(n40251), .B1(n50490),
        .C0(n40349), .C1(n50489), .Y(n15965) );
  AOI222XL U53172 ( .A0(net265036), .A1(n50490), .B0(n40251), .B1(n50489),
        .C0(n40382), .C1(n50488), .Y(n15941) );
  AOI222XL U53173 ( .A0(net265017), .A1(n50489), .B0(n40252), .B1(n50488),
        .C0(n40382), .C1(n37252), .Y(n15917) );
  AOI222XL U53174 ( .A0(net265017), .A1(n50488), .B0(n40252), .B1(n37252),
        .C0(n40382), .C1(n50487), .Y(n15893) );
  AOI222XL U53175 ( .A0(net265017), .A1(n37252), .B0(n40253), .B1(n50487),
        .C0(n40350), .C1(n50486), .Y(n15869) );
  AOI222XL U53176 ( .A0(net264998), .A1(n50487), .B0(n40253), .B1(n50486),
        .C0(n40350), .C1(n50485), .Y(n15845) );
  AOI222XL U53177 ( .A0(net264998), .A1(n50486), .B0(n40253), .B1(n50485),
        .C0(n40350), .C1(n50484), .Y(n15821) );
  AOI222XL U53178 ( .A0(net264998), .A1(n50485), .B0(n40254), .B1(n50484),
        .C0(net217036), .C1(n50483), .Y(n15797) );
  AOI222XL U53179 ( .A0(net264979), .A1(n50484), .B0(n40254), .B1(n50483),
        .C0(net217036), .C1(n50482), .Y(n15773) );
  AOI222XL U53180 ( .A0(net264979), .A1(n50483), .B0(n40255), .B1(n50482),
        .C0(n40351), .C1(n50481), .Y(n15749) );
  AOI222XL U53181 ( .A0(net264979), .A1(n50482), .B0(n40255), .B1(n50481),
        .C0(n40351), .C1(n50480), .Y(n15725) );
  AOI222XL U53182 ( .A0(net264960), .A1(n50481), .B0(n40255), .B1(n50480),
        .C0(n40351), .C1(n50479), .Y(n15701) );
  AOI222XL U53183 ( .A0(net264960), .A1(n50480), .B0(n40250), .B1(n50479),
        .C0(n40352), .C1(n50478), .Y(n15677) );
  AOI222XL U53184 ( .A0(net265967), .A1(n50479), .B0(n40193), .B1(n50478),
        .C0(n40352), .C1(n50477), .Y(n15653) );
  AOI222XL U53185 ( .A0(net265967), .A1(n50478), .B0(n40193), .B1(n50477),
        .C0(n40352), .C1(n50476), .Y(n15629) );
  AOI222XL U53186 ( .A0(net265967), .A1(n50477), .B0(n40194), .B1(n50476),
        .C0(n40353), .C1(n50475), .Y(n15605) );
  AOI222XL U53187 ( .A0(net265948), .A1(n50476), .B0(n40194), .B1(n50475),
        .C0(n40353), .C1(n50474), .Y(n15581) );
  AOI222XL U53188 ( .A0(net265948), .A1(n50475), .B0(n40195), .B1(n50474),
        .C0(n40353), .C1(n50473), .Y(n15557) );
  AOI222XL U53189 ( .A0(net265948), .A1(n50474), .B0(n40195), .B1(n50473),
        .C0(n40354), .C1(n50472), .Y(n15533) );
  AOI222XL U53190 ( .A0(net265929), .A1(n50473), .B0(n40195), .B1(n50472),
        .C0(n40354), .C1(n50471), .Y(n15509) );
  AOI222XL U53191 ( .A0(net265929), .A1(n50472), .B0(n40196), .B1(n50471),
        .C0(n40354), .C1(n50470), .Y(n15485) );
  AOI222XL U53192 ( .A0(net265929), .A1(n50471), .B0(n40196), .B1(n50470),
        .C0(n40355), .C1(n50469), .Y(n15461) );
  AOI222XL U53193 ( .A0(net265910), .A1(n50470), .B0(n40197), .B1(n50469),
        .C0(n40355), .C1(n50468), .Y(n15437) );
  AOI222XL U53194 ( .A0(net265910), .A1(n50469), .B0(n40197), .B1(n50468),
        .C0(n40355), .C1(n50467), .Y(n15413) );
  AOI222XL U53195 ( .A0(net265910), .A1(n50468), .B0(n40197), .B1(n50467),
        .C0(n40356), .C1(n50466), .Y(n15389) );
  AOI222XL U53196 ( .A0(net265891), .A1(n50467), .B0(n40198), .B1(n50466),
        .C0(n40356), .C1(n50465), .Y(n15365) );
  AOI222XL U53197 ( .A0(net265891), .A1(n50466), .B0(n40198), .B1(n50465),
        .C0(n40357), .C1(n50464), .Y(n15341) );
  AOI222XL U53198 ( .A0(net265891), .A1(n50465), .B0(n40199), .B1(n50464),
        .C0(n40357), .C1(n50463), .Y(n15317) );
  AOI222XL U53199 ( .A0(net265872), .A1(n50464), .B0(n40199), .B1(n50463),
        .C0(n40357), .C1(n50462), .Y(n15293) );
  AOI222XL U53200 ( .A0(net265872), .A1(n50463), .B0(n40199), .B1(n50462),
        .C0(n40358), .C1(n50461), .Y(n15269) );
  AOI222XL U53201 ( .A0(net265872), .A1(n50462), .B0(n40200), .B1(n50461),
        .C0(n40358), .C1(n50460), .Y(n15245) );
  AOI222XL U53202 ( .A0(net265853), .A1(n50461), .B0(n40200), .B1(n50460),
        .C0(n40358), .C1(n50459), .Y(n15221) );
  AOI222XL U53203 ( .A0(net265853), .A1(n50460), .B0(n40201), .B1(n50459),
        .C0(n40359), .C1(n50458), .Y(n15197) );
  AOI222XL U53204 ( .A0(net265853), .A1(n50459), .B0(n40201), .B1(n50458),
        .C0(n40359), .C1(n50457), .Y(n15173) );
  AOI222XL U53205 ( .A0(net265834), .A1(n50458), .B0(n40201), .B1(n50457),
        .C0(n40359), .C1(n50456), .Y(n15149) );
  AOI222XL U53206 ( .A0(net265834), .A1(n50457), .B0(n40202), .B1(n50456),
        .C0(n40360), .C1(n37243), .Y(n15125) );
  AOI222XL U53207 ( .A0(net265834), .A1(n50456), .B0(n40202), .B1(n37243),
        .C0(n40360), .C1(n37019), .Y(n15101) );
  AOI222XL U53208 ( .A0(net265815), .A1(n37243), .B0(n40203), .B1(n37019),
        .C0(n40360), .C1(n36930), .Y(n15077) );
  AOI222XL U53209 ( .A0(net265815), .A1(n37019), .B0(n40203), .B1(n36930),
        .C0(net217026), .C1(n50455), .Y(n15053) );
  AOI222XL U53210 ( .A0(net221892), .A1(n50454), .B0(n40184), .B1(n50453),
        .C0(n40361), .C1(n36931), .Y(n14981) );
  AOI222XL U53211 ( .A0(net266119), .A1(n50453), .B0(n40184), .B1(n36931),
        .C0(n40361), .C1(n37244), .Y(n14957) );
  AOI222XL U53212 ( .A0(net266119), .A1(n36931), .B0(n40185), .B1(n37244),
        .C0(n40362), .C1(n37020), .Y(n14933) );
  AOI222XL U53213 ( .A0(net266119), .A1(n37244), .B0(n40185), .B1(n37020),
        .C0(n40362), .C1(n36925), .Y(n14909) );
  OA22X1 U53214 ( .A0(net263767), .A1(n32969), .B0(n32977), .B1(n40053), .Y(
        n14884) );
  AOI222XL U53215 ( .A0(net266100), .A1(n37020), .B0(n40185), .B1(n36925),
        .C0(n40362), .C1(n37245), .Y(n14885) );
  OA22X1 U53216 ( .A0(net263767), .A1(n32961), .B0(n32969), .B1(n40052), .Y(
        n14860) );
  AOI222XL U53217 ( .A0(net266100), .A1(n36925), .B0(net218110), .B1(n37245),
        .C0(n40363), .C1(n36946), .Y(n14861) );
  OA22X1 U53218 ( .A0(net218472), .A1(n32953), .B0(n32961), .B1(n40052), .Y(
        n14836) );
  AOI222XL U53219 ( .A0(net266100), .A1(n37245), .B0(net218132), .B1(n36946),
        .C0(n40363), .C1(n50452), .Y(n14837) );
  OA22X1 U53220 ( .A0(net218468), .A1(n32945), .B0(n32953), .B1(n40051), .Y(
        n14812) );
  AOI222XL U53221 ( .A0(net266081), .A1(n36946), .B0(n40186), .B1(n50452),
        .C0(n40363), .C1(n50451), .Y(n14813) );
  OAI211X1 U53222 ( .A0(n32953), .A1(n42974), .B0(n14788), .C0(n14789), .Y(
        n35102) );
  OA22X1 U53223 ( .A0(net262912), .A1(n32937), .B0(n32945), .B1(n40051), .Y(
        n14788) );
  AOI222XL U53224 ( .A0(net266081), .A1(n50452), .B0(n40186), .B1(n50451),
        .C0(n40365), .C1(n50450), .Y(n14789) );
  OAI211X1 U53225 ( .A0(n32937), .A1(n42961), .B0(n14740), .C0(n14741), .Y(
        n35086) );
  OA22X1 U53226 ( .A0(net263805), .A1(n32921), .B0(n32929), .B1(n40050), .Y(
        n14740) );
  AOI222XL U53227 ( .A0(net266062), .A1(n50450), .B0(n40187), .B1(n50449),
        .C0(n40364), .C1(n50448), .Y(n14741) );
  OAI211X1 U53228 ( .A0(n32929), .A1(n42962), .B0(n14716), .C0(n14717), .Y(
        n35078) );
  OA22X1 U53229 ( .A0(net263824), .A1(n32913), .B0(n32921), .B1(n40049), .Y(
        n14716) );
  AOI222XL U53230 ( .A0(net266062), .A1(n50449), .B0(n40187), .B1(n50448),
        .C0(n40364), .C1(n50447), .Y(n14717) );
  OAI211X1 U53231 ( .A0(n32921), .A1(n42963), .B0(n14692), .C0(n14693), .Y(
        n35070) );
  OA22X1 U53232 ( .A0(net263824), .A1(n32905), .B0(n32913), .B1(n40049), .Y(
        n14692) );
  AOI222XL U53233 ( .A0(net266062), .A1(n50448), .B0(n40188), .B1(n50447),
        .C0(n40364), .C1(n50446), .Y(n14693) );
  OAI211X1 U53234 ( .A0(n32913), .A1(n42964), .B0(n14668), .C0(n14669), .Y(
        n35062) );
  OA22X1 U53235 ( .A0(net263843), .A1(n32897), .B0(n32905), .B1(n40048), .Y(
        n14668) );
  AOI222XL U53236 ( .A0(net266043), .A1(n50447), .B0(n40188), .B1(n50446),
        .C0(n40364), .C1(n50445), .Y(n14669) );
  OAI211X1 U53237 ( .A0(n32905), .A1(n42965), .B0(n14644), .C0(n14645), .Y(
        n35054) );
  OA22X1 U53238 ( .A0(net263843), .A1(n32889), .B0(n32897), .B1(n40048), .Y(
        n14644) );
  AOI222XL U53239 ( .A0(net266043), .A1(n50446), .B0(n40189), .B1(n50445),
        .C0(n40365), .C1(n50444), .Y(n14645) );
  OA22X1 U53240 ( .A0(net263862), .A1(n32881), .B0(n32889), .B1(n40047), .Y(
        n14620) );
  AOI222XL U53241 ( .A0(net266043), .A1(n50445), .B0(n40189), .B1(n50444),
        .C0(n40365), .C1(n50443), .Y(n14621) );
  OA22X1 U53242 ( .A0(net263862), .A1(n32873), .B0(n32881), .B1(n40047), .Y(
        n14596) );
  AOI222XL U53243 ( .A0(net266024), .A1(n50444), .B0(n40189), .B1(n50443),
        .C0(n40365), .C1(n50442), .Y(n14597) );
  OA22X1 U53244 ( .A0(net218564), .A1(n32865), .B0(n32873), .B1(n40084), .Y(
        n14572) );
  AOI222XL U53245 ( .A0(net266024), .A1(n50443), .B0(n40190), .B1(n50442),
        .C0(n40366), .C1(n50441), .Y(n14573) );
  OAI211X1 U53246 ( .A0(n32873), .A1(n42970), .B0(n14548), .C0(n14549), .Y(
        n35022) );
  OA22X1 U53247 ( .A0(net263064), .A1(n32857), .B0(n32865), .B1(n40092), .Y(
        n14548) );
  AOI222XL U53248 ( .A0(net266024), .A1(n50442), .B0(n40190), .B1(n50441),
        .C0(n40366), .C1(n50440), .Y(n14549) );
  OA22X1 U53249 ( .A0(net263083), .A1(n32849), .B0(n32857), .B1(n40091), .Y(
        n14524) );
  AOI222XL U53250 ( .A0(net266005), .A1(n50441), .B0(n40191), .B1(n50440),
        .C0(n40367), .C1(n50439), .Y(n14525) );
  OAI211X1 U53251 ( .A0(n32857), .A1(n42972), .B0(n14500), .C0(n14501), .Y(
        n35006) );
  OA22X1 U53252 ( .A0(net263083), .A1(n32841), .B0(n32849), .B1(n40091), .Y(
        n14500) );
  AOI222XL U53253 ( .A0(net266005), .A1(n50440), .B0(n40191), .B1(n50439),
        .C0(n40367), .C1(n50438), .Y(n14501) );
  OAI211X1 U53254 ( .A0(n32849), .A1(n42973), .B0(n14476), .C0(n14477), .Y(
        n34998) );
  OA22X1 U53255 ( .A0(net263102), .A1(n32833), .B0(n32841), .B1(n40090), .Y(
        n14476) );
  AOI222XL U53256 ( .A0(net266005), .A1(n50439), .B0(n40191), .B1(n50438),
        .C0(n40367), .C1(n50437), .Y(n14477) );
  OAI211X1 U53257 ( .A0(n32841), .A1(n42975), .B0(n14452), .C0(n14453), .Y(
        n34990) );
  OA22X1 U53258 ( .A0(net263102), .A1(n32825), .B0(n32833), .B1(n40090), .Y(
        n14452) );
  AOI222XL U53259 ( .A0(net221852), .A1(n50438), .B0(n40192), .B1(n50437),
        .C0(n40368), .C1(n50436), .Y(n14453) );
  OAI211X1 U53260 ( .A0(n32833), .A1(n42976), .B0(n14428), .C0(n14429), .Y(
        n34982) );
  OA22X1 U53261 ( .A0(net263102), .A1(n32817), .B0(n32825), .B1(n40089), .Y(
        n14428) );
  AOI222XL U53262 ( .A0(net221834), .A1(n50437), .B0(n40192), .B1(n50436),
        .C0(n40368), .C1(n50435), .Y(n14429) );
  OAI211X1 U53263 ( .A0(n32825), .A1(n42880), .B0(n14404), .C0(n14405), .Y(
        n34974) );
  OA22X1 U53264 ( .A0(net263121), .A1(n32809), .B0(n32817), .B1(n40089), .Y(
        n14404) );
  AOI222XL U53265 ( .A0(net221832), .A1(n50436), .B0(n40193), .B1(n50435),
        .C0(n40368), .C1(n50434), .Y(n14405) );
  OAI211X1 U53266 ( .A0(n32817), .A1(n42881), .B0(n14380), .C0(n14381), .Y(
        n34966) );
  OA22X1 U53267 ( .A0(net263121), .A1(n32801), .B0(n32809), .B1(n40088), .Y(
        n14380) );
  AOI222XL U53268 ( .A0(net265644), .A1(n50435), .B0(n40214), .B1(n50434),
        .C0(n40369), .C1(n50433), .Y(n14381) );
  OAI211X1 U53269 ( .A0(n32809), .A1(n42882), .B0(n14356), .C0(n14357), .Y(
        n34958) );
  OA22X1 U53270 ( .A0(net263140), .A1(n32793), .B0(n32801), .B1(n40088), .Y(
        n14356) );
  AOI222XL U53271 ( .A0(net265625), .A1(n50434), .B0(n40215), .B1(n50433),
        .C0(n40369), .C1(n50432), .Y(n14357) );
  OA22X1 U53272 ( .A0(net263140), .A1(n32785), .B0(n32793), .B1(n40087), .Y(
        n14332) );
  AOI222XL U53273 ( .A0(net265625), .A1(n50433), .B0(n40215), .B1(n50432),
        .C0(n40369), .C1(n50431), .Y(n14333) );
  OAI211X1 U53274 ( .A0(n32793), .A1(n42884), .B0(n14308), .C0(n14309), .Y(
        n34942) );
  OA22X1 U53275 ( .A0(net263159), .A1(n32777), .B0(n32785), .B1(n40087), .Y(
        n14308) );
  AOI222XL U53276 ( .A0(net265625), .A1(n50432), .B0(n40215), .B1(n50431),
        .C0(n40370), .C1(n50430), .Y(n14309) );
  OAI211X1 U53277 ( .A0(n32785), .A1(n42885), .B0(n14284), .C0(n14285), .Y(
        n34934) );
  OA22X1 U53278 ( .A0(net263159), .A1(n32769), .B0(n32777), .B1(n40086), .Y(
        n14284) );
  AOI222XL U53279 ( .A0(net265606), .A1(n50431), .B0(n40216), .B1(n50430),
        .C0(n40370), .C1(n50429), .Y(n14285) );
  OAI211X1 U53280 ( .A0(n32777), .A1(n42887), .B0(n14260), .C0(n14261), .Y(
        n34926) );
  OA22X1 U53281 ( .A0(net263178), .A1(n32761), .B0(n32769), .B1(n40086), .Y(
        n14260) );
  AOI222XL U53282 ( .A0(net265606), .A1(n50430), .B0(n40216), .B1(n50429),
        .C0(n40370), .C1(n50428), .Y(n14261) );
  OA22X1 U53283 ( .A0(net263178), .A1(n32753), .B0(n32761), .B1(n40085), .Y(
        n14236) );
  AOI222XL U53284 ( .A0(net265606), .A1(n50429), .B0(n40217), .B1(n50428),
        .C0(n40371), .C1(n50427), .Y(n14237) );
  OA22X1 U53285 ( .A0(net263178), .A1(n32745), .B0(n32753), .B1(n40085), .Y(
        n14212) );
  AOI222XL U53286 ( .A0(net265587), .A1(n50428), .B0(n40217), .B1(n50427),
        .C0(n40371), .C1(n50426), .Y(n14213) );
  OA22X1 U53287 ( .A0(net262988), .A1(n32737), .B0(n32745), .B1(n40096), .Y(
        n14188) );
  AOI222XL U53288 ( .A0(net265587), .A1(n50427), .B0(n40217), .B1(n50426),
        .C0(n40371), .C1(n50425), .Y(n14189) );
  OAI211X1 U53289 ( .A0(n32745), .A1(n42891), .B0(n14164), .C0(n14165), .Y(
        n34894) );
  OA22X1 U53290 ( .A0(net262931), .A1(n32729), .B0(n32737), .B1(n40100), .Y(
        n14164) );
  AOI222XL U53291 ( .A0(net265587), .A1(n50426), .B0(n40218), .B1(n50425),
        .C0(n40372), .C1(n50424), .Y(n14165) );
  OAI211X1 U53292 ( .A0(n32737), .A1(n42892), .B0(n14140), .C0(n14141), .Y(
        n34886) );
  OA22X1 U53293 ( .A0(net262950), .A1(n32721), .B0(n32729), .B1(n40099), .Y(
        n14140) );
  AOI222XL U53294 ( .A0(net265568), .A1(n50425), .B0(n40218), .B1(n50424),
        .C0(n40372), .C1(n50423), .Y(n14141) );
  OAI211X1 U53295 ( .A0(n32729), .A1(n42894), .B0(n14116), .C0(n14117), .Y(
        n34878) );
  OA22X1 U53296 ( .A0(net262950), .A1(n32713), .B0(n32721), .B1(n40099), .Y(
        n14116) );
  AOI222XL U53297 ( .A0(net265568), .A1(n50424), .B0(n40219), .B1(n50423),
        .C0(n40373), .C1(n50422), .Y(n14117) );
  OAI211X1 U53298 ( .A0(n32721), .A1(n42895), .B0(n14092), .C0(n14093), .Y(
        n34870) );
  OA22X1 U53299 ( .A0(net262950), .A1(n32705), .B0(n32713), .B1(n40098), .Y(
        n14092) );
  AOI222XL U53300 ( .A0(net265568), .A1(n50423), .B0(n40219), .B1(n50422),
        .C0(n40373), .C1(n50421), .Y(n14093) );
  OA22X1 U53301 ( .A0(net262969), .A1(n32697), .B0(n32705), .B1(n40098), .Y(
        n14068) );
  AOI222XL U53302 ( .A0(net265549), .A1(n50422), .B0(n40219), .B1(n50421),
        .C0(n40373), .C1(n50420), .Y(n14069) );
  OAI211X1 U53303 ( .A0(n32705), .A1(n42865), .B0(n14044), .C0(n14045), .Y(
        n34854) );
  OA22X1 U53304 ( .A0(net262969), .A1(n32689), .B0(n32697), .B1(n40097), .Y(
        n14044) );
  AOI222XL U53305 ( .A0(net265549), .A1(n50421), .B0(n40220), .B1(n50420),
        .C0(n40374), .C1(n50419), .Y(n14045) );
  OAI211X1 U53306 ( .A0(n32697), .A1(n42866), .B0(n14020), .C0(n14021), .Y(
        n34846) );
  OA22X1 U53307 ( .A0(net262988), .A1(n32681), .B0(n32689), .B1(n40097), .Y(
        n14020) );
  AOI222XL U53308 ( .A0(net265549), .A1(n50420), .B0(n40220), .B1(n50419),
        .C0(n40374), .C1(n50418), .Y(n14021) );
  OAI211X1 U53309 ( .A0(n32689), .A1(n42867), .B0(n13996), .C0(n13997), .Y(
        n34838) );
  OA22X1 U53310 ( .A0(net262988), .A1(n32673), .B0(n32681), .B1(n40096), .Y(
        n13996) );
  AOI222XL U53311 ( .A0(net265530), .A1(n50419), .B0(n40221), .B1(n50418),
        .C0(n40374), .C1(n50417), .Y(n13997) );
  OAI211X1 U53312 ( .A0(n32681), .A1(n42868), .B0(n13972), .C0(n13973), .Y(
        n34830) );
  OA22X1 U53313 ( .A0(net263007), .A1(n32665), .B0(n32673), .B1(n40096), .Y(
        n13972) );
  AOI222XL U53314 ( .A0(net265530), .A1(n50418), .B0(n40221), .B1(n50417),
        .C0(n40375), .C1(n50416), .Y(n13973) );
  OAI211X1 U53315 ( .A0(n32673), .A1(n42869), .B0(n13948), .C0(n13949), .Y(
        n34822) );
  OA22X1 U53316 ( .A0(net263007), .A1(n32657), .B0(n32665), .B1(n40095), .Y(
        n13948) );
  AOI222XL U53317 ( .A0(net265530), .A1(n50417), .B0(n40221), .B1(n50416),
        .C0(n40375), .C1(n50415), .Y(n13949) );
  OAI211X1 U53318 ( .A0(n32665), .A1(n42871), .B0(n13924), .C0(n13925), .Y(
        n34814) );
  OA22X1 U53319 ( .A0(net263026), .A1(n32649), .B0(n32657), .B1(n40095), .Y(
        n13924) );
  AOI222XL U53320 ( .A0(net265511), .A1(n50416), .B0(n40222), .B1(n50415),
        .C0(n40375), .C1(n50414), .Y(n13925) );
  OAI211X1 U53321 ( .A0(n32657), .A1(n42872), .B0(n13900), .C0(n13901), .Y(
        n34806) );
  OA22X1 U53322 ( .A0(net263026), .A1(n32641), .B0(n32649), .B1(n40094), .Y(
        n13900) );
  AOI222XL U53323 ( .A0(net265511), .A1(n50415), .B0(n40222), .B1(n50414),
        .C0(n40376), .C1(n50413), .Y(n13901) );
  OAI211X1 U53324 ( .A0(n32649), .A1(n42873), .B0(n13876), .C0(n13877), .Y(
        n34798) );
  OA22X1 U53325 ( .A0(net263045), .A1(n32633), .B0(n32641), .B1(n40094), .Y(
        n13876) );
  AOI222XL U53326 ( .A0(net265511), .A1(n50414), .B0(n40223), .B1(n50413),
        .C0(n40376), .C1(n50412), .Y(n13877) );
  OA22X1 U53327 ( .A0(net263045), .A1(n32625), .B0(n32633), .B1(n40093), .Y(
        n13852) );
  AOI222XL U53328 ( .A0(net265492), .A1(n50413), .B0(n40223), .B1(n50412),
        .C0(n40376), .C1(n50411), .Y(n13853) );
  OA22X1 U53329 ( .A0(net263045), .A1(n32617), .B0(n32625), .B1(n40093), .Y(
        n13828) );
  AOI222XL U53330 ( .A0(net265492), .A1(n50412), .B0(n40223), .B1(n50411),
        .C0(n40377), .C1(n50410), .Y(n13829) );
  OA22X1 U53331 ( .A0(net263406), .A1(n32609), .B0(n32617), .B1(n40073), .Y(
        n13804) );
  AOI222XL U53332 ( .A0(net265492), .A1(n50411), .B0(n40224), .B1(n50410),
        .C0(n40377), .C1(n50409), .Y(n13805) );
  OA22X1 U53333 ( .A0(net263330), .A1(n32601), .B0(n32609), .B1(n40077), .Y(
        n13780) );
  AOI222XL U53334 ( .A0(net265473), .A1(n50410), .B0(n40224), .B1(n50409),
        .C0(n40377), .C1(n50408), .Y(n13781) );
  OA22X1 U53335 ( .A0(net263349), .A1(n32593), .B0(n32601), .B1(n40076), .Y(
        n13756) );
  AOI222XL U53336 ( .A0(net265473), .A1(n50409), .B0(n40225), .B1(n50408),
        .C0(n40378), .C1(n50407), .Y(n13757) );
  OA22X1 U53337 ( .A0(net263349), .A1(n32585), .B0(n32593), .B1(n40076), .Y(
        n13732) );
  AOI222XL U53338 ( .A0(net265796), .A1(n50408), .B0(n40204), .B1(n50407),
        .C0(n40378), .C1(n50406), .Y(n13733) );
  OA22X1 U53339 ( .A0(net263368), .A1(n32577), .B0(n32585), .B1(n40075), .Y(
        n13708) );
  AOI222XL U53340 ( .A0(net265796), .A1(n50407), .B0(n40204), .B1(n50406),
        .C0(n40379), .C1(n50405), .Y(n13709) );
  OA22X1 U53341 ( .A0(net263368), .A1(n32569), .B0(n32577), .B1(n40075), .Y(
        n13684) );
  AOI222XL U53342 ( .A0(net265796), .A1(n50406), .B0(n40205), .B1(n50405),
        .C0(n40379), .C1(n50404), .Y(n13685) );
  OAI211X1 U53343 ( .A0(n32577), .A1(n42915), .B0(n13660), .C0(n13661), .Y(
        n34726) );
  OA22X1 U53344 ( .A0(net263387), .A1(n32561), .B0(n32569), .B1(n40074), .Y(
        n13660) );
  AOI222XL U53345 ( .A0(net265777), .A1(n50405), .B0(n40205), .B1(n50404),
        .C0(n40379), .C1(n50403), .Y(n13661) );
  OA22X1 U53346 ( .A0(net263387), .A1(n32553), .B0(n32561), .B1(n40074), .Y(
        n13636) );
  AOI222XL U53347 ( .A0(net265777), .A1(n50404), .B0(n40205), .B1(n50403),
        .C0(n40380), .C1(n50402), .Y(n13637) );
  OA22X1 U53348 ( .A0(net263406), .A1(n32545), .B0(n32553), .B1(n40073), .Y(
        n13612) );
  AOI222XL U53349 ( .A0(net265777), .A1(n50403), .B0(n40206), .B1(n50402),
        .C0(n40380), .C1(n50401), .Y(n13613) );
  OA22X1 U53350 ( .A0(net263406), .A1(n32537), .B0(n32545), .B1(n40073), .Y(
        n13588) );
  AOI222XL U53351 ( .A0(net265758), .A1(n50402), .B0(n40206), .B1(n50401),
        .C0(n40380), .C1(n50400), .Y(n13589) );
  OAI211X1 U53352 ( .A0(n32545), .A1(n42920), .B0(n13564), .C0(n13565), .Y(
        n34694) );
  OA22X1 U53353 ( .A0(net218368), .A1(n32529), .B0(n32537), .B1(n40072), .Y(
        n13564) );
  AOI222XL U53354 ( .A0(net265758), .A1(n50401), .B0(n40207), .B1(n50400),
        .C0(n40381), .C1(n50399), .Y(n13565) );
  OAI211X1 U53355 ( .A0(n32537), .A1(n42921), .B0(n13540), .C0(n13541), .Y(
        n34686) );
  OA22X1 U53356 ( .A0(net218336), .A1(n32521), .B0(n32529), .B1(n40072), .Y(
        n13540) );
  AOI222XL U53357 ( .A0(net265758), .A1(n50400), .B0(n40207), .B1(n50399),
        .C0(n40381), .C1(n50398), .Y(n13541) );
  OAI211X1 U53358 ( .A0(n32529), .A1(n42922), .B0(n13516), .C0(n13517), .Y(
        n34678) );
  OA22X1 U53359 ( .A0(net218350), .A1(n32513), .B0(n32521), .B1(n40071), .Y(
        n13516) );
  AOI222XL U53360 ( .A0(net265739), .A1(n50399), .B0(n40207), .B1(n50398),
        .C0(n40381), .C1(n50397), .Y(n13517) );
  OAI211X1 U53361 ( .A0(n32521), .A1(n42923), .B0(n13492), .C0(n13493), .Y(
        n34670) );
  OA22X1 U53362 ( .A0(net263444), .A1(n32505), .B0(n32513), .B1(n40071), .Y(
        n13492) );
  AOI222XL U53363 ( .A0(net265739), .A1(n50398), .B0(n40208), .B1(n50397),
        .C0(n40382), .C1(n50396), .Y(n13493) );
  OA22X1 U53364 ( .A0(net263444), .A1(n32497), .B0(n32505), .B1(n40070), .Y(
        n13468) );
  AOI222XL U53365 ( .A0(net265739), .A1(n50397), .B0(n40208), .B1(n50396),
        .C0(n40382), .C1(n50395), .Y(n13469) );
  OA22X1 U53366 ( .A0(net263463), .A1(n32489), .B0(n32497), .B1(n40070), .Y(
        n13444) );
  AOI222XL U53367 ( .A0(net265720), .A1(n50396), .B0(n40209), .B1(n50395),
        .C0(n40382), .C1(n50394), .Y(n13445) );
  OA22X1 U53368 ( .A0(net218380), .A1(n32481), .B0(n32489), .B1(n40084), .Y(
        n13420) );
  AOI222XL U53369 ( .A0(net265720), .A1(n50395), .B0(n40209), .B1(n50394),
        .C0(n40383), .C1(n50393), .Y(n13421) );
  OA22X1 U53370 ( .A0(net218392), .A1(n32473), .B0(n32481), .B1(n40084), .Y(
        n13396) );
  AOI222XL U53371 ( .A0(net265720), .A1(n50394), .B0(n40209), .B1(n50393),
        .C0(n40383), .C1(n50392), .Y(n13397) );
  OAI211X1 U53372 ( .A0(n32481), .A1(n42897), .B0(n13372), .C0(n13373), .Y(
        n34630) );
  OA22X1 U53373 ( .A0(net263216), .A1(n32465), .B0(n32473), .B1(n40083), .Y(
        n13372) );
  AOI222XL U53374 ( .A0(net265701), .A1(n50393), .B0(n40210), .B1(n50392),
        .C0(n40383), .C1(n50391), .Y(n13373) );
  OAI211X1 U53375 ( .A0(n32473), .A1(n42898), .B0(n13348), .C0(n13349), .Y(
        n34622) );
  OA22X1 U53376 ( .A0(net263216), .A1(n32457), .B0(n32465), .B1(n40083), .Y(
        n13348) );
  AOI222XL U53377 ( .A0(net265701), .A1(n50392), .B0(n40210), .B1(n50391),
        .C0(n40384), .C1(n50390), .Y(n13349) );
  OAI211X1 U53378 ( .A0(n32465), .A1(n42899), .B0(n13324), .C0(n13325), .Y(
        n34614) );
  OA22X1 U53379 ( .A0(net263235), .A1(n32449), .B0(n32457), .B1(n40082), .Y(
        n13324) );
  AOI222XL U53380 ( .A0(net265701), .A1(n50391), .B0(n40211), .B1(n50390),
        .C0(n40384), .C1(n50389), .Y(n13325) );
  OAI211X1 U53381 ( .A0(n32457), .A1(n42900), .B0(n13300), .C0(n13301), .Y(
        n34606) );
  OA22X1 U53382 ( .A0(net263235), .A1(n32441), .B0(n32449), .B1(n40082), .Y(
        n13300) );
  AOI222XL U53383 ( .A0(net265682), .A1(n50390), .B0(n40211), .B1(n50389),
        .C0(n40385), .C1(n50388), .Y(n13301) );
  OA22X1 U53384 ( .A0(net263254), .A1(n32433), .B0(n32441), .B1(n40081), .Y(
        n13276) );
  AOI222XL U53385 ( .A0(net265682), .A1(n50389), .B0(n40211), .B1(n50388),
        .C0(n40385), .C1(n50387), .Y(n13277) );
  OA22X1 U53386 ( .A0(net263254), .A1(n32425), .B0(n32433), .B1(n40081), .Y(
        n13252) );
  AOI222XL U53387 ( .A0(net265682), .A1(n50388), .B0(n40212), .B1(n50387),
        .C0(n40385), .C1(n50386), .Y(n13253) );
  OA22X1 U53388 ( .A0(net218314), .A1(n32417), .B0(n32425), .B1(n40080), .Y(
        n13228) );
  AOI222XL U53389 ( .A0(net221830), .A1(n50387), .B0(n40212), .B1(n50386),
        .C0(net217012), .C1(n50385), .Y(n13229) );
  OA22X1 U53390 ( .A0(net218312), .A1(n32409), .B0(n32417), .B1(n40080), .Y(
        n13204) );
  AOI222XL U53391 ( .A0(net221800), .A1(n50386), .B0(n40213), .B1(n50385),
        .C0(net217052), .C1(n50384), .Y(n13205) );
  OA22X1 U53392 ( .A0(net218300), .A1(n32401), .B0(n32409), .B1(n40079), .Y(
        n13180) );
  AOI222XL U53393 ( .A0(net221806), .A1(n50385), .B0(n40213), .B1(n50384),
        .C0(net217050), .C1(n50383), .Y(n13181) );
  OAI211X1 U53394 ( .A0(n32409), .A1(n42907), .B0(n13156), .C0(n13157), .Y(
        n34558) );
  AOI222XL U53395 ( .A0(net265644), .A1(n50384), .B0(n40213), .B1(n50383),
        .C0(n40381), .C1(n50382), .Y(n13157) );
  OAI211X1 U53396 ( .A0(n32401), .A1(n42908), .B0(n13132), .C0(n13133), .Y(
        n34550) );
  AOI222XL U53397 ( .A0(net265644), .A1(n50383), .B0(n40214), .B1(n50382),
        .C0(n40381), .C1(n50381), .Y(n13133) );
  OAI211X1 U53398 ( .A0(n34418), .A1(n42910), .B0(n13046), .C0(n50075), .Y(
        n34524) );
  OAI222XL U53399 ( .A0(net266654), .A1(n9658), .B0(n40159), .B1(n9657), .C0(
        n40292), .C1(n34426), .Y(n13048) );
  CLKINVX1 U53400 ( .A(n19161), .Y(n49564) );
  OAI222XL U53401 ( .A0(net266381), .A1(n9657), .B0(n40174), .B1(n34426), .C0(
        n40303), .C1(n34418), .Y(n19161) );
  AOI222XL U53402 ( .A0(net265302), .A1(n49510), .B0(n40235), .B1(n50379),
        .C0(net217108), .C1(n50378), .Y(n18224) );
  OAI211X1 U53403 ( .A0(n34090), .A1(n42828), .B0(n18199), .C0(n18200), .Y(
        n36239) );
  AOI222XL U53404 ( .A0(net265302), .A1(n50379), .B0(n40188), .B1(n50378),
        .C0(n40368), .C1(n50377), .Y(n18200) );
  OAI211X1 U53405 ( .A0(n34082), .A1(n42829), .B0(n18175), .C0(n18176), .Y(
        n36231) );
  AOI222XL U53406 ( .A0(net265283), .A1(n50378), .B0(n40198), .B1(n50377),
        .C0(n40318), .C1(n50376), .Y(n18176) );
  AOI222XL U53407 ( .A0(net265283), .A1(n50377), .B0(n40236), .B1(n50376),
        .C0(n40318), .C1(n50375), .Y(n18152) );
  AOI222XL U53408 ( .A0(net265283), .A1(n50376), .B0(n40236), .B1(n50375),
        .C0(n40319), .C1(n50374), .Y(n18128) );
  AOI222XL U53409 ( .A0(net265264), .A1(n50375), .B0(n40236), .B1(n50374),
        .C0(n40319), .C1(n50373), .Y(n18104) );
  OAI211X1 U53410 ( .A0(n34050), .A1(n42801), .B0(n18079), .C0(n18080), .Y(
        n36199) );
  AOI222XL U53411 ( .A0(net265264), .A1(n50374), .B0(n40237), .B1(n50373),
        .C0(n40319), .C1(n50372), .Y(n18080) );
  OAI211X1 U53412 ( .A0(n34042), .A1(n42803), .B0(n18055), .C0(n18056), .Y(
        n36191) );
  AOI222XL U53413 ( .A0(net265264), .A1(n50373), .B0(n40237), .B1(n50372),
        .C0(n40320), .C1(n50371), .Y(n18056) );
  OAI211X1 U53414 ( .A0(n34034), .A1(n42804), .B0(n18031), .C0(n18032), .Y(
        n36183) );
  OA22X1 U53415 ( .A0(net262931), .A1(n34018), .B0(n34026), .B1(n40100), .Y(
        n18031) );
  AOI222XL U53416 ( .A0(net265245), .A1(n50372), .B0(n40238), .B1(n50371),
        .C0(n40320), .C1(n50370), .Y(n18032) );
  OA22X1 U53417 ( .A0(net262665), .A1(n34010), .B0(n34018), .B1(n40086), .Y(
        n18007) );
  AOI222XL U53418 ( .A0(net265245), .A1(n50371), .B0(n40238), .B1(n50370),
        .C0(n40320), .C1(n50369), .Y(n18008) );
  AOI222XL U53419 ( .A0(net265245), .A1(n50370), .B0(n40238), .B1(n50369),
        .C0(n40321), .C1(n50368), .Y(n17984) );
  AOI222XL U53420 ( .A0(net265226), .A1(n50369), .B0(n40239), .B1(n50368),
        .C0(n40321), .C1(n50367), .Y(n17960) );
  OAI211X1 U53421 ( .A0(n34002), .A1(n42808), .B0(n17935), .C0(n17936), .Y(
        n36151) );
  AOI222XL U53422 ( .A0(net265226), .A1(n50368), .B0(n40239), .B1(n50367),
        .C0(n40321), .C1(n50366), .Y(n17936) );
  OA22X1 U53423 ( .A0(net262703), .A1(n33978), .B0(n33986), .B1(n40110), .Y(
        n17911) );
  AOI222XL U53424 ( .A0(net265226), .A1(n50367), .B0(n40240), .B1(n50366),
        .C0(n40322), .C1(n50365), .Y(n17912) );
  AOI222XL U53425 ( .A0(net265207), .A1(n50366), .B0(n40240), .B1(n50365),
        .C0(n40322), .C1(n50364), .Y(n17888) );
  AOI222XL U53426 ( .A0(net265207), .A1(n50365), .B0(n40240), .B1(n50364),
        .C0(n40322), .C1(n50363), .Y(n17864) );
  OAI211X1 U53427 ( .A0(n33970), .A1(n42813), .B0(n17839), .C0(n17840), .Y(
        n36119) );
  AOI222XL U53428 ( .A0(net265188), .A1(n50364), .B0(n40241), .B1(n50363),
        .C0(n40323), .C1(n50362), .Y(n17840) );
  OAI211X1 U53429 ( .A0(n33962), .A1(n42814), .B0(n17815), .C0(n17816), .Y(
        n36111) );
  AOI222XL U53430 ( .A0(net265188), .A1(n50363), .B0(n40241), .B1(n50362),
        .C0(n40323), .C1(n50361), .Y(n17816) );
  AOI222XL U53431 ( .A0(net265188), .A1(n50362), .B0(n40242), .B1(n50361),
        .C0(n40323), .C1(n50360), .Y(n17792) );
  AOI222XL U53432 ( .A0(net265169), .A1(n50361), .B0(n40242), .B1(n50360),
        .C0(n40324), .C1(n50359), .Y(n17768) );
  AOI222XL U53433 ( .A0(net265169), .A1(n50360), .B0(n40242), .B1(n50359),
        .C0(n40324), .C1(n50358), .Y(n17744) );
  AOI222XL U53434 ( .A0(net265169), .A1(n50359), .B0(n40243), .B1(n50358),
        .C0(n40325), .C1(n50357), .Y(n17720) );
  AOI222XL U53435 ( .A0(net265150), .A1(n50358), .B0(n40243), .B1(n50357),
        .C0(n40325), .C1(n50356), .Y(n17696) );
  AOI222XL U53436 ( .A0(net265150), .A1(n50357), .B0(n40244), .B1(n50356),
        .C0(n40325), .C1(n50355), .Y(n17672) );
  OAI211X1 U53437 ( .A0(n33906), .A1(n42854), .B0(n17647), .C0(n17648), .Y(
        n36055) );
  OA22X1 U53438 ( .A0(net262798), .A1(n33890), .B0(n33898), .B1(n40106), .Y(
        n17647) );
  AOI222XL U53439 ( .A0(net265150), .A1(n50356), .B0(n40244), .B1(n50355),
        .C0(n40349), .C1(n50354), .Y(n17648) );
  OAI211X1 U53440 ( .A0(n33898), .A1(n42856), .B0(n17623), .C0(n17624), .Y(
        n36047) );
  OA22X1 U53441 ( .A0(net261981), .A1(n33882), .B0(n33890), .B1(n40144), .Y(
        n17623) );
  AOI222XL U53442 ( .A0(net265131), .A1(n50355), .B0(n40244), .B1(n50354),
        .C0(n40348), .C1(n50353), .Y(n17624) );
  OAI211X1 U53443 ( .A0(n33890), .A1(n42857), .B0(n17599), .C0(n17600), .Y(
        n36039) );
  OA22X1 U53444 ( .A0(net262000), .A1(n33874), .B0(n33882), .B1(n40143), .Y(
        n17599) );
  AOI222XL U53445 ( .A0(net265131), .A1(n50354), .B0(n40245), .B1(n50353),
        .C0(n40350), .C1(n50352), .Y(n17600) );
  OAI211X1 U53446 ( .A0(n33882), .A1(n42858), .B0(n17575), .C0(n17576), .Y(
        n36031) );
  AOI222XL U53447 ( .A0(net265473), .A1(n50353), .B0(n40225), .B1(n50352),
        .C0(n40326), .C1(n50351), .Y(n17576) );
  OAI211X1 U53448 ( .A0(n33874), .A1(n42859), .B0(n17551), .C0(n17552), .Y(
        n36023) );
  AOI222XL U53449 ( .A0(net265454), .A1(n50352), .B0(n40225), .B1(n50351),
        .C0(n40326), .C1(n50350), .Y(n17552) );
  AOI222XL U53450 ( .A0(net265454), .A1(n50351), .B0(n40226), .B1(n50350),
        .C0(n40326), .C1(n50349), .Y(n17528) );
  AOI222XL U53451 ( .A0(net265454), .A1(n50350), .B0(n40226), .B1(n50349),
        .C0(n40327), .C1(n50348), .Y(n17504) );
  AOI222XL U53452 ( .A0(net265435), .A1(n50349), .B0(n40227), .B1(n50348),
        .C0(n40327), .C1(n50347), .Y(n17480) );
  AOI222XL U53453 ( .A0(net265435), .A1(n50348), .B0(n40227), .B1(n50347),
        .C0(n40327), .C1(n50346), .Y(n17456) );
  AOI222XL U53454 ( .A0(net265435), .A1(n50347), .B0(n40227), .B1(n50346),
        .C0(n40328), .C1(n50345), .Y(n17432) );
  AOI222XL U53455 ( .A0(net265416), .A1(n50346), .B0(n40228), .B1(n50345),
        .C0(n40328), .C1(n50344), .Y(n17408) );
  AOI222XL U53456 ( .A0(net265416), .A1(n50345), .B0(n40228), .B1(n50344),
        .C0(n40328), .C1(n50343), .Y(n17384) );
  AOI222XL U53457 ( .A0(net265416), .A1(n50344), .B0(n40229), .B1(n50343),
        .C0(n40329), .C1(n50342), .Y(n17360) );
  AOI222XL U53458 ( .A0(net265397), .A1(n50343), .B0(n40229), .B1(n50342),
        .C0(n40329), .C1(n50341), .Y(n17336) );
  AOI222XL U53459 ( .A0(net265397), .A1(n50342), .B0(n40229), .B1(n50341),
        .C0(n40330), .C1(n50340), .Y(n17312) );
  AOI222XL U53460 ( .A0(net265397), .A1(n50341), .B0(n40230), .B1(n50340),
        .C0(n40330), .C1(n50339), .Y(n17288) );
  AOI222XL U53461 ( .A0(net265378), .A1(n50340), .B0(n40230), .B1(n50339),
        .C0(n40330), .C1(n50338), .Y(n17264) );
  AOI222XL U53462 ( .A0(net265378), .A1(n50339), .B0(n40231), .B1(n50338),
        .C0(n40331), .C1(n50337), .Y(n17240) );
  AOI222XL U53463 ( .A0(net265378), .A1(n50338), .B0(n40231), .B1(n50337),
        .C0(n40331), .C1(n50336), .Y(n17216) );
  AOI222XL U53464 ( .A0(net265359), .A1(n50337), .B0(n40231), .B1(n50336),
        .C0(n40331), .C1(n50335), .Y(n17192) );
  OA22X1 U53465 ( .A0(net261867), .A1(n33730), .B0(n33738), .B1(n40150), .Y(
        n17167) );
  AOI222XL U53466 ( .A0(net265359), .A1(n50336), .B0(n40232), .B1(n50335),
        .C0(n40332), .C1(n50334), .Y(n17168) );
  OA22X1 U53467 ( .A0(net261886), .A1(n33722), .B0(n33730), .B1(n40150), .Y(
        n17143) );
  AOI222XL U53468 ( .A0(net265359), .A1(n50335), .B0(n40232), .B1(n50334),
        .C0(n40332), .C1(n50333), .Y(n17144) );
  OA22X1 U53469 ( .A0(net261886), .A1(n33714), .B0(n33722), .B1(n40149), .Y(
        n17119) );
  AOI222XL U53470 ( .A0(net265340), .A1(n50334), .B0(n40233), .B1(n50333),
        .C0(n40332), .C1(n50332), .Y(n17120) );
  OAI211X1 U53471 ( .A0(n33722), .A1(n42752), .B0(n17095), .C0(n17096), .Y(
        n35871) );
  AOI222XL U53472 ( .A0(net265340), .A1(n50333), .B0(n40233), .B1(n50332),
        .C0(n40333), .C1(n50331), .Y(n17096) );
  AOI222XL U53473 ( .A0(net265340), .A1(n50332), .B0(n40233), .B1(n50331),
        .C0(n40333), .C1(n50330), .Y(n17072) );
  AOI222XL U53474 ( .A0(net265321), .A1(n50331), .B0(n40234), .B1(n50330),
        .C0(n40333), .C1(n50329), .Y(n17048) );
  AOI222XL U53475 ( .A0(net265321), .A1(n50330), .B0(n40234), .B1(n50329),
        .C0(n40334), .C1(n50328), .Y(n17024) );
  AOI222XL U53476 ( .A0(net265321), .A1(n50329), .B0(n40235), .B1(n50328),
        .C0(n40334), .C1(n50327), .Y(n17000) );
  AOI222XL U53477 ( .A0(net265302), .A1(n50328), .B0(n40235), .B1(n50327),
        .C0(n40334), .C1(n50326), .Y(n16976) );
  AOI222XL U53478 ( .A0(net265302), .A1(n50327), .B0(n40230), .B1(n50326),
        .C0(n40335), .C1(n50325), .Y(n16952) );
  AOI222XL U53479 ( .A0(net264960), .A1(n50326), .B0(n40256), .B1(n50325),
        .C0(n40335), .C1(n50324), .Y(n16928) );
  AOI222XL U53480 ( .A0(net264941), .A1(n50325), .B0(n40256), .B1(n50324),
        .C0(n40336), .C1(n50323), .Y(n16904) );
  OAI211X1 U53481 ( .A0(n33650), .A1(n42762), .B0(n16879), .C0(n16880), .Y(
        n35799) );
  OA22X1 U53482 ( .A0(net261981), .A1(n33634), .B0(n33642), .B1(n40144), .Y(
        n16879) );
  AOI222XL U53483 ( .A0(net264941), .A1(n50324), .B0(n40257), .B1(n50323),
        .C0(n40336), .C1(n50322), .Y(n16880) );
  OA22X1 U53484 ( .A0(net262247), .A1(n33626), .B0(n33634), .B1(n40130), .Y(
        n16855) );
  AOI222XL U53485 ( .A0(net264941), .A1(n50323), .B0(n40257), .B1(n50322),
        .C0(n40336), .C1(n50321), .Y(n16856) );
  OAI211X1 U53486 ( .A0(n33634), .A1(n42764), .B0(n16831), .C0(n16832), .Y(
        n35783) );
  OA22X1 U53487 ( .A0(net262266), .A1(n33618), .B0(n33626), .B1(n40129), .Y(
        n16831) );
  AOI222XL U53488 ( .A0(net264922), .A1(n50322), .B0(n40258), .B1(n50321),
        .C0(n40337), .C1(n50320), .Y(n16832) );
  OAI211X1 U53489 ( .A0(n33626), .A1(n42765), .B0(n16807), .C0(n16808), .Y(
        n35775) );
  OA22X1 U53490 ( .A0(net262266), .A1(n33610), .B0(n33618), .B1(n40129), .Y(
        n16807) );
  AOI222XL U53491 ( .A0(net264922), .A1(n50321), .B0(n40258), .B1(n50320),
        .C0(n40337), .C1(n50319), .Y(n16808) );
  AOI222XL U53492 ( .A0(net264903), .A1(n50319), .B0(n40259), .B1(n50318),
        .C0(n40338), .C1(n50317), .Y(n16760) );
  AOI222XL U53493 ( .A0(net264903), .A1(n50318), .B0(n40259), .B1(n50317),
        .C0(n40338), .C1(n50316), .Y(n16736) );
  AOI222XL U53494 ( .A0(net264903), .A1(n50317), .B0(n40260), .B1(n50316),
        .C0(n40338), .C1(n50315), .Y(n16712) );
  OAI211X1 U53495 ( .A0(n33586), .A1(n42739), .B0(n16687), .C0(n16688), .Y(
        n35735) );
  OA22X1 U53496 ( .A0(net262323), .A1(n33570), .B0(n33578), .B1(n40127), .Y(
        n16687) );
  AOI222XL U53497 ( .A0(net264903), .A1(n50316), .B0(n40260), .B1(n50315),
        .C0(n40339), .C1(n50314), .Y(n16688) );
  AOI222XL U53498 ( .A0(net264884), .A1(n50315), .B0(n40260), .B1(n50314),
        .C0(n40339), .C1(n50313), .Y(n16664) );
  AOI222XL U53499 ( .A0(net264884), .A1(n50314), .B0(n40261), .B1(n50313),
        .C0(n40339), .C1(n50312), .Y(n16640) );
  AOI222XL U53500 ( .A0(net265036), .A1(n50313), .B0(n40266), .B1(n50312),
        .C0(n40340), .C1(n50311), .Y(n16616) );
  AOI222XL U53501 ( .A0(net264808), .A1(n50312), .B0(n40266), .B1(n50311),
        .C0(n40340), .C1(n50310), .Y(n16592) );
  AOI222XL U53502 ( .A0(net264808), .A1(n50311), .B0(n40265), .B1(n50310),
        .C0(n40340), .C1(n50309), .Y(n16568) );
  OA22X1 U53503 ( .A0(net262361), .A1(n33522), .B0(n33530), .B1(n40124), .Y(
        n16543) );
  AOI222XL U53504 ( .A0(net264808), .A1(n50310), .B0(n40265), .B1(n50309),
        .C0(n40341), .C1(n50308), .Y(n16544) );
  OAI211X1 U53505 ( .A0(n33530), .A1(n42747), .B0(n16519), .C0(n16520), .Y(
        n35679) );
  OA22X1 U53506 ( .A0(net262380), .A1(n33514), .B0(n33522), .B1(n40124), .Y(
        n16519) );
  AOI222XL U53507 ( .A0(net264827), .A1(n50309), .B0(n40265), .B1(n50308),
        .C0(n40341), .C1(n50307), .Y(n16520) );
  OAI211X1 U53508 ( .A0(n33522), .A1(n42748), .B0(n16495), .C0(n16496), .Y(
        n35671) );
  AOI222XL U53509 ( .A0(net264827), .A1(n50308), .B0(n40264), .B1(n50307),
        .C0(n40342), .C1(n50306), .Y(n16496) );
  OAI211X1 U53510 ( .A0(n33514), .A1(n42749), .B0(n16471), .C0(n16472), .Y(
        n35663) );
  AOI222XL U53511 ( .A0(net264827), .A1(n50307), .B0(n40266), .B1(n50306),
        .C0(n40342), .C1(n50305), .Y(n16472) );
  OAI211X1 U53512 ( .A0(n33506), .A1(n42783), .B0(n16447), .C0(n16448), .Y(
        n35655) );
  AOI222XL U53513 ( .A0(net264846), .A1(n50306), .B0(n40263), .B1(n50305),
        .C0(n40342), .C1(n50304), .Y(n16448) );
  AOI222XL U53514 ( .A0(net264846), .A1(n50305), .B0(n40263), .B1(n50304),
        .C0(n40343), .C1(n50303), .Y(n16424) );
  AOI222XL U53515 ( .A0(net264846), .A1(n50304), .B0(n40263), .B1(n50303),
        .C0(n40343), .C1(n50302), .Y(n16400) );
  AOI222XL U53516 ( .A0(net264865), .A1(n50303), .B0(n40262), .B1(n50302),
        .C0(n40343), .C1(n50301), .Y(n16376) );
  AOI222XL U53517 ( .A0(net264865), .A1(n50302), .B0(n40262), .B1(n50301),
        .C0(n40344), .C1(n50300), .Y(n16352) );
  AOI222XL U53518 ( .A0(net264865), .A1(n50301), .B0(n40261), .B1(n50300),
        .C0(n40344), .C1(n50299), .Y(n16328) );
  OAI211X1 U53519 ( .A0(n33458), .A1(n42790), .B0(n16303), .C0(n16304), .Y(
        n35607) );
  OA22X1 U53520 ( .A0(net262190), .A1(n33442), .B0(n33450), .B1(n40134), .Y(
        n16303) );
  AOI222XL U53521 ( .A0(net265131), .A1(n50300), .B0(n40245), .B1(n50299),
        .C0(n40344), .C1(n50298), .Y(n16304) );
  OA22X1 U53522 ( .A0(net262190), .A1(n33434), .B0(n33442), .B1(n40134), .Y(
        n16279) );
  AOI222XL U53523 ( .A0(net265131), .A1(n50299), .B0(n40246), .B1(n50298),
        .C0(n40345), .C1(n50297), .Y(n16280) );
  OAI211X1 U53524 ( .A0(n33442), .A1(n42792), .B0(n16255), .C0(n16256), .Y(
        n35591) );
  AOI222XL U53525 ( .A0(net265112), .A1(n50298), .B0(n40246), .B1(n50297),
        .C0(n40345), .C1(n50296), .Y(n16256) );
  OAI211X1 U53526 ( .A0(n33434), .A1(n42793), .B0(n16231), .C0(n16232), .Y(
        n35583) );
  AOI222XL U53527 ( .A0(net265112), .A1(n50297), .B0(n40246), .B1(n50296),
        .C0(n40345), .C1(n50295), .Y(n16232) );
  OAI211X1 U53528 ( .A0(n33426), .A1(n42794), .B0(n16207), .C0(n16208), .Y(
        n35575) );
  AOI222XL U53529 ( .A0(net265112), .A1(n50296), .B0(n40247), .B1(n50295),
        .C0(n40346), .C1(n50294), .Y(n16208) );
  OA22X1 U53530 ( .A0(net262228), .A1(n33402), .B0(n33410), .B1(n40132), .Y(
        n16183) );
  AOI222XL U53531 ( .A0(net221812), .A1(n50295), .B0(n40247), .B1(n50294),
        .C0(n40346), .C1(n50293), .Y(n16184) );
  OA22X1 U53532 ( .A0(net262228), .A1(n33394), .B0(n33402), .B1(n40131), .Y(
        n16159) );
  AOI222XL U53533 ( .A0(net221802), .A1(n50294), .B0(n40248), .B1(n50293),
        .C0(n40346), .C1(n50292), .Y(n16160) );
  OAI211X1 U53534 ( .A0(n33402), .A1(n42798), .B0(n16135), .C0(n16136), .Y(
        n35551) );
  AOI222XL U53535 ( .A0(net221820), .A1(n50293), .B0(n40248), .B1(n50292),
        .C0(n40347), .C1(n50291), .Y(n16136) );
  OAI211X1 U53536 ( .A0(n33394), .A1(n42767), .B0(n16111), .C0(n16112), .Y(
        n35543) );
  AOI222XL U53537 ( .A0(net265074), .A1(n50292), .B0(n40248), .B1(n50291),
        .C0(n40347), .C1(n50290), .Y(n16112) );
  AOI222XL U53538 ( .A0(net265074), .A1(n50291), .B0(n40249), .B1(n50290),
        .C0(n40348), .C1(n50289), .Y(n16088) );
  OA22X1 U53539 ( .A0(net263615), .A1(n33362), .B0(n33370), .B1(n40060), .Y(
        n16063) );
  AOI222XL U53540 ( .A0(net265074), .A1(n50290), .B0(n40249), .B1(n50289),
        .C0(n40348), .C1(n50288), .Y(n16064) );
  OAI211X1 U53541 ( .A0(n33370), .A1(n42770), .B0(n16039), .C0(n16040), .Y(
        n35519) );
  OA22X1 U53542 ( .A0(net263615), .A1(n33354), .B0(n33362), .B1(n40060), .Y(
        n16039) );
  AOI222XL U53543 ( .A0(net265055), .A1(n50289), .B0(n40250), .B1(n50288),
        .C0(n40348), .C1(n50287), .Y(n16040) );
  OAI211X1 U53544 ( .A0(n33362), .A1(n42771), .B0(n16015), .C0(n16016), .Y(
        n35511) );
  AOI222XL U53545 ( .A0(net265055), .A1(n50288), .B0(n40250), .B1(n50287),
        .C0(n40349), .C1(n50286), .Y(n16016) );
  OAI211X1 U53546 ( .A0(n33354), .A1(n42772), .B0(n15991), .C0(n15992), .Y(
        n35503) );
  AOI222XL U53547 ( .A0(net265055), .A1(n50287), .B0(n40250), .B1(n50286),
        .C0(n40349), .C1(n50285), .Y(n15992) );
  OAI211X1 U53548 ( .A0(n33346), .A1(n42773), .B0(n15967), .C0(n15968), .Y(
        n35495) );
  OA22X1 U53549 ( .A0(net263653), .A1(n33330), .B0(n33338), .B1(n40058), .Y(
        n15967) );
  AOI222XL U53550 ( .A0(net265036), .A1(n50286), .B0(n40251), .B1(n50285),
        .C0(n40349), .C1(n50284), .Y(n15968) );
  OA22X1 U53551 ( .A0(net263653), .A1(n33322), .B0(n33330), .B1(n40058), .Y(
        n15943) );
  AOI222XL U53552 ( .A0(net265036), .A1(n50285), .B0(n40251), .B1(n50284),
        .C0(n40382), .C1(n50283), .Y(n15944) );
  OAI211X1 U53553 ( .A0(n33330), .A1(n42776), .B0(n15919), .C0(n15920), .Y(
        n35479) );
  AOI222XL U53554 ( .A0(net265036), .A1(n50284), .B0(n40252), .B1(n50283),
        .C0(net216968), .C1(n50282), .Y(n15920) );
  AOI222XL U53555 ( .A0(net265017), .A1(n50283), .B0(n40252), .B1(n50282),
        .C0(n40382), .C1(n50281), .Y(n15896) );
  AOI222XL U53556 ( .A0(net265017), .A1(n50282), .B0(n40252), .B1(n50281),
        .C0(n40350), .C1(n50280), .Y(n15872) );
  OA22X1 U53557 ( .A0(net263691), .A1(n33290), .B0(n33298), .B1(n40057), .Y(
        n15847) );
  AOI222XL U53558 ( .A0(net265017), .A1(n50281), .B0(n40253), .B1(n50280),
        .C0(n40350), .C1(n50279), .Y(n15848) );
  OAI211X1 U53559 ( .A0(n33298), .A1(n42780), .B0(n15823), .C0(n15824), .Y(
        n35447) );
  AOI222XL U53560 ( .A0(net264998), .A1(n50280), .B0(n40253), .B1(n50279),
        .C0(n40350), .C1(n50278), .Y(n15824) );
  OAI211X1 U53561 ( .A0(n33290), .A1(n42782), .B0(n15799), .C0(n15800), .Y(
        n35439) );
  AOI222XL U53562 ( .A0(net264998), .A1(n50279), .B0(n40254), .B1(n50278),
        .C0(n40341), .C1(n50277), .Y(n15800) );
  OAI211X1 U53563 ( .A0(n33282), .A1(n42960), .B0(n15775), .C0(n15776), .Y(
        n35431) );
  AOI222XL U53564 ( .A0(net264998), .A1(n50278), .B0(n40254), .B1(n50277),
        .C0(n40345), .C1(n50276), .Y(n15776) );
  OA22X1 U53565 ( .A0(net218418), .A1(n33258), .B0(n33266), .B1(n40055), .Y(
        n15751) );
  AOI222XL U53566 ( .A0(net264979), .A1(n50277), .B0(n40254), .B1(n50276),
        .C0(net217036), .C1(n50275), .Y(n15752) );
  OAI211X1 U53567 ( .A0(n33266), .A1(n42946), .B0(n15727), .C0(n15728), .Y(
        n35415) );
  OA22X1 U53568 ( .A0(net263558), .A1(n33250), .B0(n33258), .B1(n40054), .Y(
        n15727) );
  AOI222XL U53569 ( .A0(net264979), .A1(n50276), .B0(n40255), .B1(n50275),
        .C0(n40351), .C1(n50274), .Y(n15728) );
  OAI211X1 U53570 ( .A0(n33258), .A1(n42947), .B0(n15703), .C0(n15704), .Y(
        n35407) );
  OA22X1 U53571 ( .A0(net263463), .A1(n33242), .B0(n33250), .B1(n40069), .Y(
        n15703) );
  AOI222XL U53572 ( .A0(net264979), .A1(n50275), .B0(n40255), .B1(n50274),
        .C0(n40351), .C1(n50273), .Y(n15704) );
  OAI211X1 U53573 ( .A0(n33250), .A1(n42948), .B0(n15679), .C0(n15680), .Y(
        n35399) );
  AOI222XL U53574 ( .A0(net264960), .A1(n50274), .B0(n40256), .B1(n50273),
        .C0(n40352), .C1(n50272), .Y(n15680) );
  AOI222XL U53575 ( .A0(net265967), .A1(n50273), .B0(n40193), .B1(n50272),
        .C0(n40352), .C1(n50271), .Y(n15656) );
  OA22X1 U53576 ( .A0(net263501), .A1(n33218), .B0(n33226), .B1(n40067), .Y(
        n15631) );
  AOI222XL U53577 ( .A0(net265967), .A1(n50272), .B0(n40193), .B1(n50271),
        .C0(n40352), .C1(n50270), .Y(n15632) );
  OA22X1 U53578 ( .A0(net263501), .A1(n33210), .B0(n33218), .B1(n40067), .Y(
        n15607) );
  AOI222XL U53579 ( .A0(net265967), .A1(n50271), .B0(n40194), .B1(n50270),
        .C0(n40353), .C1(n50269), .Y(n15608) );
  OAI211X1 U53580 ( .A0(n33218), .A1(n42953), .B0(n15583), .C0(n15584), .Y(
        n35367) );
  OA22X1 U53581 ( .A0(net218322), .A1(n33202), .B0(n33210), .B1(n40066), .Y(
        n15583) );
  AOI222XL U53582 ( .A0(net265948), .A1(n50270), .B0(n40194), .B1(n50269),
        .C0(n40353), .C1(n50268), .Y(n15584) );
  OAI211X1 U53583 ( .A0(n33210), .A1(n42954), .B0(n15559), .C0(n15560), .Y(
        n35359) );
  OA22X1 U53584 ( .A0(net218398), .A1(n33194), .B0(n33202), .B1(n40066), .Y(
        n15559) );
  AOI222XL U53585 ( .A0(net265948), .A1(n50269), .B0(n40195), .B1(n50268),
        .C0(n40353), .C1(n50267), .Y(n15560) );
  OAI211X1 U53586 ( .A0(n33202), .A1(n42955), .B0(n15535), .C0(n15536), .Y(
        n35351) );
  AOI222XL U53587 ( .A0(net265948), .A1(n50268), .B0(n40195), .B1(n50267),
        .C0(n40354), .C1(n50266), .Y(n15536) );
  AOI222XL U53588 ( .A0(net265929), .A1(n50267), .B0(n40195), .B1(n50266),
        .C0(n40354), .C1(n50265), .Y(n15512) );
  OA22X1 U53589 ( .A0(net263558), .A1(n33170), .B0(n33178), .B1(n40064), .Y(
        n15487) );
  AOI222XL U53590 ( .A0(net265929), .A1(n50266), .B0(n40196), .B1(n50265),
        .C0(n40354), .C1(n50264), .Y(n15488) );
  OA22X1 U53591 ( .A0(net263558), .A1(n33162), .B0(n33170), .B1(n40064), .Y(
        n15463) );
  AOI222XL U53592 ( .A0(net265929), .A1(n50265), .B0(n40196), .B1(n50264),
        .C0(n40355), .C1(n50263), .Y(n15464) );
  OAI211X1 U53593 ( .A0(n33170), .A1(n42960), .B0(n15439), .C0(n15440), .Y(
        n35319) );
  OA22X1 U53594 ( .A0(net263558), .A1(n33154), .B0(n33162), .B1(n40063), .Y(
        n15439) );
  AOI222XL U53595 ( .A0(net265910), .A1(n50264), .B0(n40197), .B1(n50263),
        .C0(n40355), .C1(n50262), .Y(n15440) );
  OAI211X1 U53596 ( .A0(n33162), .A1(n42928), .B0(n15415), .C0(n15416), .Y(
        n35311) );
  OA22X1 U53597 ( .A0(net263577), .A1(n33146), .B0(n33154), .B1(n40063), .Y(
        n15415) );
  AOI222XL U53598 ( .A0(net265910), .A1(n50263), .B0(n40197), .B1(n50262),
        .C0(n40355), .C1(n50261), .Y(n15416) );
  OAI211X1 U53599 ( .A0(n33154), .A1(n42930), .B0(n15391), .C0(n15392), .Y(
        n35303) );
  OA22X1 U53600 ( .A0(net263577), .A1(n33138), .B0(n33146), .B1(n40062), .Y(
        n15391) );
  AOI222XL U53601 ( .A0(net265910), .A1(n50262), .B0(n40197), .B1(n50261),
        .C0(n40356), .C1(n50260), .Y(n15392) );
  OA22X1 U53602 ( .A0(net263596), .A1(n33130), .B0(n33138), .B1(n40062), .Y(
        n15367) );
  AOI222XL U53603 ( .A0(net265891), .A1(n50261), .B0(n40198), .B1(n50260),
        .C0(n40356), .C1(n50259), .Y(n15368) );
  OA22X1 U53604 ( .A0(net263596), .A1(n33122), .B0(n33130), .B1(n40061), .Y(
        n15343) );
  AOI222XL U53605 ( .A0(net265891), .A1(n50260), .B0(n40198), .B1(n50259),
        .C0(n40356), .C1(n50258), .Y(n15344) );
  OAI211X1 U53606 ( .A0(n33130), .A1(n42933), .B0(n15319), .C0(n15320), .Y(
        n35279) );
  AOI222XL U53607 ( .A0(net265891), .A1(n50259), .B0(n40199), .B1(n50258),
        .C0(n40357), .C1(n50257), .Y(n15320) );
  AOI222XL U53608 ( .A0(net265872), .A1(n50258), .B0(n40199), .B1(n50257),
        .C0(n40357), .C1(n50256), .Y(n15296) );
  AOI222XL U53609 ( .A0(net265872), .A1(n50257), .B0(n40199), .B1(n50256),
        .C0(n40358), .C1(n50255), .Y(n15272) );
  AOI222XL U53610 ( .A0(net265872), .A1(n50256), .B0(n40200), .B1(n50255),
        .C0(n40358), .C1(n50254), .Y(n15248) );
  OAI211X1 U53611 ( .A0(n33098), .A1(n42938), .B0(n15223), .C0(n15224), .Y(
        n35247) );
  OA22X1 U53612 ( .A0(net263919), .A1(n33082), .B0(n33090), .B1(n40044), .Y(
        n15223) );
  AOI222XL U53613 ( .A0(net265853), .A1(n50255), .B0(n40200), .B1(n50254),
        .C0(n40358), .C1(n50253), .Y(n15224) );
  OAI211X1 U53614 ( .A0(n33090), .A1(n42939), .B0(n15199), .C0(n15200), .Y(
        n35239) );
  OA22X1 U53615 ( .A0(net263919), .A1(n33074), .B0(n33082), .B1(n40043), .Y(
        n15199) );
  AOI222XL U53616 ( .A0(net265853), .A1(n50254), .B0(n40201), .B1(n50253),
        .C0(n40359), .C1(n50252), .Y(n15200) );
  OAI211X1 U53617 ( .A0(n33082), .A1(n42940), .B0(n15175), .C0(n15176), .Y(
        n35231) );
  OA22X1 U53618 ( .A0(net263919), .A1(n33066), .B0(n33074), .B1(n40043), .Y(
        n15175) );
  AOI222XL U53619 ( .A0(net265853), .A1(n50253), .B0(n40201), .B1(n50252),
        .C0(n40359), .C1(n50251), .Y(n15176) );
  OAI211X1 U53620 ( .A0(n33074), .A1(n42941), .B0(n15151), .C0(n15152), .Y(
        n35223) );
  AOI222XL U53621 ( .A0(net265834), .A1(n50252), .B0(n40201), .B1(n50251),
        .C0(n40359), .C1(n50250), .Y(n15152) );
  AOI222XL U53622 ( .A0(net265834), .A1(n50251), .B0(n40202), .B1(n50250),
        .C0(n40360), .C1(n50249), .Y(n15128) );
  AOI222XL U53623 ( .A0(net265834), .A1(n50250), .B0(n40202), .B1(n50249),
        .C0(n40360), .C1(n50248), .Y(n15104) );
  OA22X1 U53624 ( .A0(net263957), .A1(n33034), .B0(n33042), .B1(n40042), .Y(
        n15079) );
  AOI222XL U53625 ( .A0(net265815), .A1(n50249), .B0(n40203), .B1(n50248),
        .C0(n40360), .C1(n50247), .Y(n15080) );
  OAI211X1 U53626 ( .A0(n33042), .A1(n42978), .B0(n15055), .C0(n15056), .Y(
        n35191) );
  OA22X1 U53627 ( .A0(net263976), .A1(n33026), .B0(n33034), .B1(n40041), .Y(
        n15055) );
  AOI222XL U53628 ( .A0(net265815), .A1(n50248), .B0(n40203), .B1(n50247),
        .C0(n40347), .C1(n50246), .Y(n15056) );
  OAI211X1 U53629 ( .A0(n33034), .A1(n42979), .B0(n15031), .C0(n15032), .Y(
        n35183) );
  OA22X1 U53630 ( .A0(net263976), .A1(n33018), .B0(n33026), .B1(n40041), .Y(
        n15031) );
  AOI222XL U53631 ( .A0(net265815), .A1(n50247), .B0(n40198), .B1(n50246),
        .C0(n40351), .C1(n50245), .Y(n15032) );
  OAI211X1 U53632 ( .A0(n33026), .A1(n42980), .B0(n15007), .C0(n15008), .Y(
        n35175) );
  OA22X1 U53633 ( .A0(net263995), .A1(n33010), .B0(n33018), .B1(n40040), .Y(
        n15007) );
  AOI222XL U53634 ( .A0(net221892), .A1(n50246), .B0(net217934), .B1(n50245),
        .C0(n40377), .C1(n50244), .Y(n15008) );
  OAI211X1 U53635 ( .A0(n33018), .A1(n42981), .B0(n14983), .C0(n14984), .Y(
        n35167) );
  OA22X1 U53636 ( .A0(net263995), .A1(n33002), .B0(n33010), .B1(n40040), .Y(
        n14983) );
  AOI222XL U53637 ( .A0(net221892), .A1(n50245), .B0(n40184), .B1(n50244),
        .C0(n40361), .C1(n50243), .Y(n14984) );
  AOI222XL U53638 ( .A0(net266119), .A1(n50244), .B0(n40184), .B1(n50243),
        .C0(n40361), .C1(n50242), .Y(n14960) );
  AOI222XL U53639 ( .A0(net266119), .A1(n50243), .B0(n40185), .B1(n50242),
        .C0(n40361), .C1(n50241), .Y(n14936) );
  AOI222XL U53640 ( .A0(net266119), .A1(n50242), .B0(n40185), .B1(n50241),
        .C0(n40362), .C1(n50240), .Y(n14912) );
  AOI222XL U53641 ( .A0(net266100), .A1(n50241), .B0(n40185), .B1(n50240),
        .C0(n40362), .C1(n50239), .Y(n14888) );
  OA22X1 U53642 ( .A0(net263767), .A1(n32962), .B0(n32970), .B1(n40052), .Y(
        n14863) );
  AOI222XL U53643 ( .A0(net266100), .A1(n50240), .B0(n40195), .B1(n50239),
        .C0(n40363), .C1(n50238), .Y(n14864) );
  OAI211X1 U53644 ( .A0(n32970), .A1(n42988), .B0(n14839), .C0(n14840), .Y(
        n35119) );
  OA22X1 U53645 ( .A0(net262646), .A1(n32954), .B0(n32962), .B1(n40052), .Y(
        n14839) );
  AOI222XL U53646 ( .A0(net266100), .A1(n50239), .B0(n40194), .B1(n50238),
        .C0(n40363), .C1(n50237), .Y(n14840) );
  OAI211X1 U53647 ( .A0(n32962), .A1(n42990), .B0(n14815), .C0(n14816), .Y(
        n35111) );
  OA22X1 U53648 ( .A0(net263558), .A1(n32946), .B0(n32954), .B1(n40051), .Y(
        n14815) );
  AOI222XL U53649 ( .A0(net266081), .A1(n50238), .B0(n40186), .B1(n50237),
        .C0(n40363), .C1(n50236), .Y(n14816) );
  OAI211X1 U53650 ( .A0(n32954), .A1(n42827), .B0(n14791), .C0(n14792), .Y(
        n35103) );
  AOI222XL U53651 ( .A0(net266081), .A1(n50237), .B0(n40186), .B1(n50236),
        .C0(n40366), .C1(n50235), .Y(n14792) );
  AOI222XL U53652 ( .A0(net266062), .A1(n50235), .B0(n40187), .B1(n50234),
        .C0(net216994), .C1(n50233), .Y(n14744) );
  AOI222XL U53653 ( .A0(net266062), .A1(n50234), .B0(n40187), .B1(n50233),
        .C0(n40364), .C1(n50232), .Y(n14720) );
  OAI211X1 U53654 ( .A0(n32922), .A1(n42963), .B0(n14695), .C0(n14696), .Y(
        n35071) );
  AOI222XL U53655 ( .A0(net266062), .A1(n50233), .B0(n40188), .B1(n50232),
        .C0(n40364), .C1(n50231), .Y(n14696) );
  OAI211X1 U53656 ( .A0(n32914), .A1(n42964), .B0(n14671), .C0(n14672), .Y(
        n35063) );
  OA22X1 U53657 ( .A0(net263843), .A1(n32898), .B0(n32906), .B1(n40048), .Y(
        n14671) );
  AOI222XL U53658 ( .A0(net266043), .A1(n50232), .B0(n40188), .B1(n50231),
        .C0(n40364), .C1(n50230), .Y(n14672) );
  OAI211X1 U53659 ( .A0(n32906), .A1(n42965), .B0(n14647), .C0(n14648), .Y(
        n35055) );
  OA22X1 U53660 ( .A0(net263843), .A1(n32890), .B0(n32898), .B1(n40048), .Y(
        n14647) );
  AOI222XL U53661 ( .A0(net266043), .A1(n50231), .B0(n40188), .B1(n50230),
        .C0(n40365), .C1(n50229), .Y(n14648) );
  OAI211X1 U53662 ( .A0(n32898), .A1(n42966), .B0(n14623), .C0(n14624), .Y(
        n35047) );
  OA22X1 U53663 ( .A0(net263862), .A1(n32882), .B0(n32890), .B1(n40047), .Y(
        n14623) );
  AOI222XL U53664 ( .A0(net266043), .A1(n50230), .B0(n40189), .B1(n50229),
        .C0(n40365), .C1(n50228), .Y(n14624) );
  OAI211X1 U53665 ( .A0(n32890), .A1(n42967), .B0(n14599), .C0(n14600), .Y(
        n35039) );
  OA22X1 U53666 ( .A0(net263862), .A1(n32874), .B0(n32882), .B1(n40047), .Y(
        n14599) );
  AOI222XL U53667 ( .A0(net266024), .A1(n50229), .B0(n40189), .B1(n50228),
        .C0(n40365), .C1(n50227), .Y(n14600) );
  OAI211X1 U53668 ( .A0(n32882), .A1(n42969), .B0(n14575), .C0(n14576), .Y(
        n35031) );
  OA22X1 U53669 ( .A0(net263862), .A1(n32866), .B0(n32874), .B1(n40046), .Y(
        n14575) );
  AOI222XL U53670 ( .A0(net266024), .A1(n50228), .B0(n40190), .B1(n50227),
        .C0(n40366), .C1(n50226), .Y(n14576) );
  AOI222XL U53671 ( .A0(net266024), .A1(n50227), .B0(n40190), .B1(n50226),
        .C0(n40366), .C1(n50225), .Y(n14552) );
  AOI222XL U53672 ( .A0(net266005), .A1(n50226), .B0(n40190), .B1(n50225),
        .C0(n40366), .C1(n50224), .Y(n14528) );
  AOI222XL U53673 ( .A0(net266005), .A1(n50225), .B0(n40191), .B1(n50224),
        .C0(n40367), .C1(n50223), .Y(n14504) );
  AOI222XL U53674 ( .A0(net266005), .A1(n50224), .B0(n40191), .B1(n50223),
        .C0(n40367), .C1(n50222), .Y(n14480) );
  OAI211X1 U53675 ( .A0(n32842), .A1(n42974), .B0(n14455), .C0(n14456), .Y(
        n34991) );
  AOI222XL U53676 ( .A0(net221848), .A1(n50223), .B0(n40192), .B1(n50222),
        .C0(n40368), .C1(n50221), .Y(n14456) );
  OAI211X1 U53677 ( .A0(n32834), .A1(n42976), .B0(n14431), .C0(n14432), .Y(
        n34983) );
  OA22X1 U53678 ( .A0(net263102), .A1(n32818), .B0(n32826), .B1(n40089), .Y(
        n14431) );
  AOI222XL U53679 ( .A0(net221824), .A1(n50222), .B0(n40192), .B1(n50221),
        .C0(n40368), .C1(n50220), .Y(n14432) );
  OAI211X1 U53680 ( .A0(n32826), .A1(n42880), .B0(n14407), .C0(n14408), .Y(
        n34975) );
  OA22X1 U53681 ( .A0(net263121), .A1(n32810), .B0(n32818), .B1(n40089), .Y(
        n14407) );
  AOI222XL U53682 ( .A0(net221846), .A1(n50221), .B0(n40192), .B1(n50220),
        .C0(n40368), .C1(n50219), .Y(n14408) );
  OAI211X1 U53683 ( .A0(n32818), .A1(n42881), .B0(n14383), .C0(n14384), .Y(
        n34967) );
  OA22X1 U53684 ( .A0(net263121), .A1(n32802), .B0(n32810), .B1(n40088), .Y(
        n14383) );
  AOI222XL U53685 ( .A0(net265644), .A1(n50220), .B0(n40214), .B1(n50219),
        .C0(n40369), .C1(n50218), .Y(n14384) );
  OAI211X1 U53686 ( .A0(n32810), .A1(n42882), .B0(n14359), .C0(n14360), .Y(
        n34959) );
  OA22X1 U53687 ( .A0(net263140), .A1(n32794), .B0(n32802), .B1(n40088), .Y(
        n14359) );
  AOI222XL U53688 ( .A0(net265625), .A1(n50219), .B0(n40215), .B1(n50218),
        .C0(n40369), .C1(n50217), .Y(n14360) );
  OAI211X1 U53689 ( .A0(n32802), .A1(n42883), .B0(n14335), .C0(n14336), .Y(
        n34951) );
  OA22X1 U53690 ( .A0(net263140), .A1(n32786), .B0(n32794), .B1(n40087), .Y(
        n14335) );
  AOI222XL U53691 ( .A0(net265625), .A1(n50218), .B0(n40215), .B1(n50217),
        .C0(n40369), .C1(n50216), .Y(n14336) );
  OA22X1 U53692 ( .A0(net263159), .A1(n32778), .B0(n32786), .B1(n40087), .Y(
        n14311) );
  AOI222XL U53693 ( .A0(net265625), .A1(n50217), .B0(n40215), .B1(n50216),
        .C0(n40370), .C1(n50215), .Y(n14312) );
  OA22X1 U53694 ( .A0(net263159), .A1(n32770), .B0(n32778), .B1(n40086), .Y(
        n14287) );
  AOI222XL U53695 ( .A0(net265606), .A1(n50216), .B0(n40216), .B1(n50215),
        .C0(n40370), .C1(n50214), .Y(n14288) );
  AOI222XL U53696 ( .A0(net265606), .A1(n50215), .B0(n40216), .B1(n50214),
        .C0(n40370), .C1(n50213), .Y(n14264) );
  AOI222XL U53697 ( .A0(net265606), .A1(n50214), .B0(n40217), .B1(n50213),
        .C0(n40371), .C1(n50212), .Y(n14240) );
  OA22X1 U53698 ( .A0(net263178), .A1(n32746), .B0(n32754), .B1(n40085), .Y(
        n14215) );
  AOI222XL U53699 ( .A0(net265587), .A1(n50213), .B0(n40217), .B1(n50212),
        .C0(n40371), .C1(n50211), .Y(n14216) );
  OA22X1 U53700 ( .A0(net218432), .A1(n32738), .B0(n32746), .B1(n40084), .Y(
        n14191) );
  AOI222XL U53701 ( .A0(net265587), .A1(n50212), .B0(n40217), .B1(n50211),
        .C0(n40371), .C1(n50210), .Y(n14192) );
  OAI211X1 U53702 ( .A0(n32746), .A1(n42891), .B0(n14167), .C0(n14168), .Y(
        n34895) );
  OA22X1 U53703 ( .A0(net262931), .A1(n32730), .B0(n32738), .B1(n40100), .Y(
        n14167) );
  AOI222XL U53704 ( .A0(net265587), .A1(n50211), .B0(n40218), .B1(n50210),
        .C0(n40372), .C1(n50209), .Y(n14168) );
  OAI211X1 U53705 ( .A0(n32738), .A1(n42892), .B0(n14143), .C0(n14144), .Y(
        n34887) );
  OA22X1 U53706 ( .A0(net262950), .A1(n32722), .B0(n32730), .B1(n40099), .Y(
        n14143) );
  AOI222XL U53707 ( .A0(net265568), .A1(n50210), .B0(n40218), .B1(n50209),
        .C0(n40372), .C1(n50208), .Y(n14144) );
  OAI211X1 U53708 ( .A0(n32730), .A1(n42893), .B0(n14119), .C0(n14120), .Y(
        n34879) );
  AOI222XL U53709 ( .A0(net265568), .A1(n50209), .B0(n40219), .B1(n50208),
        .C0(n40372), .C1(n50207), .Y(n14120) );
  AOI222XL U53710 ( .A0(net265568), .A1(n50208), .B0(n40219), .B1(n50207),
        .C0(n40373), .C1(n50206), .Y(n14096) );
  AOI222XL U53711 ( .A0(net265549), .A1(n50207), .B0(n40219), .B1(n50206),
        .C0(n40373), .C1(n50205), .Y(n14072) );
  AOI222XL U53712 ( .A0(net265549), .A1(n50206), .B0(n40220), .B1(n50205),
        .C0(n40374), .C1(n50204), .Y(n14048) );
  OAI211X1 U53713 ( .A0(n32698), .A1(n42866), .B0(n14023), .C0(n14024), .Y(
        n34847) );
  OA22X1 U53714 ( .A0(net262988), .A1(n32682), .B0(n32690), .B1(n40097), .Y(
        n14023) );
  AOI222XL U53715 ( .A0(net265549), .A1(n50205), .B0(n40220), .B1(n50204),
        .C0(n40374), .C1(n50203), .Y(n14024) );
  OAI211X1 U53716 ( .A0(n32690), .A1(n42867), .B0(n13999), .C0(n14000), .Y(
        n34839) );
  OA22X1 U53717 ( .A0(net262988), .A1(n32674), .B0(n32682), .B1(n40096), .Y(
        n13999) );
  AOI222XL U53718 ( .A0(net265530), .A1(n50204), .B0(n40221), .B1(n50203),
        .C0(n40374), .C1(n50202), .Y(n14000) );
  OAI211X1 U53719 ( .A0(n32682), .A1(n42868), .B0(n13975), .C0(n13976), .Y(
        n34831) );
  OA22X1 U53720 ( .A0(net263007), .A1(n32666), .B0(n32674), .B1(n40096), .Y(
        n13975) );
  AOI222XL U53721 ( .A0(net265530), .A1(n50203), .B0(n40221), .B1(n50202),
        .C0(n40375), .C1(n50201), .Y(n13976) );
  OAI211X1 U53722 ( .A0(n32674), .A1(n42869), .B0(n13951), .C0(n13952), .Y(
        n34823) );
  OA22X1 U53723 ( .A0(net263007), .A1(n32658), .B0(n32666), .B1(n40095), .Y(
        n13951) );
  AOI222XL U53724 ( .A0(net265530), .A1(n50202), .B0(n40221), .B1(n50201),
        .C0(n40375), .C1(n50200), .Y(n13952) );
  OAI211X1 U53725 ( .A0(n32666), .A1(n42870), .B0(n13927), .C0(n13928), .Y(
        n34815) );
  OA22X1 U53726 ( .A0(net263026), .A1(n32650), .B0(n32658), .B1(n40095), .Y(
        n13927) );
  AOI222XL U53727 ( .A0(net265511), .A1(n50201), .B0(n40222), .B1(n50200),
        .C0(n40375), .C1(n50199), .Y(n13928) );
  AOI222XL U53728 ( .A0(net265511), .A1(n50200), .B0(n40222), .B1(n50199),
        .C0(n40376), .C1(n50198), .Y(n13904) );
  AOI222XL U53729 ( .A0(net265511), .A1(n50199), .B0(n40223), .B1(n50198),
        .C0(n40376), .C1(n50197), .Y(n13880) );
  AOI222XL U53730 ( .A0(net265492), .A1(n50198), .B0(n40223), .B1(n50197),
        .C0(n40376), .C1(n50196), .Y(n13856) );
  AOI222XL U53731 ( .A0(net265492), .A1(n50197), .B0(n40223), .B1(n50196),
        .C0(n40377), .C1(n50195), .Y(n13832) );
  OAI211X1 U53732 ( .A0(n32626), .A1(n42876), .B0(n13807), .C0(n13808), .Y(
        n34775) );
  OA22X1 U53733 ( .A0(net263064), .A1(n32610), .B0(n32618), .B1(n40092), .Y(
        n13807) );
  AOI222XL U53734 ( .A0(net265492), .A1(n50196), .B0(n40224), .B1(n50195),
        .C0(n40377), .C1(n50194), .Y(n13808) );
  OAI211X1 U53735 ( .A0(n32618), .A1(n42877), .B0(n13783), .C0(n13784), .Y(
        n34767) );
  OA22X1 U53736 ( .A0(net263330), .A1(n32602), .B0(n32610), .B1(n40077), .Y(
        n13783) );
  AOI222XL U53737 ( .A0(net265473), .A1(n50195), .B0(n40224), .B1(n50194),
        .C0(n40377), .C1(n50193), .Y(n13784) );
  OAI211X1 U53738 ( .A0(n32610), .A1(n42879), .B0(n13759), .C0(n13760), .Y(
        n34759) );
  OA22X1 U53739 ( .A0(net263349), .A1(n32594), .B0(n32602), .B1(n40076), .Y(
        n13759) );
  AOI222XL U53740 ( .A0(net265473), .A1(n50194), .B0(n40225), .B1(n50193),
        .C0(n40378), .C1(n50192), .Y(n13760) );
  OAI211X1 U53741 ( .A0(n32602), .A1(n42912), .B0(n13735), .C0(n13736), .Y(
        n34751) );
  OA22X1 U53742 ( .A0(net263349), .A1(n32586), .B0(n32594), .B1(n40076), .Y(
        n13735) );
  AOI222XL U53743 ( .A0(net265796), .A1(n50193), .B0(n40204), .B1(n50192),
        .C0(n40378), .C1(n50191), .Y(n13736) );
  OAI211X1 U53744 ( .A0(n32594), .A1(n42913), .B0(n13711), .C0(n13712), .Y(
        n34743) );
  AOI222XL U53745 ( .A0(net265796), .A1(n50192), .B0(n40204), .B1(n50191),
        .C0(n40378), .C1(n50190), .Y(n13712) );
  AOI222XL U53746 ( .A0(net265796), .A1(n50191), .B0(n40204), .B1(n50190),
        .C0(n40379), .C1(n50189), .Y(n13688) );
  OA22X1 U53747 ( .A0(net263387), .A1(n32562), .B0(n32570), .B1(n40074), .Y(
        n13663) );
  AOI222XL U53748 ( .A0(net265777), .A1(n50190), .B0(n40205), .B1(n50189),
        .C0(n40379), .C1(n50188), .Y(n13664) );
  OA22X1 U53749 ( .A0(net263387), .A1(n32554), .B0(n32562), .B1(n40074), .Y(
        n13639) );
  AOI222XL U53750 ( .A0(net265777), .A1(n50189), .B0(n40205), .B1(n50188),
        .C0(n40380), .C1(n50187), .Y(n13640) );
  OAI211X1 U53751 ( .A0(n32562), .A1(n42917), .B0(n13615), .C0(n13616), .Y(
        n34711) );
  OA22X1 U53752 ( .A0(net263406), .A1(n32546), .B0(n32554), .B1(n40073), .Y(
        n13615) );
  AOI222XL U53753 ( .A0(net265777), .A1(n50188), .B0(n40206), .B1(n50187),
        .C0(n40380), .C1(n50186), .Y(n13616) );
  OAI211X1 U53754 ( .A0(n32554), .A1(n42919), .B0(n13591), .C0(n13592), .Y(
        n34703) );
  OA22X1 U53755 ( .A0(net263406), .A1(n32538), .B0(n32546), .B1(n40073), .Y(
        n13591) );
  AOI222XL U53756 ( .A0(net265758), .A1(n50187), .B0(n40206), .B1(n50186),
        .C0(n40380), .C1(n50185), .Y(n13592) );
  OAI211X1 U53757 ( .A0(n32546), .A1(n42920), .B0(n13567), .C0(n13568), .Y(
        n34695) );
  OA22X1 U53758 ( .A0(net263406), .A1(n32530), .B0(n32538), .B1(n40072), .Y(
        n13567) );
  AOI222XL U53759 ( .A0(net265758), .A1(n50186), .B0(n40206), .B1(n50185),
        .C0(n40381), .C1(n50184), .Y(n13568) );
  AOI222XL U53760 ( .A0(net265758), .A1(n50185), .B0(n40207), .B1(n50184),
        .C0(n40381), .C1(n50183), .Y(n13544) );
  AOI222XL U53761 ( .A0(net265739), .A1(n50184), .B0(n40207), .B1(n50183),
        .C0(n40381), .C1(n50182), .Y(n13520) );
  OA22X1 U53762 ( .A0(net263444), .A1(n32506), .B0(n32514), .B1(n40071), .Y(
        n13495) );
  AOI222XL U53763 ( .A0(net265739), .A1(n50183), .B0(n40208), .B1(n50182),
        .C0(n40382), .C1(n50181), .Y(n13496) );
  OA22X1 U53764 ( .A0(net263444), .A1(n32498), .B0(n32506), .B1(n40070), .Y(
        n13471) );
  AOI222XL U53765 ( .A0(net265739), .A1(n50182), .B0(n40208), .B1(n50181),
        .C0(n40382), .C1(n50180), .Y(n13472) );
  OAI211X1 U53766 ( .A0(n32506), .A1(n42926), .B0(n13447), .C0(n13448), .Y(
        n34655) );
  OA22X1 U53767 ( .A0(net263463), .A1(n32490), .B0(n32498), .B1(n40070), .Y(
        n13447) );
  AOI222XL U53768 ( .A0(net265720), .A1(n50181), .B0(n40208), .B1(n50180),
        .C0(n40382), .C1(n50179), .Y(n13448) );
  OAI211X1 U53769 ( .A0(n32498), .A1(n42927), .B0(n13423), .C0(n13424), .Y(
        n34647) );
  OA22X1 U53770 ( .A0(net263254), .A1(n32482), .B0(n32490), .B1(n40080), .Y(
        n13423) );
  AOI222XL U53771 ( .A0(net265720), .A1(n50180), .B0(n40209), .B1(n50179),
        .C0(n40383), .C1(n50178), .Y(n13424) );
  OAI211X1 U53772 ( .A0(n32490), .A1(n42896), .B0(n13399), .C0(n13400), .Y(
        n34639) );
  AOI222XL U53773 ( .A0(net265720), .A1(n50179), .B0(n40209), .B1(n50178),
        .C0(n40383), .C1(n50177), .Y(n13400) );
  AOI222XL U53774 ( .A0(net265701), .A1(n50178), .B0(n40210), .B1(n50177),
        .C0(n40383), .C1(n50176), .Y(n13376) );
  AOI222XL U53775 ( .A0(net265701), .A1(n50177), .B0(n40210), .B1(n50176),
        .C0(n40384), .C1(n50175), .Y(n13352) );
  AOI222XL U53776 ( .A0(net265701), .A1(n50176), .B0(n40211), .B1(n50175),
        .C0(n40384), .C1(n50174), .Y(n13328) );
  OAI211X1 U53777 ( .A0(n32458), .A1(n42900), .B0(n13303), .C0(n13304), .Y(
        n34607) );
  OA22X1 U53778 ( .A0(net263235), .A1(n32442), .B0(n32450), .B1(n40082), .Y(
        n13303) );
  AOI222XL U53779 ( .A0(net265682), .A1(n50175), .B0(n40211), .B1(n50174),
        .C0(n40384), .C1(n50173), .Y(n13304) );
  OAI211X1 U53780 ( .A0(n32450), .A1(n42901), .B0(n13279), .C0(n13280), .Y(
        n34599) );
  OA22X1 U53781 ( .A0(net263254), .A1(n32434), .B0(n32442), .B1(n40081), .Y(
        n13279) );
  AOI222XL U53782 ( .A0(net265682), .A1(n50174), .B0(n40211), .B1(n50173),
        .C0(n40385), .C1(n50172), .Y(n13280) );
  OAI211X1 U53783 ( .A0(n32442), .A1(n42902), .B0(n13255), .C0(n13256), .Y(
        n34591) );
  OA22X1 U53784 ( .A0(net263254), .A1(n32426), .B0(n32434), .B1(n40081), .Y(
        n13255) );
  AOI222XL U53785 ( .A0(net265682), .A1(n50173), .B0(n40212), .B1(n50172),
        .C0(n40385), .C1(n50171), .Y(n13256) );
  OAI211X1 U53786 ( .A0(n32434), .A1(n42904), .B0(n13231), .C0(n13232), .Y(
        n34583) );
  OA22X1 U53787 ( .A0(net218416), .A1(n32418), .B0(n32426), .B1(n40080), .Y(
        n13231) );
  AOI222XL U53788 ( .A0(net221816), .A1(n50172), .B0(n40212), .B1(n50171),
        .C0(net216982), .C1(n50170), .Y(n13232) );
  OAI211X1 U53789 ( .A0(n32426), .A1(n42905), .B0(n13207), .C0(n13208), .Y(
        n34575) );
  AOI222XL U53790 ( .A0(net221812), .A1(n50171), .B0(n40213), .B1(n50170),
        .C0(net217010), .C1(n50169), .Y(n13208) );
  AOI222XL U53791 ( .A0(net221800), .A1(n50170), .B0(n40213), .B1(n50169),
        .C0(net216996), .C1(n50168), .Y(n13184) );
  AOI222XL U53792 ( .A0(net265644), .A1(n50169), .B0(n40213), .B1(n50168),
        .C0(net216970), .C1(n50167), .Y(n13160) );
  AOI222XL U53793 ( .A0(net265644), .A1(n50168), .B0(n40214), .B1(n50167),
        .C0(net216978), .C1(n50166), .Y(n13136) );
  OAI211X1 U53794 ( .A0(n34419), .A1(n42911), .B0(n13043), .C0(n50076), .Y(
        n34523) );
  OAI222XL U53795 ( .A0(net266654), .A1(n9656), .B0(n40159), .B1(n9655), .C0(
        n40292), .C1(n34427), .Y(n13045) );
  CLKINVX1 U53796 ( .A(n19164), .Y(n49563) );
  OAI222XL U53797 ( .A0(net266381), .A1(n9655), .B0(n40174), .B1(n34427), .C0(
        n40303), .C1(n34419), .Y(n19164) );
  CLKINVX1 U53798 ( .A(n19140), .Y(n49567) );
  OAI222XL U53799 ( .A0(net266402), .A1(n34427), .B0(n40174), .B1(n34419),
        .C0(n40303), .C1(n42064), .Y(n19140) );
  OAI222XL U53800 ( .A0(net266402), .A1(n34419), .B0(n40174), .B1(n42064),
        .C0(n40303), .C1(n42065), .Y(n19116) );
  NOR4X1 U53801 ( .A(n20023), .B(n20022), .C(n20021), .D(n20020), .Y(net211456) );
  NOR2X1 U53802 ( .A(n21214), .B(n21213), .Y(net211785) );
  NOR2X1 U53803 ( .A(n22043), .B(n22042), .Y(net212171) );
  NOR4X1 U53804 ( .A(n22041), .B(n22040), .C(n22039), .D(n22038), .Y(net212172) );
  NOR4X1 U53805 ( .A(n21777), .B(n21776), .C(n21775), .D(n21774), .Y(net212020) );
  NAND4X1 U53806 ( .A(n43506), .B(n43505), .C(n43504), .D(n43503), .Y(n12634)
         );
  NOR2X1 U53807 ( .A(n30119), .B(n30118), .Y(n43504) );
  NOR4X1 U53808 ( .A(n30117), .B(n30116), .C(n30115), .D(n30114), .Y(n43503)
         );
  NAND4X1 U53809 ( .A(n43526), .B(n43525), .C(n43524), .D(n43523), .Y(n12629)
         );
  NOR2X1 U53810 ( .A(n29759), .B(n29758), .Y(n43524) );
  NOR4X1 U53811 ( .A(n29757), .B(n29756), .C(n29755), .D(n29754), .Y(n43523)
         );
  CLKINVX1 U53812 ( .A(n19176), .Y(n49559) );
  OAI222XL U53813 ( .A0(net266444), .A1(n9663), .B0(n40182), .B1(n34431), .C0(
        n40313), .C1(n34423), .Y(n19176) );
  OAI211X1 U53814 ( .A0(n33618), .A1(n42735), .B0(n16783), .C0(n16784), .Y(
        n35767) );
  AOI222XL U53815 ( .A0(net264922), .A1(n50320), .B0(n40258), .B1(n50319),
        .C0(n40337), .C1(n50318), .Y(n16784) );
  NAND4X1 U53816 ( .A(n43481), .B(n43480), .C(n43479), .D(n43478), .Y(n12640)
         );
  NOR2X1 U53817 ( .A(n30300), .B(n30299), .Y(n43479) );
  NOR4X1 U53818 ( .A(n30298), .B(n30297), .C(n30296), .D(n30295), .Y(n43478)
         );
  NAND4X1 U53819 ( .A(n44367), .B(n44366), .C(n44365), .D(n44364), .Y(n12618)
         );
  NOR2X1 U53820 ( .A(n26148), .B(n26147), .Y(n44365) );
  NOR4X1 U53821 ( .A(n26146), .B(n26145), .C(n26144), .D(n26143), .Y(n44364)
         );
  NAND4X1 U53822 ( .A(n43533), .B(n43532), .C(n43531), .D(n43530), .Y(n12624)
         );
  NOR2X1 U53823 ( .A(n29578), .B(n29577), .Y(n43531) );
  NOR4X1 U53824 ( .A(n29576), .B(n29575), .C(n29574), .D(n29573), .Y(n43530)
         );
  NAND4X1 U53825 ( .A(n45546), .B(n45545), .C(n45544), .D(n45543), .Y(
        net209101) );
  NOR2X1 U53826 ( .A(n24640), .B(n24638), .Y(n45544) );
  NOR4X1 U53827 ( .A(n24637), .B(n24636), .C(n24635), .D(n24634), .Y(n45543)
         );
  XNOR2X1 U53828 ( .A(n36734), .B(n32722), .Y(net212059) );
  NOR2X1 U53829 ( .A(n21841), .B(n21840), .Y(net212060) );
  NOR4X1 U53830 ( .A(n21839), .B(n21838), .C(n21837), .D(n21836), .Y(net212061) );
  NAND4X1 U53831 ( .A(n43446), .B(n43445), .C(n43444), .D(n43443), .Y(n12643)
         );
  NOR2X1 U53832 ( .A(n30542), .B(n30541), .Y(n43444) );
  NOR4X1 U53833 ( .A(n30540), .B(n30539), .C(n30538), .D(n30537), .Y(n43443)
         );
  NOR4X1 U53834 ( .A(n24303), .B(n24302), .C(n24301), .D(n24300), .Y(net213500) );
  NOR2X1 U53835 ( .A(n24215), .B(n24214), .Y(net212080) );
  NOR4X1 U53836 ( .A(n24213), .B(n24212), .C(n24211), .D(n24210), .Y(net212081) );
  NOR2X1 U53837 ( .A(n24285), .B(n24284), .Y(net212050) );
  NOR4X1 U53838 ( .A(n24283), .B(n24282), .C(n24281), .D(n24280), .Y(net212051) );
  NOR2X1 U53839 ( .A(n26178), .B(n26177), .Y(net213207) );
  NOR4X1 U53840 ( .A(n26176), .B(n26175), .C(n26174), .D(n26173), .Y(net213208) );
  NAND4X1 U53841 ( .A(n47279), .B(n47278), .C(n47277), .D(n47276), .Y(n12183)
         );
  NOR2X1 U53842 ( .A(n23646), .B(n23645), .Y(n47277) );
  NOR4X1 U53843 ( .A(n23644), .B(n23643), .C(n23642), .D(n23641), .Y(n47276)
         );
  NOR4X1 U53844 ( .A(n24405), .B(n24404), .C(n24403), .D(n24402), .Y(net213540) );
  NOR4X1 U53845 ( .A(n24263), .B(n24262), .C(n24261), .D(n24260), .Y(net213480) );
  NOR4X1 U53846 ( .A(n24617), .B(n24616), .C(n24615), .D(n24614), .Y(net213636) );
  NAND4X1 U53847 ( .A(n44389), .B(n44388), .C(n44387), .D(n44386), .Y(
        net209701) );
  NOR2X1 U53848 ( .A(n25968), .B(n25967), .Y(n44387) );
  NOR4X1 U53849 ( .A(n25966), .B(n25965), .C(n25964), .D(n25963), .Y(n44386)
         );
  NOR4X1 U53850 ( .A(n23624), .B(n23623), .C(n23622), .D(n23621), .Y(net213320) );
  NOR2X1 U53851 ( .A(n25848), .B(n25847), .Y(net215017) );
  NOR4X1 U53852 ( .A(n25846), .B(n25845), .C(n25844), .D(n25843), .Y(net215018) );
  NOR2X1 U53853 ( .A(n26238), .B(n26237), .Y(net215098) );
  NOR4X1 U53854 ( .A(n26236), .B(n26235), .C(n26234), .D(n26233), .Y(net215099) );
  NOR4X1 U53855 ( .A(n24415), .B(n24414), .C(n24413), .D(n24412), .Y(net213545) );
  NOR2X1 U53856 ( .A(n26028), .B(n26027), .Y(net215053) );
  NOR4X1 U53857 ( .A(n26026), .B(n26025), .C(n26024), .D(n26023), .Y(net215054) );
  NOR2X1 U53858 ( .A(n23321), .B(n23320), .Y(net213233) );
  NOR4X1 U53859 ( .A(n23319), .B(n23318), .C(n23317), .D(n23316), .Y(net213234) );
  NOR2X1 U53860 ( .A(n22073), .B(n22072), .Y(net212186) );
  NOR4X1 U53861 ( .A(n22071), .B(n22070), .C(n22069), .D(n22068), .Y(net212187) );
  NOR4X1 U53862 ( .A(n21809), .B(n21808), .C(n21807), .D(n21806), .Y(net212041) );
  NAND4X1 U53863 ( .A(n46703), .B(n46702), .C(n46701), .D(n46700), .Y(n11519)
         );
  NOR2X1 U53864 ( .A(n21668), .B(n21667), .Y(n46701) );
  NOR4X1 U53865 ( .A(n21666), .B(n21665), .C(n21664), .D(n21663), .Y(n46700)
         );
  NOR2X1 U53866 ( .A(n21224), .B(n21223), .Y(net211790) );
  NOR2X1 U53867 ( .A(n22053), .B(n22052), .Y(net212176) );
  NOR4X1 U53868 ( .A(n22051), .B(n22050), .C(n22049), .D(n22048), .Y(net212177) );
  XNOR2X1 U53869 ( .A(n36733), .B(n32738), .Y(net212069) );
  NOR2X1 U53870 ( .A(n21861), .B(n21860), .Y(net212070) );
  NOR4X1 U53871 ( .A(n21859), .B(n21858), .C(n21857), .D(n21856), .Y(net212071) );
  NOR2X1 U53872 ( .A(n21658), .B(n21657), .Y(net210499) );
  XNOR2X1 U53873 ( .A(n36736), .B(n32818), .Y(net212130) );
  NOR2X1 U53874 ( .A(n21983), .B(n21982), .Y(net212131) );
  NOR4X1 U53875 ( .A(n21981), .B(n21980), .C(n21979), .D(n21978), .Y(net212132) );
  NOR2X1 U53876 ( .A(n21254), .B(n21253), .Y(net210623) );
  NOR2X1 U53877 ( .A(n21851), .B(n21850), .Y(net212065) );
  OA22X1 U53878 ( .A0(net263805), .A1(n32932), .B0(n32940), .B1(n40050), .Y(
        n14773) );
  AOI222XL U53879 ( .A0(net266081), .A1(n51296), .B0(n40186), .B1(n51295),
        .C0(net216982), .C1(n51294), .Y(n14774) );
  AOI222XL U53880 ( .A0(net266081), .A1(n50236), .B0(n40186), .B1(n50235),
        .C0(net216980), .C1(n50234), .Y(n14768) );
  NAND4X1 U53881 ( .A(n45581), .B(n45580), .C(n45579), .D(n45578), .Y(n12230)
         );
  XNOR2X1 U53882 ( .A(n36841), .B(n32874), .Y(n45580) );
  NOR2X1 U53883 ( .A(n24427), .B(n24426), .Y(n45579) );
  NOR4X1 U53884 ( .A(n24425), .B(n24424), .C(n24423), .D(n24422), .Y(n45578)
         );
  NAND4X1 U53885 ( .A(n43461), .B(n43460), .C(n43459), .D(n43458), .Y(n12648)
         );
  NOR2X1 U53886 ( .A(n30512), .B(n30511), .Y(n43459) );
  NOR4X1 U53887 ( .A(n30510), .B(n30509), .C(n30508), .D(n30507), .Y(n43458)
         );
  NAND4X1 U53888 ( .A(n43441), .B(n43440), .C(n43439), .D(n43438), .Y(n12639)
         );
  NOR2X1 U53889 ( .A(n30572), .B(n30571), .Y(n43439) );
  NOR4X1 U53890 ( .A(n30570), .B(n30569), .C(n30568), .D(n30567), .Y(n43438)
         );
  NOR4X1 U53891 ( .A(n24313), .B(n24312), .C(n24311), .D(n24310), .Y(net213505) );
  NAND4X1 U53892 ( .A(n46657), .B(n46656), .C(n46655), .D(n46654), .Y(n10644)
         );
  XNOR2X1 U53893 ( .A(n36734), .B(n32706), .Y(n46656) );
  NOR2X1 U53894 ( .A(n21913), .B(n21911), .Y(n46655) );
  NOR4X1 U53895 ( .A(n21910), .B(n21909), .C(n21908), .D(n21907), .Y(n46654)
         );
  INVX3 U53896 ( .A(n33028), .Y(n51303) );
  INVX3 U53897 ( .A(n33020), .Y(n51302) );
  INVX3 U53898 ( .A(n33012), .Y(n51301) );
  INVX3 U53899 ( .A(n33004), .Y(n51300) );
  NOR2X1 U53900 ( .A(n22023), .B(n22022), .Y(net212161) );
  NOR4X1 U53901 ( .A(n22021), .B(n22020), .C(n22019), .D(n22018), .Y(net212162) );
  XNOR2X1 U53902 ( .A(n36734), .B(n32746), .Y(net212044) );
  NOR2X1 U53903 ( .A(n21821), .B(n21820), .Y(net212045) );
  NOR4X1 U53904 ( .A(n21819), .B(n21818), .C(n21817), .D(n21816), .Y(net212046) );
  OAI211X1 U53905 ( .A0(n9678), .A1(net266780), .B0(n9807), .C0(n9808), .Y(
        n34510) );
  AOI221XL U53906 ( .A0(n9759), .A1(n9809), .B0(n9770), .B1(n9810), .C0(n9811),
        .Y(n9808) );
  NAND2BX1 U53907 ( .AN(n9878), .B(n9771), .Y(n9873) );
  NOR2X1 U53908 ( .A(n22013), .B(n22012), .Y(net212146) );
  NOR4X1 U53909 ( .A(n22011), .B(n22010), .C(n22009), .D(n22008), .Y(net212147) );
  NOR2X1 U53910 ( .A(n21993), .B(n21992), .Y(net212136) );
  NOR4X1 U53911 ( .A(n21991), .B(n21990), .C(n21989), .D(n21988), .Y(net212137) );
  NAND4X1 U53912 ( .A(n47911), .B(n47910), .C(n47909), .D(n47908), .Y(n12847)
         );
  NOR2X1 U53913 ( .A(n21963), .B(n21962), .Y(n47909) );
  NOR4X1 U53914 ( .A(n21961), .B(n21960), .C(n21959), .D(n21958), .Y(n47908)
         );
  NAND4X1 U53915 ( .A(n47864), .B(n47863), .C(n47862), .D(n47861), .Y(n12831)
         );
  NOR2X1 U53916 ( .A(n20918), .B(n20917), .Y(n47862) );
  NOR4X1 U53917 ( .A(n20916), .B(n20915), .C(n20914), .D(n20913), .Y(n47861)
         );
  NAND4X1 U53918 ( .A(n47876), .B(n47875), .C(n47874), .D(n47873), .Y(n12811)
         );
  NOR2X1 U53919 ( .A(n20444), .B(n20443), .Y(n47874) );
  NOR4X1 U53920 ( .A(n20442), .B(n20441), .C(n20440), .D(n20439), .Y(n47873)
         );
  NOR2X1 U53921 ( .A(n22094), .B(n22093), .Y(net212196) );
  NAND4X1 U53922 ( .A(n45602), .B(n45601), .C(n45600), .D(n45599), .Y(
        net212037) );
  NOR2X1 U53923 ( .A(n24275), .B(n24274), .Y(n45600) );
  NOR4X1 U53924 ( .A(n24273), .B(n24272), .C(n24271), .D(n24270), .Y(n45599)
         );
  NAND4X1 U53925 ( .A(n45611), .B(n45610), .C(n45609), .D(n45608), .Y(
        net212088) );
  NOR2X1 U53926 ( .A(n24205), .B(n24204), .Y(n45609) );
  NOR4X1 U53927 ( .A(n24203), .B(n24202), .C(n24201), .D(n24200), .Y(n45608)
         );
  NAND4X1 U53928 ( .A(n45557), .B(n45556), .C(n45555), .D(n45554), .Y(
        net211640) );
  XNOR2X1 U53929 ( .A(n36839), .B(n32650), .Y(n45556) );
  NOR2X1 U53930 ( .A(n24609), .B(n24608), .Y(n45555) );
  NOR4X1 U53931 ( .A(n24607), .B(n24606), .C(n24605), .D(n24604), .Y(n45554)
         );
  NAND4X1 U53932 ( .A(n45536), .B(n45535), .C(n45534), .D(n45533), .Y(
        net211602) );
  NOR2X1 U53933 ( .A(n24661), .B(n24660), .Y(n45534) );
  NOR4X1 U53934 ( .A(n24659), .B(n24658), .C(n24657), .D(n24656), .Y(n45533)
         );
  NAND4X1 U53935 ( .A(n45551), .B(n45550), .C(n45549), .D(n45548), .Y(
        net211584) );
  XNOR2X1 U53936 ( .A(n36843), .B(n32562), .Y(n45550) );
  NOR2X1 U53937 ( .A(n24629), .B(n24628), .Y(n45549) );
  NOR4X1 U53938 ( .A(n24627), .B(n24626), .C(n24625), .D(n24624), .Y(n45548)
         );
  NAND4X1 U53939 ( .A(n45714), .B(n45713), .C(n45712), .D(n45711), .Y(
        net211568) );
  NOR2X1 U53940 ( .A(n23636), .B(n23635), .Y(n45712) );
  NOR4X1 U53941 ( .A(n23634), .B(n23633), .C(n23632), .D(n23631), .Y(n45711)
         );
  NAND4X1 U53942 ( .A(n44361), .B(n44360), .C(n44359), .D(n44358), .Y(
        net213230) );
  NOR2X1 U53943 ( .A(n26268), .B(n26267), .Y(n44359) );
  NOR4X1 U53944 ( .A(n26266), .B(n26265), .C(n26264), .D(n26263), .Y(n44358)
         );
  XNOR2X1 U53945 ( .A(n36735), .B(n32690), .Y(net212105) );
  NOR2X1 U53946 ( .A(n21923), .B(n21922), .Y(net212106) );
  NOR4X1 U53947 ( .A(n21921), .B(n21920), .C(n21919), .D(n21918), .Y(net212107) );
  NAND4X1 U53948 ( .A(n46622), .B(n46621), .C(n46620), .D(n46619), .Y(n13023)
         );
  NOR2X1 U53949 ( .A(n22063), .B(n22062), .Y(n46620) );
  NOR4X1 U53950 ( .A(n22061), .B(n22060), .C(n22059), .D(n22058), .Y(n46619)
         );
  NAND4X1 U53951 ( .A(n46671), .B(n46670), .C(n46669), .D(n46668), .Y(n13025)
         );
  NOR2X1 U53952 ( .A(n21801), .B(n21799), .Y(n46669) );
  NOR4X1 U53953 ( .A(n21798), .B(n21797), .C(n21796), .D(n21795), .Y(n46668)
         );
  NAND4X1 U53954 ( .A(n46853), .B(n46852), .C(n46851), .D(n46850), .Y(n13022)
         );
  NOR2X1 U53955 ( .A(n21244), .B(n21243), .Y(n46851) );
  NOR4X1 U53956 ( .A(n21242), .B(n21241), .C(n21240), .D(n21239), .Y(n46850)
         );
  NOR2X1 U53957 ( .A(n21831), .B(n21830), .Y(net212055) );
  NOR4X1 U53958 ( .A(n20853), .B(n20852), .C(n20851), .D(n20850), .Y(net211606) );
  NOR4X1 U53959 ( .A(n20885), .B(n20884), .C(n20883), .D(n20882), .Y(net211626) );
  NAND4X1 U53960 ( .A(n46989), .B(n46988), .C(n46987), .D(n46986), .Y(
        net209974) );
  NOR2X1 U53961 ( .A(n20476), .B(n20475), .Y(n46987) );
  NOR4X1 U53962 ( .A(n20474), .B(n20473), .C(n20472), .D(n20471), .Y(n46986)
         );
  OAI22XL U53963 ( .A0(n50145), .A1(n9690), .B0(n9693), .B1(n50144), .Y(
        nxt_state[0]) );
  NOR4X1 U53964 ( .A(n9695), .B(n9696), .C(n9697), .D(n9698), .Y(n9693) );
  XNOR2X1 U53965 ( .A(n42316), .B(nxt_data_num[0]), .Y(n9698) );
  XNOR2X1 U53966 ( .A(n32398), .B(nxt_data_num[2]), .Y(n9696) );
  NAND4X1 U53967 ( .A(n47916), .B(n47915), .C(n47914), .D(n47913), .Y(n12851)
         );
  NOR2X1 U53968 ( .A(n21973), .B(n21972), .Y(n47914) );
  NOR4X1 U53969 ( .A(n21971), .B(n21970), .C(n21969), .D(n21968), .Y(n47913)
         );
  NOR4X1 U53970 ( .A(n20926), .B(n20925), .C(n20924), .D(n20923), .Y(net210356) );
  NOR2X1 U53971 ( .A(n20455), .B(n20453), .Y(net210350) );
  XNOR2X1 U53972 ( .A(n36735), .B(n32698), .Y(net212115) );
  NOR2X1 U53973 ( .A(n21933), .B(n21932), .Y(net212116) );
  NOR4X1 U53974 ( .A(n21931), .B(n21930), .C(n21929), .D(n21928), .Y(net212117) );
  NOR4X1 U53975 ( .A(n22081), .B(n22080), .C(n22079), .D(n22078), .Y(net212192) );
  NOR2X1 U53976 ( .A(n20466), .B(n20464), .Y(net211565) );
  XNOR2X1 U53977 ( .A(n36770), .B(n32609), .Y(net211630) );
  NOR2X1 U53978 ( .A(n20897), .B(n20896), .Y(net211631) );
  XNOR2X1 U53979 ( .A(n36735), .B(n32802), .Y(net212125) );
  NOR2X1 U53980 ( .A(n21953), .B(n21952), .Y(net212126) );
  NOR2X1 U53981 ( .A(n22033), .B(n22032), .Y(net212166) );
  NAND4X1 U53982 ( .A(n46638), .B(n46637), .C(n46636), .D(n46635), .Y(n13024)
         );
  NOR2X1 U53983 ( .A(n22003), .B(n22002), .Y(n46636) );
  NOR4X1 U53984 ( .A(n22001), .B(n22000), .C(n21999), .D(n21998), .Y(n46635)
         );
  NOR2X1 U53985 ( .A(n10965), .B(n47907), .Y(n47911) );
  NOR2X1 U53986 ( .A(n10966), .B(n46666), .Y(net212038) );
  NOR2X1 U53987 ( .A(net260527), .B(n43486), .Y(net216364) );
  NOR2X1 U53988 ( .A(n10064), .B(n44352), .Y(net215114) );
  XOR2X1 U53989 ( .A(n32484), .B(n36821), .Y(n44352) );
  NOR2X1 U53990 ( .A(n10776), .B(n47048), .Y(net211453) );
  NOR2X1 U53991 ( .A(n10434), .B(n44405), .Y(net214997) );
  XOR2X1 U53992 ( .A(n32572), .B(n36825), .Y(n44405) );
  NOR2X1 U53993 ( .A(n10485), .B(n46085), .Y(net212836) );
  NOR2X1 U53994 ( .A(n10436), .B(n44399), .Y(net215015) );
  XOR2X1 U53995 ( .A(n32580), .B(n36825), .Y(n44399) );
  NOR2X1 U53996 ( .A(n10206), .B(n46649), .Y(net212104) );
  NOR2X1 U53997 ( .A(n10471), .B(n45604), .Y(net213472) );
  NOR2X1 U53998 ( .A(n10433), .B(n43535), .Y(net216175) );
  NOR2X1 U53999 ( .A(n10905), .B(n46617), .Y(net212184) );
  NOR2X1 U54000 ( .A(n10904), .B(n46857), .Y(net211778) );
  NOR2X1 U54001 ( .A(n10487), .B(n46080), .Y(n46084) );
  AOI222XL U54002 ( .A0(n36928), .A1(n50135), .B0(n9732), .B1(n50147), .C0(
        n32398), .C1(n9733), .Y(n9728) );
  OA21XL U54003 ( .A0(n9730), .A1(n43042), .B0(n9712), .Y(n9727) );
  OAI21XL U54004 ( .A0(n9689), .A1(n9721), .B0(n32398), .Y(n9729) );
  NOR2X1 U54005 ( .A(n10469), .B(n45605), .Y(net213467) );
  NOR2X1 U54006 ( .A(n39470), .B(n43442), .Y(n43446) );
  NOR2X1 U54007 ( .A(n10205), .B(n46643), .Y(net212114) );
  NOR2X1 U54008 ( .A(n10470), .B(n45607), .Y(n45611) );
  NOR2X1 U54009 ( .A(n_cell_303546_net275987), .B(n46610), .Y(n46614) );
  NOR2X1 U54010 ( .A(n10302), .B(n43516), .Y(net216238) );
  NAND4X1 U54011 ( .A(n48556), .B(n9983), .C(n48555), .D(n48554), .Y(n34512)
         );
  AOI21XL U54012 ( .A0(codeword[5]), .A1(net264532), .B0(n48553), .Y(n48556)
         );
  AOI2BB1X1 U54013 ( .A0N(n42991), .A1N(n10059), .B0(n10060), .Y(n9983) );
  NOR2X1 U54014 ( .A(n11915), .B(n45591), .Y(net213497) );
  NOR2X1 U54015 ( .A(n11551), .B(n44345), .Y(net215141) );
  XOR2X1 U54016 ( .A(n32476), .B(n36830), .Y(n44345) );
  NOR2X1 U54017 ( .A(n_cell_303546_net275967), .B(n45583), .Y(net213537) );
  XOR2X1 U54018 ( .A(n32865), .B(n36785), .Y(n45583) );
  NOR2X1 U54019 ( .A(n10480), .B(n45573), .Y(net213567) );
  NOR2X1 U54020 ( .A(n10983), .B(n46623), .Y(net212174) );
  NOR2X1 U54021 ( .A(n10448), .B(n47275), .Y(n47279) );
  NOR2X1 U54022 ( .A(n_cell_303546_net275959), .B(n46624), .Y(net212169) );
  NOR2X1 U54023 ( .A(n11567), .B(n44384), .Y(net215042) );
  XOR2X1 U54024 ( .A(n32604), .B(n36827), .Y(n44384) );
  NOR2X1 U54025 ( .A(n11901), .B(n45547), .Y(n45551) );
  XOR2X1 U54026 ( .A(n32561), .B(n36779), .Y(n45547) );
  NOR2X1 U54027 ( .A(n10923), .B(n47049), .Y(net211448) );
  NOR2X1 U54028 ( .A(n10960), .B(n46661), .Y(net212063) );
  NOR2X1 U54029 ( .A(n10992), .B(n46855), .Y(net211788) );
  NOR2X1 U54030 ( .A(n11943), .B(n45576), .Y(net213552) );
  XOR2X1 U54031 ( .A(n32881), .B(n36777), .Y(n45576) );
  NOR2X1 U54032 ( .A(n11578), .B(n44615), .Y(n44619) );
  NOR2X1 U54033 ( .A(n11916), .B(n46658), .Y(net212078) );
  NOR2X1 U54034 ( .A(net260299), .B(n45590), .Y(net213502) );
  NOR2X1 U54035 ( .A(net259645), .B(n43418), .Y(n43422) );
  NOR2X1 U54036 ( .A(n11550), .B(n44321), .Y(n44325) );
  XOR2X1 U54037 ( .A(n32452), .B(n36829), .Y(n44321) );
  NOR2X1 U54038 ( .A(n11924), .B(n46664), .Y(net212048) );
  NOR2X1 U54039 ( .A(n10969), .B(n47912), .Y(n47916) );
  NOR2X1 U54040 ( .A(n11935), .B(n45572), .Y(net213572) );
  XOR2X1 U54041 ( .A(n32817), .B(n36785), .Y(n45572) );
  NOR2X1 U54042 ( .A(n11595), .B(n43514), .Y(net216256) );
  NOR2X1 U54043 ( .A(n11601), .B(n43502), .Y(n43506) );
  NOR2X1 U54044 ( .A(n10958), .B(n46662), .Y(net212058) );
  NOR2X1 U54045 ( .A(n10990), .B(n46856), .Y(net211783) );
  NOR2X1 U54046 ( .A(net259641), .B(n43457), .Y(n43461) );
  NOR2X1 U54047 ( .A(n10976), .B(n46639), .Y(net212134) );
  NOR2X1 U54048 ( .A(n11600), .B(n43495), .Y(net216319) );
  NOR2X1 U54049 ( .A(n11886), .B(n45788), .Y(net213236) );
  NOR2X1 U54050 ( .A(n11874), .B(n44362), .Y(net215096) );
  XOR2X1 U54051 ( .A(n32516), .B(n36830), .Y(n44362) );
  NOR2X1 U54052 ( .A(net259661), .B(n43540), .Y(net216166) );
  NOR2X1 U54053 ( .A(n11594), .B(n43513), .Y(net216265) );
  NOR2X1 U54054 ( .A(n_cell_303546_net276365), .B(n44620), .Y(net214688) );
  NOR2X1 U54055 ( .A(n10991), .B(n46849), .Y(n46853) );
  NOR2X1 U54056 ( .A(n12392), .B(n46652), .Y(net212089) );
  NOR2X1 U54057 ( .A(n10974), .B(n46640), .Y(net212129) );
  NOR2X1 U54058 ( .A(n_cell_303546_net275923), .B(n46626), .Y(net212159) );
  NOR2X1 U54059 ( .A(n10447), .B(n47867), .Y(n47871) );
  NAND4BX1 U54060 ( .AN(n47950), .B(n49490), .C(n47949), .D(n9777), .Y(n34509)
         );
  NAND3X1 U54061 ( .A(n9773), .B(n9771), .C(n9802), .Y(n47949) );
  NOR2X1 U54062 ( .A(n9778), .B(n9779), .Y(n9777) );
  NOR2X1 U54063 ( .A(n11549), .B(n47270), .Y(n47274) );
  NOR2X1 U54064 ( .A(n11558), .B(n45791), .Y(net213220) );
  NOR2X1 U54065 ( .A(n11883), .B(n45789), .Y(net213231) );
  NOR2X1 U54066 ( .A(n11605), .B(n46627), .Y(net212154) );
  NOR2X1 U54067 ( .A(n11606), .B(n43493), .Y(net216337) );
  NOR2X1 U54068 ( .A(n12804), .B(n45575), .Y(net213557) );
  XOR2X1 U54069 ( .A(n32825), .B(n36776), .Y(n45575) );
  NOR2X1 U54070 ( .A(n_cell_303546_net276178), .B(n46673), .Y(net212022) );
  NOR2X1 U54071 ( .A(n40415), .B(n43501), .Y(net216301) );
  NOR2X1 U54072 ( .A(net260295), .B(n45553), .Y(n45557) );
  NOR2X1 U54073 ( .A(n10968), .B(n46641), .Y(net212124) );
  NOR2X1 U54074 ( .A(n11907), .B(n45559), .Y(net213618) );
  XOR2X1 U54075 ( .A(n32625), .B(n36786), .Y(n45559) );
  NOR2X1 U54076 ( .A(n_cell_303546_net275998), .B(n46634), .Y(n46638) );
  NOR2X1 U54077 ( .A(n10801), .B(n47758), .Y(net210621) );
  NOR2X1 U54078 ( .A(net260431), .B(n46078), .Y(net212851) );
  NOR2X1 U54079 ( .A(n10483), .B(n47753), .Y(n47757) );
  NOR2X1 U54080 ( .A(n11917), .B(n45592), .Y(n45596) );
  NOR2X1 U54081 ( .A(n11942), .B(n45577), .Y(n45581) );
  XOR2X1 U54082 ( .A(n32873), .B(n36777), .Y(n45577) );
  NOR2X1 U54083 ( .A(n11885), .B(n45796), .Y(net213195) );
  NOR2X1 U54084 ( .A(net260247), .B(n46079), .Y(net212846) );
  NOR2X1 U54085 ( .A(n12803), .B(n45585), .Y(net213527) );
  NOR2X1 U54086 ( .A(n12807), .B(n45558), .Y(net213623) );
  NOR2X1 U54087 ( .A(n12806), .B(n46644), .Y(n46648) );
  NOR2X1 U54088 ( .A(n40411), .B(n43507), .Y(net216283) );
  NOR2X1 U54089 ( .A(n10957), .B(n46663), .Y(net212053) );
  NOR2X1 U54090 ( .A(n11934), .B(n45586), .Y(net213522) );
  NOR2X1 U54091 ( .A(n11925), .B(n45617), .Y(net213447) );
  NOR2X1 U54092 ( .A(n10946), .B(n47860), .Y(n47864) );
  NOR2X1 U54093 ( .A(n12165), .B(n46628), .Y(n46632) );
  NOR2X1 U54094 ( .A(n_cell_303546_net275934), .B(n43448), .Y(n43452) );
  NOR2X1 U54095 ( .A(n11620), .B(n43409), .Y(n43413) );
  NOR2X1 U54096 ( .A(n11565), .B(n44383), .Y(net215051) );
  XOR2X1 U54097 ( .A(n32596), .B(n36828), .Y(n44383) );
  NOR2X1 U54098 ( .A(net259649), .B(n43437), .Y(n43441) );
  NOR2X1 U54099 ( .A(net259653), .B(n43477), .Y(n43481) );
  NOR2X1 U54100 ( .A(net259626), .B(n43521), .Y(net216229) );
  NOR2X1 U54101 ( .A(n11869), .B(n43527), .Y(net216211) );
  NOR2X1 U54102 ( .A(n11870), .B(n43534), .Y(net216184) );
  NOR2X1 U54103 ( .A(n11568), .B(n44385), .Y(n44389) );
  XOR2X1 U54104 ( .A(n32612), .B(n36829), .Y(n44385) );
  NOR2X1 U54105 ( .A(n40422), .B(n43522), .Y(n43526) );
  NOR2X1 U54106 ( .A(n11556), .B(n44351), .Y(net215123) );
  XOR2X1 U54107 ( .A(n32492), .B(n36821), .Y(n44351) );
  NOR2X1 U54108 ( .A(n11576), .B(n44363), .Y(n44367) );
  XOR2X1 U54109 ( .A(n32652), .B(n36828), .Y(n44363) );
  NOR2X1 U54110 ( .A(n10973), .B(n46642), .Y(net212119) );
  NOR2X1 U54111 ( .A(n11884), .B(n45710), .Y(n45714) );
  NOR2X1 U54112 ( .A(n40418), .B(n43515), .Y(net216247) );
  NOR2X1 U54113 ( .A(n11555), .B(n45794), .Y(net213205) );
  NOR2X1 U54114 ( .A(n11575), .B(n44610), .Y(n44614) );
  NOR2X1 U54115 ( .A(n11932), .B(n45587), .Y(net213517) );
  NOR2X1 U54116 ( .A(n11906), .B(n45561), .Y(net213608) );
  NOR2X1 U54117 ( .A(n12166), .B(n45598), .Y(n45602) );
  NOR2X1 U54118 ( .A(net259873), .B(n46633), .Y(net212144) );
  NOR2X1 U54119 ( .A(n12168), .B(n45606), .Y(net213462) );
  NOR2X1 U54120 ( .A(net259747), .B(n47792), .Y(n47796) );
  NOR2X1 U54121 ( .A(n10464), .B(n45597), .Y(net213487) );
  NOR2X1 U54122 ( .A(n10947), .B(n46975), .Y(net211623) );
  NOR2X1 U54123 ( .A(n10940), .B(n46974), .Y(net211629) );
  NOR2X1 U54124 ( .A(n10959), .B(n46660), .Y(net212068) );
  NOR2X1 U54125 ( .A(n10319), .B(n43494), .Y(net216328) );
  NOR2X1 U54126 ( .A(n10938), .B(n46979), .Y(net211603) );
  NAND4X1 U54127 ( .A(n19141), .B(n48560), .C(n48559), .D(n48558), .Y(n36553)
         );
  NAND2X1 U54128 ( .A(n43000), .B(n48568), .Y(n48559) );
  NAND4X1 U54129 ( .A(n19117), .B(n48564), .C(n48563), .D(n48562), .Y(n36545)
         );
  NAND2X1 U54130 ( .A(n43000), .B(n41387), .Y(n48563) );
  NAND4X1 U54131 ( .A(n19093), .B(n48567), .C(n48566), .D(n48565), .Y(n36537)
         );
  NAND2X1 U54132 ( .A(n43000), .B(n48575), .Y(n48566) );
  NAND4X1 U54133 ( .A(n19069), .B(n48571), .C(n48570), .D(n48569), .Y(n36529)
         );
  NAND2X1 U54134 ( .A(n43000), .B(n48579), .Y(n48570) );
  NAND4X1 U54135 ( .A(n19045), .B(n48574), .C(n48573), .D(n48572), .Y(n36521)
         );
  NAND2X1 U54136 ( .A(n43000), .B(n48583), .Y(n48573) );
  NAND4X1 U54137 ( .A(n19021), .B(n48578), .C(n48577), .D(n48576), .Y(n36513)
         );
  NAND2X1 U54138 ( .A(n42999), .B(n41270), .Y(n48577) );
  NAND4X1 U54139 ( .A(n18997), .B(n48582), .C(n48581), .D(n48580), .Y(n36505)
         );
  NAND2X1 U54140 ( .A(n42999), .B(n48590), .Y(n48581) );
  NAND4X1 U54141 ( .A(n18973), .B(n48586), .C(n48585), .D(n48584), .Y(n36497)
         );
  NAND2X1 U54142 ( .A(n42999), .B(n48594), .Y(n48585) );
  NAND4X1 U54143 ( .A(n18949), .B(n48589), .C(n48588), .D(n48587), .Y(n36489)
         );
  NAND2X1 U54144 ( .A(n42999), .B(n48598), .Y(n48588) );
  NAND4X1 U54145 ( .A(n18925), .B(n48593), .C(n48592), .D(n48591), .Y(n36481)
         );
  NAND2X1 U54146 ( .A(n42999), .B(n48602), .Y(n48592) );
  NAND4X1 U54147 ( .A(n18901), .B(n48597), .C(n48596), .D(n48595), .Y(n36473)
         );
  NAND2X1 U54148 ( .A(n42999), .B(n48606), .Y(n48596) );
  NAND4X1 U54149 ( .A(n18877), .B(n48601), .C(n48600), .D(n48599), .Y(n36465)
         );
  NAND2X1 U54150 ( .A(n42999), .B(n48610), .Y(n48600) );
  NAND4X1 U54151 ( .A(n18853), .B(n48605), .C(n48604), .D(n48603), .Y(n36457)
         );
  NAND2X1 U54152 ( .A(n42999), .B(n48614), .Y(n48604) );
  NAND4X1 U54153 ( .A(n18829), .B(n48609), .C(n48608), .D(n48607), .Y(n36449)
         );
  NAND2X1 U54154 ( .A(n42999), .B(n48618), .Y(n48608) );
  NAND4X1 U54155 ( .A(n18805), .B(n48613), .C(n48612), .D(n48611), .Y(n36441)
         );
  NAND2X1 U54156 ( .A(n42999), .B(n48622), .Y(n48612) );
  NAND4X1 U54157 ( .A(n18781), .B(n48617), .C(n48616), .D(n48615), .Y(n36433)
         );
  NAND2X1 U54158 ( .A(n42999), .B(n48626), .Y(n48616) );
  NAND4X1 U54159 ( .A(n18757), .B(n48621), .C(n48620), .D(n48619), .Y(n36425)
         );
  NAND2X1 U54160 ( .A(n42999), .B(n48630), .Y(n48620) );
  NAND4X1 U54161 ( .A(n18733), .B(n48625), .C(n48624), .D(n48623), .Y(n36417)
         );
  NAND2X1 U54162 ( .A(n42999), .B(n48634), .Y(n48624) );
  NAND4X1 U54163 ( .A(n18709), .B(n48629), .C(n48628), .D(n48627), .Y(n36409)
         );
  NAND2X1 U54164 ( .A(n42993), .B(n48638), .Y(n48628) );
  NAND4X1 U54165 ( .A(n18685), .B(n48633), .C(n48632), .D(n48631), .Y(n36401)
         );
  NAND2X1 U54166 ( .A(n43001), .B(n48642), .Y(n48632) );
  NAND4X1 U54167 ( .A(n18661), .B(n48637), .C(n48636), .D(n48635), .Y(n36393)
         );
  NAND2X1 U54168 ( .A(n42997), .B(n48646), .Y(n48636) );
  NAND4X1 U54169 ( .A(n18637), .B(n48641), .C(n48640), .D(n48639), .Y(n36385)
         );
  NAND2X1 U54170 ( .A(n42993), .B(n48650), .Y(n48640) );
  NAND4X1 U54171 ( .A(n18613), .B(n48645), .C(n48644), .D(n48643), .Y(n36377)
         );
  NAND2X1 U54172 ( .A(n43005), .B(n48654), .Y(n48644) );
  NAND4X1 U54173 ( .A(n18589), .B(n48649), .C(n48648), .D(n48647), .Y(n36369)
         );
  NAND2X1 U54174 ( .A(n42999), .B(n48658), .Y(n48648) );
  NAND4X1 U54175 ( .A(n18565), .B(n48653), .C(n48652), .D(n48651), .Y(n36361)
         );
  NAND2X1 U54176 ( .A(n43004), .B(n48662), .Y(n48652) );
  NAND4X1 U54177 ( .A(n18541), .B(n48657), .C(n48656), .D(n48655), .Y(n36353)
         );
  NAND2X1 U54178 ( .A(n43002), .B(n48666), .Y(n48656) );
  NAND4X1 U54179 ( .A(n18517), .B(n48661), .C(n48660), .D(n48659), .Y(n36345)
         );
  NAND2X1 U54180 ( .A(n43007), .B(n48670), .Y(n48660) );
  NAND4X1 U54181 ( .A(n18493), .B(n48665), .C(n48664), .D(n48663), .Y(n36337)
         );
  NAND2X1 U54182 ( .A(n43008), .B(n48674), .Y(n48664) );
  NAND4X1 U54183 ( .A(n18469), .B(n48669), .C(n48668), .D(n48667), .Y(n36329)
         );
  NAND2X1 U54184 ( .A(n42994), .B(n48678), .Y(n48668) );
  NAND4X1 U54185 ( .A(n18445), .B(n48673), .C(n48672), .D(n48671), .Y(n36321)
         );
  NAND2X1 U54186 ( .A(n43001), .B(n48682), .Y(n48672) );
  NAND4X1 U54187 ( .A(n18421), .B(n48677), .C(n48676), .D(n48675), .Y(n36313)
         );
  NAND2X1 U54188 ( .A(n42997), .B(n48686), .Y(n48676) );
  NAND4X1 U54189 ( .A(n18397), .B(n48681), .C(n48680), .D(n48679), .Y(n36305)
         );
  NAND2X1 U54190 ( .A(n42998), .B(n48690), .Y(n48680) );
  NAND4X1 U54191 ( .A(n18373), .B(n48685), .C(n48684), .D(n48683), .Y(n36297)
         );
  NAND2X1 U54192 ( .A(n42998), .B(n48694), .Y(n48684) );
  NAND4X1 U54193 ( .A(n18259), .B(n49019), .C(n49018), .D(n49017), .Y(n36259)
         );
  NAND2X1 U54194 ( .A(n42992), .B(n51010), .Y(n49018) );
  NAND4X1 U54195 ( .A(n19153), .B(n49028), .C(n49027), .D(n49026), .Y(n36557)
         );
  NAND4X1 U54196 ( .A(n19129), .B(n49032), .C(n49031), .D(n49030), .Y(n36549)
         );
  NAND4X1 U54197 ( .A(n19105), .B(n49035), .C(n49034), .D(n49033), .Y(n36541)
         );
  NAND4X1 U54198 ( .A(n19081), .B(n49038), .C(n49037), .D(n49036), .Y(n36533)
         );
  NAND4X1 U54199 ( .A(n19057), .B(n49042), .C(n49041), .D(n49040), .Y(n36525)
         );
  NAND4X1 U54200 ( .A(n19033), .B(n49046), .C(n49045), .D(n49044), .Y(n36517)
         );
  NAND4X1 U54201 ( .A(n19009), .B(n49050), .C(n49049), .D(n49048), .Y(n36509)
         );
  NAND4X1 U54202 ( .A(n18985), .B(n49054), .C(n49053), .D(n49052), .Y(n36501)
         );
  NAND4X1 U54203 ( .A(n18961), .B(n49057), .C(n49056), .D(n49055), .Y(n36493)
         );
  NAND2X1 U54204 ( .A(n43008), .B(n49066), .Y(n49056) );
  NAND4X1 U54205 ( .A(n18937), .B(n49061), .C(n49060), .D(n49059), .Y(n36485)
         );
  NAND4X1 U54206 ( .A(n18913), .B(n49065), .C(n49064), .D(n49063), .Y(n36477)
         );
  NAND2X1 U54207 ( .A(n43008), .B(n49074), .Y(n49064) );
  NAND4X1 U54208 ( .A(n18889), .B(n49069), .C(n49068), .D(n49067), .Y(n36469)
         );
  NAND2X1 U54209 ( .A(n43008), .B(n49078), .Y(n49068) );
  NAND4X1 U54210 ( .A(n18865), .B(n49073), .C(n49072), .D(n49071), .Y(n36461)
         );
  NAND2X1 U54211 ( .A(n43008), .B(n49082), .Y(n49072) );
  NAND4X1 U54212 ( .A(n18841), .B(n49077), .C(n49076), .D(n49075), .Y(n36453)
         );
  NAND2X1 U54213 ( .A(n43008), .B(n49086), .Y(n49076) );
  NAND4X1 U54214 ( .A(n18817), .B(n49081), .C(n49080), .D(n49079), .Y(n36445)
         );
  NAND2X1 U54215 ( .A(n43008), .B(n49090), .Y(n49080) );
  NAND4X1 U54216 ( .A(n18793), .B(n49085), .C(n49084), .D(n49083), .Y(n36437)
         );
  NAND2X1 U54217 ( .A(n43008), .B(n49094), .Y(n49084) );
  NAND4X1 U54218 ( .A(n18769), .B(n49089), .C(n49088), .D(n49087), .Y(n36429)
         );
  NAND2X1 U54219 ( .A(n43008), .B(n49098), .Y(n49088) );
  NAND4X1 U54220 ( .A(n18745), .B(n49093), .C(n49092), .D(n49091), .Y(n36421)
         );
  NAND2X1 U54221 ( .A(n43008), .B(n49102), .Y(n49092) );
  NAND4X1 U54222 ( .A(n18721), .B(n49097), .C(n49096), .D(n49095), .Y(n36413)
         );
  NAND2X1 U54223 ( .A(n43008), .B(n49106), .Y(n49096) );
  NAND4X1 U54224 ( .A(n18697), .B(n49101), .C(n49100), .D(n49099), .Y(n36405)
         );
  NAND2X1 U54225 ( .A(n43008), .B(n49110), .Y(n49100) );
  NAND4X1 U54226 ( .A(n18673), .B(n49105), .C(n49104), .D(n49103), .Y(n36397)
         );
  NAND2X1 U54227 ( .A(n43007), .B(n49114), .Y(n49104) );
  NAND4X1 U54228 ( .A(n18649), .B(n49109), .C(n49108), .D(n49107), .Y(n36389)
         );
  NAND2X1 U54229 ( .A(n43008), .B(n49118), .Y(n49108) );
  NAND4X1 U54230 ( .A(n18625), .B(n49113), .C(n49112), .D(n49111), .Y(n36381)
         );
  NAND2X1 U54231 ( .A(n43007), .B(n49122), .Y(n49112) );
  NAND4X1 U54232 ( .A(n18601), .B(n49117), .C(n49116), .D(n49115), .Y(n36373)
         );
  NAND2X1 U54233 ( .A(n43008), .B(n49126), .Y(n49116) );
  NAND4X1 U54234 ( .A(n18577), .B(n49121), .C(n49120), .D(n49119), .Y(n36365)
         );
  NAND2X1 U54235 ( .A(n43007), .B(n49130), .Y(n49120) );
  NAND4X1 U54236 ( .A(n18553), .B(n49125), .C(n49124), .D(n49123), .Y(n36357)
         );
  NAND2X1 U54237 ( .A(n43007), .B(n41231), .Y(n49124) );
  NAND4X1 U54238 ( .A(n18529), .B(n49129), .C(n49128), .D(n49127), .Y(n36349)
         );
  NAND2X1 U54239 ( .A(n43007), .B(n49137), .Y(n49128) );
  NAND4X1 U54240 ( .A(n18505), .B(n49133), .C(n49132), .D(n49131), .Y(n36341)
         );
  NAND2X1 U54241 ( .A(n43007), .B(n49141), .Y(n49132) );
  NAND4X1 U54242 ( .A(n18481), .B(n49136), .C(n49135), .D(n49134), .Y(n36333)
         );
  NAND2X1 U54243 ( .A(n43007), .B(n41259), .Y(n49135) );
  NAND4X1 U54244 ( .A(n18457), .B(n49140), .C(n49139), .D(n49138), .Y(n36325)
         );
  NAND2X1 U54245 ( .A(n43007), .B(n49148), .Y(n49139) );
  NAND4X1 U54246 ( .A(n18433), .B(n49144), .C(n49143), .D(n49142), .Y(n36317)
         );
  NAND2X1 U54247 ( .A(n43007), .B(n49152), .Y(n49143) );
  NAND4X1 U54248 ( .A(n18409), .B(n49147), .C(n49146), .D(n49145), .Y(n36309)
         );
  NAND2X1 U54249 ( .A(n43007), .B(n49156), .Y(n49146) );
  NAND4X1 U54250 ( .A(n18385), .B(n49151), .C(n49150), .D(n49149), .Y(n36301)
         );
  NAND2X1 U54251 ( .A(n43007), .B(n49160), .Y(n49150) );
  NAND4X1 U54252 ( .A(n18361), .B(n49155), .C(n49154), .D(n49153), .Y(n36293)
         );
  NAND2X1 U54253 ( .A(n43007), .B(n49164), .Y(n49154) );
  NAND4X1 U54254 ( .A(n18337), .B(n49159), .C(n49158), .D(n49157), .Y(n36285)
         );
  NAND2X1 U54255 ( .A(n43007), .B(n37541), .Y(n49158) );
  NAND4X1 U54256 ( .A(n18313), .B(n49163), .C(n49162), .D(n49161), .Y(n36277)
         );
  NAND2X1 U54257 ( .A(n43006), .B(n49171), .Y(n49162) );
  NAND4X1 U54258 ( .A(n18289), .B(n49167), .C(n49166), .D(n49165), .Y(n36269)
         );
  NAND4X1 U54259 ( .A(n18265), .B(n49170), .C(n49169), .D(n49168), .Y(n36261)
         );
  NAND2X1 U54260 ( .A(n43006), .B(n50796), .Y(n49169) );
  NAND4X1 U54261 ( .A(n18241), .B(n49174), .C(n49173), .D(n49172), .Y(n36253)
         );
  NAND2X1 U54262 ( .A(n43006), .B(n50795), .Y(n49173) );
  NAND4X1 U54263 ( .A(n19132), .B(n49184), .C(n49183), .D(n49182), .Y(n36550)
         );
  NAND2X1 U54264 ( .A(n43006), .B(n49192), .Y(n49183) );
  NAND4X1 U54265 ( .A(n19108), .B(n49188), .C(n49187), .D(n49186), .Y(n36542)
         );
  NAND2X1 U54266 ( .A(n43006), .B(n49196), .Y(n49187) );
  NAND4X1 U54267 ( .A(n19084), .B(n49191), .C(n49190), .D(n49189), .Y(n36534)
         );
  NAND2X1 U54268 ( .A(n43006), .B(n49200), .Y(n49190) );
  NAND4X1 U54269 ( .A(n19060), .B(n49195), .C(n49194), .D(n49193), .Y(n36526)
         );
  NAND2X1 U54270 ( .A(n43006), .B(n49204), .Y(n49194) );
  NAND4X1 U54271 ( .A(n19036), .B(n49199), .C(n49198), .D(n49197), .Y(n36518)
         );
  NAND2X1 U54272 ( .A(n43006), .B(n49208), .Y(n49198) );
  NAND4X1 U54273 ( .A(n19012), .B(n49203), .C(n49202), .D(n49201), .Y(n36510)
         );
  NAND2X1 U54274 ( .A(n43006), .B(n49212), .Y(n49202) );
  NAND4X1 U54275 ( .A(n18988), .B(n49207), .C(n49206), .D(n49205), .Y(n36502)
         );
  NAND2X1 U54276 ( .A(n43005), .B(n49216), .Y(n49206) );
  NAND4X1 U54277 ( .A(n18964), .B(n49211), .C(n49210), .D(n49209), .Y(n36494)
         );
  NAND2X1 U54278 ( .A(n43006), .B(n49220), .Y(n49210) );
  NAND4X1 U54279 ( .A(n18940), .B(n49215), .C(n49214), .D(n49213), .Y(n36486)
         );
  NAND2X1 U54280 ( .A(n43005), .B(n49224), .Y(n49214) );
  NAND4X1 U54281 ( .A(n18916), .B(n49219), .C(n49218), .D(n49217), .Y(n36478)
         );
  NAND2X1 U54282 ( .A(n43005), .B(n49228), .Y(n49218) );
  NAND4X1 U54283 ( .A(n18892), .B(n49223), .C(n49222), .D(n49221), .Y(n36470)
         );
  NAND2X1 U54284 ( .A(n43005), .B(n49232), .Y(n49222) );
  NAND4X1 U54285 ( .A(n18868), .B(n49227), .C(n49226), .D(n49225), .Y(n36462)
         );
  NAND2X1 U54286 ( .A(n43005), .B(n49236), .Y(n49226) );
  NAND4X1 U54287 ( .A(n18844), .B(n49231), .C(n49230), .D(n49229), .Y(n36454)
         );
  NAND2X1 U54288 ( .A(n43005), .B(n49240), .Y(n49230) );
  NAND4X1 U54289 ( .A(n18820), .B(n49235), .C(n49234), .D(n49233), .Y(n36446)
         );
  NAND2X1 U54290 ( .A(n43005), .B(n49244), .Y(n49234) );
  NAND4X1 U54291 ( .A(n18796), .B(n49239), .C(n49238), .D(n49237), .Y(n36438)
         );
  NAND2X1 U54292 ( .A(n43005), .B(n49248), .Y(n49238) );
  NAND4X1 U54293 ( .A(n18772), .B(n49243), .C(n49242), .D(n49241), .Y(n36430)
         );
  NAND2X1 U54294 ( .A(n43005), .B(n49252), .Y(n49242) );
  NAND4X1 U54295 ( .A(n18748), .B(n49247), .C(n49246), .D(n49245), .Y(n36422)
         );
  NAND2X1 U54296 ( .A(n43005), .B(n49256), .Y(n49246) );
  NAND4X1 U54297 ( .A(n18724), .B(n49251), .C(n49250), .D(n49249), .Y(n36414)
         );
  NAND2X1 U54298 ( .A(n43005), .B(n49260), .Y(n49250) );
  NAND4X1 U54299 ( .A(n18700), .B(n49255), .C(n49254), .D(n49253), .Y(n36406)
         );
  NAND2X1 U54300 ( .A(n43005), .B(n49264), .Y(n49254) );
  NAND4X1 U54301 ( .A(n18676), .B(n49259), .C(n49258), .D(n49257), .Y(n36398)
         );
  NAND2X1 U54302 ( .A(n43004), .B(n49268), .Y(n49258) );
  NAND4X1 U54303 ( .A(n18652), .B(n49263), .C(n49262), .D(n49261), .Y(n36390)
         );
  NAND2X1 U54304 ( .A(n43004), .B(n49272), .Y(n49262) );
  NAND4X1 U54305 ( .A(n18628), .B(n49267), .C(n49266), .D(n49265), .Y(n36382)
         );
  NAND2X1 U54306 ( .A(n43004), .B(n49276), .Y(n49266) );
  NAND4X1 U54307 ( .A(n18604), .B(n49271), .C(n49270), .D(n49269), .Y(n36374)
         );
  NAND2X1 U54308 ( .A(n43004), .B(n49280), .Y(n49270) );
  NAND4X1 U54309 ( .A(n18580), .B(n49275), .C(n49274), .D(n49273), .Y(n36366)
         );
  NAND2X1 U54310 ( .A(n43004), .B(n49284), .Y(n49274) );
  NAND4X1 U54311 ( .A(n18556), .B(n49279), .C(n49278), .D(n49277), .Y(n36358)
         );
  NAND2X1 U54312 ( .A(n43004), .B(n49288), .Y(n49278) );
  NAND4X1 U54313 ( .A(n18532), .B(n49283), .C(n49282), .D(n49281), .Y(n36350)
         );
  NAND2X1 U54314 ( .A(n43004), .B(n41227), .Y(n49282) );
  NAND4X1 U54315 ( .A(n18508), .B(n49287), .C(n49286), .D(n49285), .Y(n36342)
         );
  NAND2X1 U54316 ( .A(n43004), .B(n49295), .Y(n49286) );
  NAND4X1 U54317 ( .A(n18484), .B(n49291), .C(n49290), .D(n49289), .Y(n36334)
         );
  NAND2X1 U54318 ( .A(n43004), .B(n49299), .Y(n49290) );
  NAND4X1 U54319 ( .A(n18460), .B(n49294), .C(n49293), .D(n49292), .Y(n36326)
         );
  NAND2X1 U54320 ( .A(n43004), .B(n49303), .Y(n49293) );
  NAND4X1 U54321 ( .A(n18436), .B(n49298), .C(n49297), .D(n49296), .Y(n36318)
         );
  NAND2X1 U54322 ( .A(n43004), .B(n49307), .Y(n49297) );
  NAND4X1 U54323 ( .A(n18412), .B(n49302), .C(n49301), .D(n49300), .Y(n36310)
         );
  NAND2X1 U54324 ( .A(n43004), .B(n49311), .Y(n49301) );
  NAND4X1 U54325 ( .A(n18388), .B(n49306), .C(n49305), .D(n49304), .Y(n36302)
         );
  NAND2X1 U54326 ( .A(n43004), .B(n49315), .Y(n49305) );
  NAND4X1 U54327 ( .A(n18364), .B(n49310), .C(n49309), .D(n49308), .Y(n36294)
         );
  NAND2X1 U54328 ( .A(n43003), .B(n49319), .Y(n49309) );
  NAND4X1 U54329 ( .A(n18340), .B(n49314), .C(n49313), .D(n49312), .Y(n36286)
         );
  NAND2X1 U54330 ( .A(n43003), .B(n37542), .Y(n49313) );
  NAND4X1 U54331 ( .A(n18316), .B(n49318), .C(n49317), .D(n49316), .Y(n36278)
         );
  NAND2X1 U54332 ( .A(n43003), .B(n37543), .Y(n49317) );
  NAND4X1 U54333 ( .A(n18292), .B(n49322), .C(n49321), .D(n49320), .Y(n36270)
         );
  NAND4X1 U54334 ( .A(n18268), .B(n49325), .C(n49324), .D(n49323), .Y(n36262)
         );
  NAND4X1 U54335 ( .A(n18244), .B(n49329), .C(n49328), .D(n49327), .Y(n36254)
         );
  NAND2X1 U54336 ( .A(n43003), .B(n49326), .Y(n49328) );
  NAND4X1 U54337 ( .A(n19135), .B(n49339), .C(n49338), .D(n49337), .Y(n36551)
         );
  NAND2X1 U54338 ( .A(n43003), .B(n49347), .Y(n49338) );
  NAND4X1 U54339 ( .A(n19111), .B(n49343), .C(n49342), .D(n49341), .Y(n36543)
         );
  NAND2X1 U54340 ( .A(n43003), .B(n49351), .Y(n49342) );
  NAND4X1 U54341 ( .A(n19087), .B(n49346), .C(n49345), .D(n49344), .Y(n36535)
         );
  NAND2X1 U54342 ( .A(n43003), .B(n49355), .Y(n49345) );
  NAND4X1 U54343 ( .A(n19063), .B(n49350), .C(n49349), .D(n49348), .Y(n36527)
         );
  NAND2X1 U54344 ( .A(n43003), .B(n49359), .Y(n49349) );
  NAND4X1 U54345 ( .A(n19039), .B(n49354), .C(n49353), .D(n49352), .Y(n36519)
         );
  NAND2X1 U54346 ( .A(n43003), .B(n49363), .Y(n49353) );
  NAND4X1 U54347 ( .A(n19015), .B(n49358), .C(n49357), .D(n49356), .Y(n36511)
         );
  NAND2X1 U54348 ( .A(n43002), .B(n49367), .Y(n49357) );
  NAND4X1 U54349 ( .A(n18991), .B(n49362), .C(n49361), .D(n49360), .Y(n36503)
         );
  NAND2X1 U54350 ( .A(n43002), .B(n49371), .Y(n49361) );
  NAND4X1 U54351 ( .A(n18967), .B(n49366), .C(n49365), .D(n49364), .Y(n36495)
         );
  NAND2X1 U54352 ( .A(n43002), .B(n49375), .Y(n49365) );
  NAND4X1 U54353 ( .A(n18943), .B(n49370), .C(n49369), .D(n49368), .Y(n36487)
         );
  NAND2X1 U54354 ( .A(n43002), .B(n49379), .Y(n49369) );
  NAND4X1 U54355 ( .A(n18919), .B(n49374), .C(n49373), .D(n49372), .Y(n36479)
         );
  NAND2X1 U54356 ( .A(n43002), .B(n49383), .Y(n49373) );
  NAND4X1 U54357 ( .A(n18895), .B(n49378), .C(n49377), .D(n49376), .Y(n36471)
         );
  NAND2X1 U54358 ( .A(n43002), .B(n49387), .Y(n49377) );
  NAND4X1 U54359 ( .A(n18871), .B(n49382), .C(n49381), .D(n49380), .Y(n36463)
         );
  NAND2X1 U54360 ( .A(n43002), .B(n49391), .Y(n49381) );
  NAND4X1 U54361 ( .A(n18847), .B(n49386), .C(n49385), .D(n49384), .Y(n36455)
         );
  NAND2X1 U54362 ( .A(n43002), .B(n49395), .Y(n49385) );
  NAND4X1 U54363 ( .A(n18823), .B(n49390), .C(n49389), .D(n49388), .Y(n36447)
         );
  NAND2X1 U54364 ( .A(n43005), .B(n49399), .Y(n49389) );
  NAND4X1 U54365 ( .A(n18799), .B(n49394), .C(n49393), .D(n49392), .Y(n36439)
         );
  NAND2X1 U54366 ( .A(n43002), .B(n49403), .Y(n49393) );
  NAND4X1 U54367 ( .A(n18775), .B(n49398), .C(n49397), .D(n49396), .Y(n36431)
         );
  NAND2X1 U54368 ( .A(n43002), .B(n49407), .Y(n49397) );
  NAND4X1 U54369 ( .A(n18751), .B(n49402), .C(n49401), .D(n49400), .Y(n36423)
         );
  NAND2X1 U54370 ( .A(n43002), .B(n49411), .Y(n49401) );
  NAND4X1 U54371 ( .A(n18727), .B(n49406), .C(n49405), .D(n49404), .Y(n36415)
         );
  NAND2X1 U54372 ( .A(n43002), .B(n49415), .Y(n49405) );
  NAND4X1 U54373 ( .A(n18703), .B(n49410), .C(n49409), .D(n49408), .Y(n36407)
         );
  NAND2X1 U54374 ( .A(n43002), .B(n49419), .Y(n49409) );
  NAND4X1 U54375 ( .A(n18679), .B(n49414), .C(n49413), .D(n49412), .Y(n36399)
         );
  NAND2X1 U54376 ( .A(n43001), .B(n49423), .Y(n49413) );
  NAND4X1 U54377 ( .A(n18655), .B(n49418), .C(n49417), .D(n49416), .Y(n36391)
         );
  NAND2X1 U54378 ( .A(n43001), .B(n41221), .Y(n49417) );
  NAND4X1 U54379 ( .A(n18631), .B(n49422), .C(n49421), .D(n49420), .Y(n36383)
         );
  NAND2X1 U54380 ( .A(n43001), .B(n49430), .Y(n49421) );
  NAND4X1 U54381 ( .A(n18607), .B(n49426), .C(n49425), .D(n49424), .Y(n36375)
         );
  NAND2X1 U54382 ( .A(n43001), .B(n49434), .Y(n49425) );
  NAND4X1 U54383 ( .A(n18583), .B(n49429), .C(n49428), .D(n49427), .Y(n36367)
         );
  NAND2X1 U54384 ( .A(n43001), .B(n49438), .Y(n49428) );
  NAND4X1 U54385 ( .A(n18559), .B(n49433), .C(n49432), .D(n49431), .Y(n36359)
         );
  NAND2X1 U54386 ( .A(n43001), .B(n49442), .Y(n49432) );
  NAND4X1 U54387 ( .A(n18535), .B(n49437), .C(n49436), .D(n49435), .Y(n36351)
         );
  NAND2X1 U54388 ( .A(n43001), .B(n49446), .Y(n49436) );
  NAND4X1 U54389 ( .A(n18511), .B(n49441), .C(n49440), .D(n49439), .Y(n36343)
         );
  NAND2X1 U54390 ( .A(n43001), .B(n49450), .Y(n49440) );
  NAND4X1 U54391 ( .A(n18487), .B(n49445), .C(n49444), .D(n49443), .Y(n36335)
         );
  NAND2X1 U54392 ( .A(n43001), .B(n49454), .Y(n49444) );
  NAND4X1 U54393 ( .A(n18463), .B(n49449), .C(n49448), .D(n49447), .Y(n36327)
         );
  NAND2X1 U54394 ( .A(n43001), .B(n49458), .Y(n49448) );
  NAND4X1 U54395 ( .A(n18439), .B(n49453), .C(n49452), .D(n49451), .Y(n36319)
         );
  NAND2X1 U54396 ( .A(n43001), .B(n49462), .Y(n49452) );
  NAND4X1 U54397 ( .A(n18415), .B(n49457), .C(n49456), .D(n49455), .Y(n36311)
         );
  NAND2X1 U54398 ( .A(n43001), .B(n49466), .Y(n49456) );
  NAND4X1 U54399 ( .A(n18391), .B(n49461), .C(n49460), .D(n49459), .Y(n36303)
         );
  NAND2X1 U54400 ( .A(n43001), .B(n49470), .Y(n49460) );
  NAND4X1 U54401 ( .A(n18367), .B(n49465), .C(n49464), .D(n49463), .Y(n36295)
         );
  NAND2X1 U54402 ( .A(n43000), .B(n49474), .Y(n49464) );
  NAND4X1 U54403 ( .A(n18343), .B(n49469), .C(n49468), .D(n49467), .Y(n36287)
         );
  NAND2X1 U54404 ( .A(n43000), .B(n49478), .Y(n49468) );
  NAND4X1 U54405 ( .A(n18319), .B(n49473), .C(n49472), .D(n49471), .Y(n36279)
         );
  NAND2X1 U54406 ( .A(n43000), .B(n37195), .Y(n49472) );
  NAND4X1 U54407 ( .A(n18295), .B(n49477), .C(n49476), .D(n49475), .Y(n36271)
         );
  NAND4X1 U54408 ( .A(n18271), .B(n49481), .C(n49480), .D(n49479), .Y(n36263)
         );
  NAND2X1 U54409 ( .A(n43000), .B(n50379), .Y(n49480) );
  NAND4X1 U54410 ( .A(n18247), .B(n49484), .C(n49483), .D(n49482), .Y(n36255)
         );
  NAND2X1 U54411 ( .A(n43000), .B(n50378), .Y(n49483) );
  NAND4X1 U54412 ( .A(n18349), .B(n48689), .C(n48688), .D(n48687), .Y(n36289)
         );
  NAND2X1 U54413 ( .A(n42998), .B(n48698), .Y(n48688) );
  NAND4X1 U54414 ( .A(n18325), .B(n48693), .C(n48692), .D(n48691), .Y(n36281)
         );
  NAND2X1 U54415 ( .A(n42998), .B(n37544), .Y(n48692) );
  NAND4X1 U54416 ( .A(n18301), .B(n48697), .C(n48696), .D(n48695), .Y(n36273)
         );
  NAND2X1 U54417 ( .A(n42998), .B(n48705), .Y(n48696) );
  NAND4X1 U54418 ( .A(n18277), .B(n48701), .C(n48700), .D(n48699), .Y(n36265)
         );
  NAND2X1 U54419 ( .A(n42998), .B(n51438), .Y(n48700) );
  NAND4X1 U54420 ( .A(n18253), .B(n48704), .C(n48703), .D(n48702), .Y(n36257)
         );
  NAND2X1 U54421 ( .A(n42998), .B(n51437), .Y(n48703) );
  NAND4X1 U54422 ( .A(n18229), .B(n48708), .C(n48707), .D(n48706), .Y(n36249)
         );
  NAND2X1 U54423 ( .A(n42998), .B(n37540), .Y(n48707) );
  AOI2BB2X1 U54424 ( .B0(net265530), .B1(n48705), .A0N(n40281), .A1N(n34108),
        .Y(n48706) );
  NAND4X1 U54425 ( .A(n19144), .B(n48719), .C(n48718), .D(n48717), .Y(n36554)
         );
  NAND2X1 U54426 ( .A(n42998), .B(n48726), .Y(n48718) );
  NAND4X1 U54427 ( .A(n19120), .B(n48722), .C(n48721), .D(n48720), .Y(n36546)
         );
  NAND2X1 U54428 ( .A(n42998), .B(n48730), .Y(n48721) );
  NAND4X1 U54429 ( .A(n19096), .B(n48725), .C(n48724), .D(n48723), .Y(n36538)
         );
  NAND2X1 U54430 ( .A(n42998), .B(n48734), .Y(n48724) );
  NAND4X1 U54431 ( .A(n19072), .B(n48729), .C(n48728), .D(n48727), .Y(n36530)
         );
  NAND2X1 U54432 ( .A(n42998), .B(n48738), .Y(n48728) );
  NAND4X1 U54433 ( .A(n19048), .B(n48733), .C(n48732), .D(n48731), .Y(n36522)
         );
  NAND2X1 U54434 ( .A(n42997), .B(n48742), .Y(n48732) );
  NAND4X1 U54435 ( .A(n19024), .B(n48737), .C(n48736), .D(n48735), .Y(n36514)
         );
  NAND2X1 U54436 ( .A(n42997), .B(n48746), .Y(n48736) );
  NAND4X1 U54437 ( .A(n19000), .B(n48741), .C(n48740), .D(n48739), .Y(n36506)
         );
  NAND2X1 U54438 ( .A(n42997), .B(n48750), .Y(n48740) );
  NAND4X1 U54439 ( .A(n18976), .B(n48745), .C(n48744), .D(n48743), .Y(n36498)
         );
  NAND2X1 U54440 ( .A(n42997), .B(n48754), .Y(n48744) );
  NAND4X1 U54441 ( .A(n18952), .B(n48749), .C(n48748), .D(n48747), .Y(n36490)
         );
  NAND2X1 U54442 ( .A(n42997), .B(n48758), .Y(n48748) );
  NAND4X1 U54443 ( .A(n18928), .B(n48753), .C(n48752), .D(n48751), .Y(n36482)
         );
  NAND2X1 U54444 ( .A(n42997), .B(n48762), .Y(n48752) );
  NAND4X1 U54445 ( .A(n18904), .B(n48757), .C(n48756), .D(n48755), .Y(n36474)
         );
  NAND2X1 U54446 ( .A(n42997), .B(n48766), .Y(n48756) );
  NAND4X1 U54447 ( .A(n18880), .B(n48761), .C(n48760), .D(n48759), .Y(n36466)
         );
  NAND2X1 U54448 ( .A(n42997), .B(n48770), .Y(n48760) );
  NAND4X1 U54449 ( .A(n18856), .B(n48765), .C(n48764), .D(n48763), .Y(n36458)
         );
  NAND2X1 U54450 ( .A(n42997), .B(n48774), .Y(n48764) );
  NAND4X1 U54451 ( .A(n18832), .B(n48769), .C(n48768), .D(n48767), .Y(n36450)
         );
  NAND2X1 U54452 ( .A(n42997), .B(n48778), .Y(n48768) );
  NAND4X1 U54453 ( .A(n18808), .B(n48773), .C(n48772), .D(n48771), .Y(n36442)
         );
  NAND2X1 U54454 ( .A(n43000), .B(n48782), .Y(n48772) );
  NAND4X1 U54455 ( .A(n18784), .B(n48777), .C(n48776), .D(n48775), .Y(n36434)
         );
  NAND2X1 U54456 ( .A(n42997), .B(n48786), .Y(n48776) );
  NAND4X1 U54457 ( .A(n18760), .B(n48781), .C(n48780), .D(n48779), .Y(n36426)
         );
  NAND2X1 U54458 ( .A(n42997), .B(n48790), .Y(n48780) );
  NAND4X1 U54459 ( .A(n18736), .B(n48785), .C(n48784), .D(n48783), .Y(n36418)
         );
  NAND2X1 U54460 ( .A(n42997), .B(n48794), .Y(n48784) );
  NAND4X1 U54461 ( .A(n18712), .B(n48789), .C(n48788), .D(n48787), .Y(n36410)
         );
  NAND2X1 U54462 ( .A(n42996), .B(n48798), .Y(n48788) );
  NAND4X1 U54463 ( .A(n18688), .B(n48793), .C(n48792), .D(n48791), .Y(n36402)
         );
  NAND2X1 U54464 ( .A(n42996), .B(n48802), .Y(n48792) );
  NAND4X1 U54465 ( .A(n18664), .B(n48797), .C(n48796), .D(n48795), .Y(n36394)
         );
  NAND2X1 U54466 ( .A(n42996), .B(n48806), .Y(n48796) );
  NAND4X1 U54467 ( .A(n18640), .B(n48801), .C(n48800), .D(n48799), .Y(n36386)
         );
  NAND2X1 U54468 ( .A(n42996), .B(n48810), .Y(n48800) );
  NAND4X1 U54469 ( .A(n18616), .B(n48805), .C(n48804), .D(n48803), .Y(n36378)
         );
  NAND2X1 U54470 ( .A(n42996), .B(n48814), .Y(n48804) );
  NAND4X1 U54471 ( .A(n18592), .B(n48809), .C(n48808), .D(n48807), .Y(n36370)
         );
  NAND2X1 U54472 ( .A(n42996), .B(n48818), .Y(n48808) );
  NAND4X1 U54473 ( .A(n18568), .B(n48813), .C(n48812), .D(n48811), .Y(n36362)
         );
  NAND2X1 U54474 ( .A(n42996), .B(n48822), .Y(n48812) );
  NAND4X1 U54475 ( .A(n18544), .B(n48817), .C(n48816), .D(n48815), .Y(n36354)
         );
  NAND2X1 U54476 ( .A(n42996), .B(n48826), .Y(n48816) );
  NAND4X1 U54477 ( .A(n18520), .B(n48821), .C(n48820), .D(n48819), .Y(n36346)
         );
  NAND2X1 U54478 ( .A(n42996), .B(n48830), .Y(n48820) );
  NAND4X1 U54479 ( .A(n18496), .B(n48825), .C(n48824), .D(n48823), .Y(n36338)
         );
  NAND2X1 U54480 ( .A(n42996), .B(n48834), .Y(n48824) );
  NAND4X1 U54481 ( .A(n18472), .B(n48829), .C(n48828), .D(n48827), .Y(n36330)
         );
  NAND2X1 U54482 ( .A(n42996), .B(n48838), .Y(n48828) );
  NAND4X1 U54483 ( .A(n18448), .B(n48833), .C(n48832), .D(n48831), .Y(n36322)
         );
  NAND2X1 U54484 ( .A(n42996), .B(n48842), .Y(n48832) );
  NAND4X1 U54485 ( .A(n18424), .B(n48837), .C(n48836), .D(n48835), .Y(n36314)
         );
  NAND2X1 U54486 ( .A(n42995), .B(n48846), .Y(n48836) );
  NAND4X1 U54487 ( .A(n18400), .B(n48841), .C(n48840), .D(n48839), .Y(n36306)
         );
  NAND2X1 U54488 ( .A(n42995), .B(n48850), .Y(n48840) );
  NAND4X1 U54489 ( .A(n18376), .B(n48845), .C(n48844), .D(n48843), .Y(n36298)
         );
  NAND2X1 U54490 ( .A(n42995), .B(n48854), .Y(n48844) );
  NAND4X1 U54491 ( .A(n18352), .B(n48849), .C(n48848), .D(n48847), .Y(n36290)
         );
  NAND2X1 U54492 ( .A(n42995), .B(n37545), .Y(n48848) );
  NAND4X1 U54493 ( .A(n18328), .B(n48853), .C(n48852), .D(n48851), .Y(n36282)
         );
  NAND2X1 U54494 ( .A(n42995), .B(n37546), .Y(n48852) );
  NAND4X1 U54495 ( .A(n18304), .B(n48857), .C(n48856), .D(n48855), .Y(n36274)
         );
  NAND2X1 U54496 ( .A(n42995), .B(n48864), .Y(n48856) );
  NAND4X1 U54497 ( .A(n18280), .B(n48860), .C(n48859), .D(n48858), .Y(n36266)
         );
  NAND4X1 U54498 ( .A(n18256), .B(n48863), .C(n48862), .D(n48861), .Y(n36258)
         );
  NAND2X1 U54499 ( .A(n42995), .B(n51224), .Y(n48862) );
  NAND4X1 U54500 ( .A(n18232), .B(n48867), .C(n48866), .D(n48865), .Y(n36250)
         );
  NAND2X1 U54501 ( .A(n42995), .B(n51223), .Y(n48866) );
  NAND4X1 U54502 ( .A(n19147), .B(n48877), .C(n48876), .D(n48875), .Y(n36555)
         );
  NAND2X1 U54503 ( .A(n42995), .B(n48884), .Y(n48876) );
  NAND4X1 U54504 ( .A(n19123), .B(n48880), .C(n48879), .D(n48878), .Y(n36547)
         );
  NAND2X1 U54505 ( .A(n42995), .B(n41367), .Y(n48879) );
  NAND4X1 U54506 ( .A(n19099), .B(n48883), .C(n48882), .D(n48881), .Y(n36539)
         );
  NAND2X1 U54507 ( .A(n42994), .B(n48891), .Y(n48882) );
  NAND4X1 U54508 ( .A(n19075), .B(n48887), .C(n48886), .D(n48885), .Y(n36531)
         );
  NAND2X1 U54509 ( .A(n42994), .B(n48895), .Y(n48886) );
  NAND4X1 U54510 ( .A(n19051), .B(n48890), .C(n48889), .D(n48888), .Y(n36523)
         );
  NAND2X1 U54511 ( .A(n42994), .B(n41655), .Y(n48889) );
  NAND4X1 U54512 ( .A(n19027), .B(n48894), .C(n48893), .D(n48892), .Y(n36515)
         );
  NAND2X1 U54513 ( .A(n42994), .B(n48902), .Y(n48893) );
  NAND4X1 U54514 ( .A(n19003), .B(n48898), .C(n48897), .D(n48896), .Y(n36507)
         );
  NAND2X1 U54515 ( .A(n42994), .B(n48906), .Y(n48897) );
  NAND4X1 U54516 ( .A(n18979), .B(n48901), .C(n48900), .D(n48899), .Y(n36499)
         );
  NAND2X1 U54517 ( .A(n42994), .B(n48910), .Y(n48900) );
  NAND4X1 U54518 ( .A(n18955), .B(n48905), .C(n48904), .D(n48903), .Y(n36491)
         );
  NAND2X1 U54519 ( .A(n42994), .B(n48914), .Y(n48904) );
  NAND4X1 U54520 ( .A(n18931), .B(n48909), .C(n48908), .D(n48907), .Y(n36483)
         );
  NAND2X1 U54521 ( .A(n42994), .B(n48918), .Y(n48908) );
  NAND4X1 U54522 ( .A(n18907), .B(n48913), .C(n48912), .D(n48911), .Y(n36475)
         );
  NAND2X1 U54523 ( .A(n42994), .B(n48922), .Y(n48912) );
  NAND4X1 U54524 ( .A(n18883), .B(n48917), .C(n48916), .D(n48915), .Y(n36467)
         );
  NAND2X1 U54525 ( .A(n42994), .B(n48926), .Y(n48916) );
  NAND4X1 U54526 ( .A(n18859), .B(n48921), .C(n48920), .D(n48919), .Y(n36459)
         );
  NAND2X1 U54527 ( .A(n42994), .B(n48930), .Y(n48920) );
  NAND4X1 U54528 ( .A(n18835), .B(n48925), .C(n48924), .D(n48923), .Y(n36451)
         );
  NAND2X1 U54529 ( .A(n42994), .B(n48934), .Y(n48924) );
  NAND4X1 U54530 ( .A(n18811), .B(n48929), .C(n48928), .D(n48927), .Y(n36443)
         );
  NAND2X1 U54531 ( .A(n42994), .B(n48938), .Y(n48928) );
  NAND4X1 U54532 ( .A(n18787), .B(n48933), .C(n48932), .D(n48931), .Y(n36435)
         );
  NAND2X1 U54533 ( .A(n42993), .B(n48942), .Y(n48932) );
  NAND4X1 U54534 ( .A(n18763), .B(n48937), .C(n48936), .D(n48935), .Y(n36427)
         );
  NAND2X1 U54535 ( .A(n42993), .B(n48946), .Y(n48936) );
  NAND4X1 U54536 ( .A(n18739), .B(n48941), .C(n48940), .D(n48939), .Y(n36419)
         );
  NAND2X1 U54537 ( .A(n42993), .B(n48950), .Y(n48940) );
  NAND4X1 U54538 ( .A(n18715), .B(n48945), .C(n48944), .D(n48943), .Y(n36411)
         );
  NAND2X1 U54539 ( .A(n42993), .B(n48954), .Y(n48944) );
  NAND4X1 U54540 ( .A(n18691), .B(n48949), .C(n48948), .D(n48947), .Y(n36403)
         );
  NAND2X1 U54541 ( .A(n42993), .B(n48958), .Y(n48948) );
  NAND4X1 U54542 ( .A(n18667), .B(n48953), .C(n48952), .D(n48951), .Y(n36395)
         );
  NAND2X1 U54543 ( .A(n42993), .B(n48962), .Y(n48952) );
  NAND4X1 U54544 ( .A(n18643), .B(n48957), .C(n48956), .D(n48955), .Y(n36387)
         );
  NAND2X1 U54545 ( .A(n42993), .B(n48966), .Y(n48956) );
  NAND4X1 U54546 ( .A(n18619), .B(n48961), .C(n48960), .D(n48959), .Y(n36379)
         );
  NAND2X1 U54547 ( .A(n42993), .B(n48970), .Y(n48960) );
  NAND4X1 U54548 ( .A(n18595), .B(n48965), .C(n48964), .D(n48963), .Y(n36371)
         );
  NAND2X1 U54549 ( .A(n42993), .B(n48974), .Y(n48964) );
  NAND4X1 U54550 ( .A(n18571), .B(n48969), .C(n48968), .D(n48967), .Y(n36363)
         );
  NAND2X1 U54551 ( .A(n42993), .B(n48978), .Y(n48968) );
  NAND4X1 U54552 ( .A(n18547), .B(n48973), .C(n48972), .D(n48971), .Y(n36355)
         );
  NAND2X1 U54553 ( .A(n42993), .B(n48982), .Y(n48972) );
  NAND4X1 U54554 ( .A(n18523), .B(n48977), .C(n48976), .D(n48975), .Y(n36347)
         );
  NAND2X1 U54555 ( .A(n42993), .B(n48986), .Y(n48976) );
  NAND4X1 U54556 ( .A(n18499), .B(n48981), .C(n48980), .D(n48979), .Y(n36339)
         );
  NAND2X1 U54557 ( .A(n42993), .B(n48990), .Y(n48980) );
  NAND4X1 U54558 ( .A(n18475), .B(n48985), .C(n48984), .D(n48983), .Y(n36331)
         );
  NAND2X1 U54559 ( .A(n42992), .B(n48994), .Y(n48984) );
  NAND4X1 U54560 ( .A(n18451), .B(n48989), .C(n48988), .D(n48987), .Y(n36323)
         );
  NAND2X1 U54561 ( .A(n42992), .B(n48998), .Y(n48988) );
  NAND4X1 U54562 ( .A(n18427), .B(n48993), .C(n48992), .D(n48991), .Y(n36315)
         );
  NAND2X1 U54563 ( .A(n42992), .B(n49002), .Y(n48992) );
  NAND4X1 U54564 ( .A(n18403), .B(n48997), .C(n48996), .D(n48995), .Y(n36307)
         );
  NAND2X1 U54565 ( .A(n42992), .B(n49006), .Y(n48996) );
  NAND4X1 U54566 ( .A(n18379), .B(n49001), .C(n49000), .D(n48999), .Y(n36299)
         );
  NAND2X1 U54567 ( .A(n42992), .B(n49010), .Y(n49000) );
  NAND4X1 U54568 ( .A(n18355), .B(n49005), .C(n49004), .D(n49003), .Y(n36291)
         );
  NAND2X1 U54569 ( .A(n42992), .B(n37547), .Y(n49004) );
  NAND4X1 U54570 ( .A(n18331), .B(n49009), .C(n49008), .D(n49007), .Y(n36283)
         );
  NAND2X1 U54571 ( .A(n42992), .B(n37548), .Y(n49008) );
  NAND4X1 U54572 ( .A(n18307), .B(n49013), .C(n49012), .D(n49011), .Y(n36275)
         );
  NAND4X1 U54573 ( .A(n18283), .B(n49016), .C(n49015), .D(n49014), .Y(n36267)
         );
  NOR2X1 U54574 ( .A(n40391), .B(n47797), .Y(net210497) );
  NOR2X1 U54575 ( .A(n12221), .B(n46674), .Y(net212017) );
  NOR2X1 U54576 ( .A(n10906), .B(n46859), .Y(net211768) );
  NOR2X1 U54577 ( .A(net260332), .B(n46615), .Y(net212194) );
  NOR2X1 U54578 ( .A(n12186), .B(n47872), .Y(n47876) );
  NOR2X1 U54579 ( .A(n12604), .B(n45792), .Y(net213215) );
  NOR2X1 U54580 ( .A(net260352), .B(n44377), .Y(net215069) );
  XOR2X1 U54581 ( .A(n32636), .B(n36822), .Y(n44377) );
  NOR2X1 U54582 ( .A(n12213), .B(n46650), .Y(net212099) );
  NOR2X1 U54583 ( .A(n12614), .B(n45560), .Y(net213613) );
  XOR2X1 U54584 ( .A(n32593), .B(n36786), .Y(n45560) );
  NOR2X1 U54585 ( .A(n12424), .B(n43528), .Y(net216202) );
  NOR2X1 U54586 ( .A(n12591), .B(n44330), .Y(n44334) );
  XOR2X1 U54587 ( .A(n32460), .B(n36823), .Y(n44330) );
  NOR2X1 U54588 ( .A(net260367), .B(n43468), .Y(n43472) );
  NOR2X1 U54589 ( .A(net260355), .B(n44372), .Y(net215078) );
  XOR2X1 U54590 ( .A(n32644), .B(n36822), .Y(n44372) );
  NOR2X1 U54591 ( .A(net271431), .B(n45715), .Y(net213317) );
  NOR2X1 U54592 ( .A(net260346), .B(n44350), .Y(net215132) );
  XOR2X1 U54593 ( .A(n32468), .B(n36825), .Y(n44350) );
  NOR2X1 U54594 ( .A(n12427), .B(n44621), .Y(net214683) );
  NOR2X1 U54595 ( .A(n10484), .B(n46087), .Y(net212826) );
  NOR2X1 U54596 ( .A(net260412), .B(n45574), .Y(net213562) );
  NOR2X1 U54597 ( .A(net271999), .B(n45603), .Y(net213477) );
  NOR2X1 U54598 ( .A(net260376), .B(n43512), .Y(net216274) );
  NOR2X1 U54599 ( .A(n12640), .B(n45584), .Y(net213532) );
  XOR2X1 U54600 ( .A(n32897), .B(n36776), .Y(n45584) );
  NOR2X1 U54601 ( .A(net260403), .B(n45552), .Y(net213633) );
  XOR2X1 U54602 ( .A(n32641), .B(n36786), .Y(n45552) );
  NOR2X1 U54603 ( .A(net271996), .B(n45612), .Y(n45616) );
  NOR2X1 U54604 ( .A(n12433), .B(n43500), .Y(net216310) );
  NOR2X1 U54605 ( .A(n12210), .B(n46651), .Y(net212094) );
  NOR2X1 U54606 ( .A(n12219), .B(n46665), .Y(net212043) );
  NOR2X1 U54607 ( .A(n12212), .B(n46659), .Y(net212073) );
  NOR2X1 U54608 ( .A(n10982), .B(n46618), .Y(n46622) );
  NOR2X1 U54609 ( .A(n12188), .B(n46985), .Y(n46989) );
  NOR2X1 U54610 ( .A(n12643), .B(n46086), .Y(net212831) );
  NOR2X1 U54611 ( .A(n12602), .B(n45795), .Y(net213200) );
  NOR2X1 U54612 ( .A(n12611), .B(n45532), .Y(n45536) );
  NOR2X1 U54613 ( .A(n11613), .B(n43462), .Y(net216400) );
  NOR2X1 U54614 ( .A(n11614), .B(n43447), .Y(net216427) );
  NOR2X1 U54615 ( .A(n11607), .B(n43487), .Y(net216355) );
  NOR2X1 U54616 ( .A(n11586), .B(n44622), .Y(net214678) );
  NOR2X1 U54617 ( .A(net271956), .B(n46625), .Y(net212164) );
  NOR2X1 U54618 ( .A(n11585), .B(n43529), .Y(n43533) );
  NOR2X1 U54619 ( .A(n40389), .B(n46077), .Y(net212856) );
  NOR2X1 U54620 ( .A(n12639), .B(n45582), .Y(net213542) );
  NOR2X1 U54621 ( .A(n43492), .B(net260900), .Y(net216346) );
  NOR2X1 U54622 ( .A(n47865), .B(net209111), .Y(net210353) );
  NOR2X1 U54623 ( .A(n47866), .B(net209087), .Y(net210348) );
  NOR2X1 U54624 ( .A(n46616), .B(net209136), .Y(net212189) );
  NOR2X1 U54625 ( .A(n45542), .B(net209697), .Y(n45546) );
  XOR2X1 U54626 ( .A(n32569), .B(n36776), .Y(n45542) );
  NOR2X1 U54627 ( .A(n45562), .B(net260925), .Y(net213603) );
  XOR2X1 U54628 ( .A(n32601), .B(n36784), .Y(n45562) );
  NOR2X1 U54629 ( .A(n45797), .B(net209689), .Y(net213190) );
  NOR2X1 U54630 ( .A(n12167), .B(n45589), .Y(net213507) );
  NOR2X1 U54631 ( .A(n46653), .B(net212088), .Y(n46657) );
  NOR2X1 U54632 ( .A(n46980), .B(net211602), .Y(net211597) );
  NOR2X1 U54633 ( .A(n46990), .B(net261069), .Y(net211563) );
  NOR2X1 U54634 ( .A(n46667), .B(net212037), .Y(n46671) );
  NOR2X1 U54635 ( .A(n46973), .B(net211640), .Y(net211635) );
  NOR2X1 U54636 ( .A(n46983), .B(net272417), .Y(net211579) );
  NOR2X1 U54637 ( .A(n11933), .B(n45588), .Y(net213512) );
  NOR2X1 U54638 ( .A(n45790), .B(net213230), .Y(net213225) );
  NOR2X1 U54639 ( .A(n44382), .B(net214783), .Y(net215060) );
  XOR2X1 U54640 ( .A(n32628), .B(n36828), .Y(n44382) );
  NOR2X1 U54641 ( .A(n44623), .B(net261422), .Y(net214672) );
  NOR2X1 U54642 ( .A(n44357), .B(net214756), .Y(n44361) );
  XOR2X1 U54643 ( .A(n32524), .B(n36828), .Y(n44357) );
  CLKBUFX3 U54644 ( .A(n32983), .Y(n41984) );
  CLKBUFX3 U54645 ( .A(n32975), .Y(n41985) );
  CLKBUFX3 U54646 ( .A(n32967), .Y(n41986) );
  CLKBUFX3 U54647 ( .A(n32959), .Y(n41987) );
  CLKBUFX3 U54648 ( .A(n32951), .Y(n41988) );
  CLKBUFX3 U54649 ( .A(n32943), .Y(n41989) );
  CLKBUFX3 U54650 ( .A(n32935), .Y(n41990) );
  CLKBUFX3 U54651 ( .A(n32927), .Y(n41991) );
  CLKBUFX3 U54652 ( .A(n32919), .Y(n41992) );
  CLKBUFX3 U54653 ( .A(n32911), .Y(n41993) );
  CLKBUFX3 U54654 ( .A(n32903), .Y(n41994) );
  CLKBUFX3 U54655 ( .A(n32895), .Y(n41995) );
  CLKBUFX3 U54656 ( .A(n32887), .Y(n41996) );
  CLKBUFX3 U54657 ( .A(n32879), .Y(n41997) );
  CLKBUFX3 U54658 ( .A(n32979), .Y(n42243) );
  CLKBUFX3 U54659 ( .A(n32971), .Y(n42244) );
  CLKBUFX3 U54660 ( .A(n32963), .Y(n42245) );
  CLKBUFX3 U54661 ( .A(n32955), .Y(n42246) );
  CLKBUFX3 U54662 ( .A(n32947), .Y(n42247) );
  CLKBUFX3 U54663 ( .A(n32939), .Y(n42248) );
  CLKBUFX3 U54664 ( .A(n32931), .Y(n42249) );
  CLKBUFX3 U54665 ( .A(n32923), .Y(n42250) );
  CLKBUFX3 U54666 ( .A(n32915), .Y(n42251) );
  CLKBUFX3 U54667 ( .A(n32907), .Y(n42252) );
  CLKBUFX3 U54668 ( .A(n32899), .Y(n42253) );
  CLKBUFX3 U54669 ( .A(n32891), .Y(n42254) );
  CLKBUFX3 U54670 ( .A(n32883), .Y(n42255) );
  CLKBUFX3 U54671 ( .A(n32875), .Y(n42256) );
  OR3X2 U54672 ( .A(n9892), .B(n9893), .C(n9894), .Y(n34511) );
  OAI221XL U54673 ( .A0(n42701), .A1(n40182), .B0(n9671), .B1(net266255), .C0(
        n9895), .Y(n9894) );
  AOI211X1 U54674 ( .A0(n50092), .A1(n9966), .B0(n9872), .C0(n9870), .Y(n9892)
         );
  OAI32X1 U54675 ( .A0(n9921), .A1(n9922), .A2(n42735), .B0(n40313), .B1(n9923), .Y(n9893) );
  OAI222XL U54676 ( .A0(n49540), .A1(n42728), .B0(n49548), .B1(n41797), .C0(
        n34475), .C1(n43044), .Y(n19483) );
  OAI222XL U54677 ( .A0(n49548), .A1(n42728), .B0(n49540), .B1(n42729), .C0(
        n34483), .C1(n43044), .Y(n19445) );
  OAI222XL U54678 ( .A0(n49548), .A1(n42729), .B0(n34475), .B1(n43039), .C0(
        n34491), .C1(n43043), .Y(n19407) );
  OAI222XL U54679 ( .A0(n49541), .A1(n42728), .B0(n49549), .B1(n41797), .C0(
        n34476), .C1(n43044), .Y(n19479) );
  OAI222XL U54680 ( .A0(n49549), .A1(n42728), .B0(n49541), .B1(n42729), .C0(
        n34484), .C1(n43044), .Y(n19441) );
  OAI222XL U54681 ( .A0(n49549), .A1(n42730), .B0(n34476), .B1(n43039), .C0(
        n34492), .C1(n43043), .Y(n19403) );
  OAI222XL U54682 ( .A0(n49542), .A1(n42728), .B0(n49550), .B1(n41797), .C0(
        n34477), .C1(n43044), .Y(n19475) );
  OAI222XL U54683 ( .A0(n49550), .A1(n42728), .B0(n49542), .B1(n42729), .C0(
        n34485), .C1(n43044), .Y(n19437) );
  OAI222XL U54684 ( .A0(n49550), .A1(n42730), .B0(n34477), .B1(n43039), .C0(
        n34493), .C1(n43044), .Y(n19399) );
  OAI222XL U54685 ( .A0(n49543), .A1(n42728), .B0(n49551), .B1(n41797), .C0(
        n34478), .C1(n43044), .Y(n19471) );
  OAI222XL U54686 ( .A0(n49551), .A1(n42728), .B0(n49543), .B1(n42729), .C0(
        n34486), .C1(n43043), .Y(n19433) );
  OAI222XL U54687 ( .A0(n49551), .A1(n42730), .B0(n34478), .B1(n43039), .C0(
        n34494), .C1(n43043), .Y(n19395) );
  OAI222XL U54688 ( .A0(n49544), .A1(n42728), .B0(n49552), .B1(n41797), .C0(
        n34479), .C1(n43044), .Y(n19467) );
  OAI222XL U54689 ( .A0(n49552), .A1(n19420), .B0(n49544), .B1(n42729), .C0(
        n34487), .C1(n43043), .Y(n19429) );
  OAI222XL U54690 ( .A0(n49552), .A1(n42729), .B0(n34479), .B1(n43040), .C0(
        n34495), .C1(n43043), .Y(n19391) );
  OAI222XL U54691 ( .A0(n49545), .A1(n19420), .B0(n49553), .B1(n41797), .C0(
        n34480), .C1(n43044), .Y(n19463) );
  OAI222XL U54692 ( .A0(n49553), .A1(n42728), .B0(n49545), .B1(n42730), .C0(
        n34488), .C1(n43043), .Y(n19425) );
  OAI222XL U54693 ( .A0(n49553), .A1(n42730), .B0(n34480), .B1(n43039), .C0(
        n34496), .C1(n43043), .Y(n19387) );
  OAI222XL U54694 ( .A0(n49546), .A1(n42728), .B0(n49554), .B1(n41797), .C0(
        n34481), .C1(n43044), .Y(n19459) );
  OAI222XL U54695 ( .A0(n49554), .A1(n42728), .B0(n49546), .B1(n42730), .C0(
        n34489), .C1(n43043), .Y(n19421) );
  OAI222XL U54696 ( .A0(n49554), .A1(n42730), .B0(n34481), .B1(n43039), .C0(
        n34497), .C1(n43043), .Y(n19383) );
  OAI222XL U54697 ( .A0(n49547), .A1(n42728), .B0(n49555), .B1(n41797), .C0(
        n34482), .C1(n43044), .Y(n19452) );
  OAI222XL U54698 ( .A0(n49555), .A1(n42730), .B0(n34482), .B1(n43040), .C0(
        n34498), .C1(n43043), .Y(n19377) );
  OAI222XL U54699 ( .A0(n49555), .A1(n19420), .B0(n49547), .B1(n42729), .C0(
        n34490), .C1(n43043), .Y(n19413) );
  NOR4X1 U54700 ( .A(n23664), .B(n23663), .C(n23662), .D(n23661), .Y(net212565) );
  NOR2X1 U54701 ( .A(n20834), .B(n20832), .Y(net211576) );
  NOR4X1 U54702 ( .A(n25696), .B(n25695), .C(n25694), .D(n25693), .Y(net214955) );
  NOR2X1 U54703 ( .A(n20434), .B(n20433), .Y(net211560) );
  NOR4X1 U54704 ( .A(n20432), .B(n20431), .C(n20430), .D(n20429), .Y(net211561) );
  NOR2X1 U54705 ( .A(n25878), .B(n25877), .Y(net214990) );
  NOR4X1 U54706 ( .A(n25876), .B(n25875), .C(n25874), .D(n25873), .Y(net214991) );
  NOR2X1 U54707 ( .A(n25788), .B(n25787), .Y(net214981) );
  NOR4X1 U54708 ( .A(n25786), .B(n25785), .C(n25784), .D(n25783), .Y(net214982) );
  NOR2X1 U54709 ( .A(n25728), .B(n25727), .Y(net214963) );
  NOR4X1 U54710 ( .A(n25726), .B(n25725), .C(n25724), .D(n25723), .Y(net214964) );
  NOR2X1 U54711 ( .A(n20486), .B(n20485), .Y(net211189) );
  NOR4X1 U54712 ( .A(n20484), .B(n20483), .C(n20482), .D(n20481), .Y(net211190) );
  NOR4X1 U54713 ( .A(n20937), .B(n20936), .C(n20935), .D(n20934), .Y(net211611) );
  NOR2X1 U54714 ( .A(n23290), .B(n23289), .Y(net213212) );
  NOR4X1 U54715 ( .A(n23288), .B(n23287), .C(n23286), .D(n23285), .Y(net213213) );
  XNOR2X1 U54716 ( .A(n36844), .B(n32610), .Y(net213598) );
  NOR2X1 U54717 ( .A(n24548), .B(n24546), .Y(net213599) );
  NOR4X1 U54718 ( .A(n25756), .B(n25755), .C(n25754), .D(n25753), .Y(net214973) );
  NOR2X1 U54719 ( .A(n20949), .B(n20948), .Y(net211615) );
  NOR4X1 U54720 ( .A(n20947), .B(n20946), .C(n20945), .D(n20944), .Y(net211616) );
  NOR4X1 U54721 ( .A(n20821), .B(n20820), .C(n20819), .D(n20818), .Y(net211594) );
  NOR2X1 U54722 ( .A(n20959), .B(n20958), .Y(net211620) );
  NOR4X1 U54723 ( .A(n20957), .B(n20956), .C(n20955), .D(n20954), .Y(net211621) );
  NOR4X1 U54724 ( .A(n20810), .B(n20809), .C(n20808), .D(n20807), .Y(net211588) );
  NOR4X1 U54725 ( .A(n23654), .B(n23653), .C(n23652), .D(n23651), .Y(net213315) );
  NOR2X1 U54726 ( .A(n20085), .B(n20084), .Y(net211440) );
  NOR4X1 U54727 ( .A(n20083), .B(n20082), .C(n20081), .D(n20080), .Y(net211441) );
  NOR2X1 U54728 ( .A(n20075), .B(n20074), .Y(net211435) );
  NOR2X1 U54729 ( .A(n20095), .B(n20094), .Y(net211445) );
  NOR4X1 U54730 ( .A(n20093), .B(n20092), .C(n20091), .D(n20090), .Y(net211446) );
  NOR4X1 U54731 ( .A(n24515), .B(n24514), .C(n24513), .D(n24512), .Y(net213595) );
  NOR2X1 U54732 ( .A(n23686), .B(n23685), .Y(net212554) );
  NOR4X1 U54733 ( .A(n23684), .B(n23683), .C(n23682), .D(n23681), .Y(net212555) );
  NOR2X1 U54734 ( .A(n23676), .B(n23675), .Y(net212559) );
  NOR4X1 U54735 ( .A(n23674), .B(n23673), .C(n23672), .D(n23671), .Y(net212560) );
  NAND4X1 U54736 ( .A(n44344), .B(n44343), .C(n44342), .D(n44341), .Y(n12597)
         );
  NOR2X1 U54737 ( .A(n26599), .B(n26598), .Y(n44342) );
  NOR4X1 U54738 ( .A(n26597), .B(n26596), .C(n26595), .D(n26594), .Y(n44341)
         );
  NAND4X1 U54739 ( .A(n44339), .B(n44338), .C(n44337), .D(n44336), .Y(n12808)
         );
  NOR2X1 U54740 ( .A(n26629), .B(n26628), .Y(n44337) );
  NOR4X1 U54741 ( .A(n26627), .B(n26626), .C(n26625), .D(n26624), .Y(n44336)
         );
  NOR2X1 U54742 ( .A(n20506), .B(n20505), .Y(net211184) );
  NOR4X1 U54743 ( .A(n20494), .B(n20493), .C(n20492), .D(n20491), .Y(net211170) );
  NOR2X1 U54744 ( .A(n26419), .B(n26418), .Y(net212569) );
  NOR4X1 U54745 ( .A(n26417), .B(n26416), .C(n26415), .D(n26414), .Y(net212570) );
  NAND4X1 U54746 ( .A(n45541), .B(n45540), .C(n45539), .D(n45538), .Y(
        net209103) );
  NOR2X1 U54747 ( .A(n24651), .B(n24649), .Y(n45539) );
  NOR4X1 U54748 ( .A(n24648), .B(n24647), .C(n24646), .D(n24645), .Y(n45538)
         );
  NOR4X1 U54749 ( .A(n24535), .B(n24534), .C(n24533), .D(n24532), .Y(net213585) );
  NOR4X1 U54750 ( .A(n24505), .B(n24504), .C(n24503), .D(n24502), .Y(net213590) );
  NOR2X1 U54751 ( .A(n20055), .B(n20054), .Y(net211470) );
  NOR4X1 U54752 ( .A(n20053), .B(n20052), .C(n20051), .D(n20050), .Y(net211471) );
  NOR4X1 U54753 ( .A(n20033), .B(n20032), .C(n20031), .D(n20030), .Y(net211461) );
  NOR4X1 U54754 ( .A(n21787), .B(n21786), .C(n21785), .D(n21784), .Y(net212030) );
  NOR4X1 U54755 ( .A(n26537), .B(n26536), .C(n26535), .D(n26534), .Y(net215189) );
  OAI22XL U54756 ( .A0(n34489), .A1(n42452), .B0(n34497), .B1(n43039), .Y(
        n19293) );
  OAI22XL U54757 ( .A0(n34488), .A1(n42452), .B0(n34496), .B1(n43039), .Y(
        n19299) );
  OAI22XL U54758 ( .A0(n34487), .A1(n42452), .B0(n34495), .B1(n43039), .Y(
        n19305) );
  OAI22XL U54759 ( .A0(n34486), .A1(n42453), .B0(n34494), .B1(n43039), .Y(
        n19311) );
  OAI22XL U54760 ( .A0(n34485), .A1(n42452), .B0(n34493), .B1(n43039), .Y(
        n19317) );
  OAI22XL U54761 ( .A0(n34484), .A1(n42453), .B0(n34492), .B1(n43039), .Y(
        n19323) );
  OAI22XL U54762 ( .A0(n34483), .A1(n42453), .B0(n34491), .B1(n43039), .Y(
        n19329) );
  OAI22XL U54763 ( .A0(n34490), .A1(n42452), .B0(n34498), .B1(n43039), .Y(
        n19284) );
  OAI22XL U54764 ( .A0(n34491), .A1(n42450), .B0(n34499), .B1(n36935), .Y(
        n19371) );
  OAI22XL U54765 ( .A0(n34492), .A1(n42450), .B0(n34500), .B1(n36935), .Y(
        n19367) );
  OAI22XL U54766 ( .A0(n34493), .A1(n42450), .B0(n34501), .B1(n36935), .Y(
        n19363) );
  OAI22XL U54767 ( .A0(n34494), .A1(n42450), .B0(n34502), .B1(n36935), .Y(
        n19359) );
  OAI22XL U54768 ( .A0(n34495), .A1(n42450), .B0(n34503), .B1(n36935), .Y(
        n19355) );
  OAI22XL U54769 ( .A0(n34496), .A1(n42450), .B0(n34504), .B1(n36935), .Y(
        n19351) );
  OAI22XL U54770 ( .A0(n34497), .A1(n42450), .B0(n34505), .B1(n36935), .Y(
        n19347) );
  OAI22XL U54771 ( .A0(n34498), .A1(n42450), .B0(n34506), .B1(n36935), .Y(
        n19339) );
  OAI22XL U54772 ( .A0(n34478), .A1(n43041), .B0(n41300), .B1(n42450), .Y(
        n19507) );
  OAI22XL U54773 ( .A0(n34479), .A1(n43041), .B0(n41331), .B1(n42450), .Y(
        n19503) );
  OAI22XL U54774 ( .A0(n34477), .A1(n43041), .B0(n36807), .B1(n42450), .Y(
        n19511) );
  OAI22XL U54775 ( .A0(n34476), .A1(n43041), .B0(n36841), .B1(n42450), .Y(
        n19515) );
  NOR4X1 U54776 ( .A(n20863), .B(n20862), .C(n20861), .D(n20860), .Y(net210366) );
  NAND4X1 U54777 ( .A(n44404), .B(n44403), .C(n44402), .D(n44401), .Y(
        net213653) );
  NOR2X1 U54778 ( .A(n25818), .B(n25817), .Y(n44402) );
  NOR4X1 U54779 ( .A(n25816), .B(n25815), .C(n25814), .D(n25813), .Y(n44401)
         );
  NAND4X1 U54780 ( .A(n44398), .B(n44397), .C(n44396), .D(n44395), .Y(
        net213602) );
  NOR2X1 U54781 ( .A(n25938), .B(n25937), .Y(n44396) );
  NOR4X1 U54782 ( .A(n25936), .B(n25935), .C(n25934), .D(n25933), .Y(n44395)
         );
  NAND4X1 U54783 ( .A(n45571), .B(n45570), .C(n45569), .D(n45568), .Y(
        net211590) );
  XNOR2X1 U54784 ( .A(n36839), .B(n32554), .Y(n45570) );
  NOR2X1 U54785 ( .A(n24527), .B(n24526), .Y(n45569) );
  NOR4X1 U54786 ( .A(n24525), .B(n24524), .C(n24523), .D(n24522), .Y(n45568)
         );
  NAND4X1 U54787 ( .A(n44319), .B(n44318), .C(n44317), .D(n44316), .Y(n12395)
         );
  NOR2X1 U54788 ( .A(n26569), .B(n26568), .Y(n44317) );
  NOR4X1 U54789 ( .A(n26567), .B(n26566), .C(n26565), .D(n26564), .Y(n44316)
         );
  NOR4X1 U54790 ( .A(n20043), .B(n20042), .C(n20041), .D(n20040), .Y(net211466) );
  NOR4X1 U54791 ( .A(n20873), .B(n20872), .C(n20871), .D(n20870), .Y(net210371) );
  OAI22XL U54792 ( .A0(net171523), .A1(net264532), .B0(n9653), .B1(n9754), .Y(
        n34516) );
  NOR2X1 U54793 ( .A(n10772), .B(n47050), .Y(net211443) );
  NOR2X1 U54794 ( .A(n10771), .B(n47052), .Y(net211433) );
  NOR2X1 U54795 ( .A(n10763), .B(n46991), .Y(net211558) );
  NOR2X1 U54796 ( .A(n10292), .B(n44422), .Y(net214952) );
  NOR2X1 U54797 ( .A(n11538), .B(n44315), .Y(n44319) );
  NOR2X1 U54798 ( .A(n11544), .B(n46306), .Y(net212567) );
  NOR2X1 U54799 ( .A(n11896), .B(n45564), .Y(net213592) );
  NOR2X1 U54800 ( .A(n10928), .B(n47047), .Y(net211458) );
  NOR2X1 U54801 ( .A(n11543), .B(n44340), .Y(n44344) );
  XOR2X1 U54802 ( .A(n32428), .B(n36823), .Y(n44340) );
  NOR2X1 U54803 ( .A(n11902), .B(n45567), .Y(n45571) );
  NOR2X1 U54804 ( .A(n11893), .B(n45565), .Y(net213587) );
  NOR2X1 U54805 ( .A(n11895), .B(n45566), .Y(net213582) );
  NOR2X1 U54806 ( .A(n11541), .B(n44320), .Y(net215186) );
  XOR2X1 U54807 ( .A(n32412), .B(n36824), .Y(n44320) );
  NOR2X1 U54808 ( .A(n10927), .B(n47046), .Y(net211463) );
  NOR2X1 U54809 ( .A(n11566), .B(n44400), .Y(n44404) );
  XOR2X1 U54810 ( .A(n32588), .B(n36825), .Y(n44400) );
  NOR2X1 U54811 ( .A(n10941), .B(n46977), .Y(net211613) );
  NOR2X1 U54812 ( .A(net259677), .B(n44410), .Y(net214988) );
  XOR2X1 U54813 ( .A(n32564), .B(n36830), .Y(n44410) );
  NOR2X1 U54814 ( .A(n11542), .B(n44335), .Y(n44339) );
  XOR2X1 U54815 ( .A(n32420), .B(n36828), .Y(n44335) );
  NOR2X1 U54816 ( .A(n11894), .B(n45793), .Y(net213210) );
  NOR2X1 U54817 ( .A(n10939), .B(n46978), .Y(net211608) );
  NOR2X1 U54818 ( .A(n12196), .B(n46981), .Y(net211591) );
  NOR2X1 U54819 ( .A(n12190), .B(n47051), .Y(net211438) );
  NOR2X1 U54820 ( .A(n12408), .B(n44411), .Y(net214979) );
  XOR2X1 U54821 ( .A(n32540), .B(n36831), .Y(n44411) );
  NOR2X1 U54822 ( .A(net260394), .B(n46309), .Y(net212552) );
  NOR2X1 U54823 ( .A(net260449), .B(n46307), .Y(net212562) );
  NOR2X1 U54824 ( .A(n12194), .B(n47045), .Y(net211468) );
  NOR2X1 U54825 ( .A(net260302), .B(n47280), .Y(net211167) );
  NOR2X1 U54826 ( .A(n12596), .B(n46308), .Y(net212557) );
  NOR2X1 U54827 ( .A(n12207), .B(n46976), .Y(net211618) );
  NOR2X1 U54828 ( .A(n47268), .B(net210555), .Y(net211187) );
  NOR2X1 U54829 ( .A(n47269), .B(net210556), .Y(net211182) );
  NOR2X1 U54830 ( .A(n12594), .B(n45716), .Y(net213312) );
  NOR2X1 U54831 ( .A(n47859), .B(net209101), .Y(net210363) );
  NOR2X1 U54832 ( .A(n47858), .B(net260830), .Y(net210368) );
  NOR2X1 U54833 ( .A(n46672), .B(net209124), .Y(net212027) );
  NOR2X1 U54834 ( .A(n46984), .B(net209099), .Y(net211574) );
  AO22X1 U54835 ( .A0(N23561), .A1(out_valid), .B0(n37191), .B1(n41791), .Y(
        n32384) );
  AO22X1 U54836 ( .A0(N23562), .A1(out_valid), .B0(n37194), .B1(n41791), .Y(
        n32395) );
  NOR2X1 U54837 ( .A(n46982), .B(net211590), .Y(net211585) );
  NOR2X1 U54838 ( .A(n45537), .B(net213653), .Y(n45541) );
  XOR2X1 U54839 ( .A(n32577), .B(n36779), .Y(n45537) );
  NOR2X1 U54840 ( .A(n45563), .B(net272583), .Y(net213597) );
  NOR2X1 U54841 ( .A(n44394), .B(net214782), .Y(n44398) );
  XOR2X1 U54842 ( .A(n32620), .B(n36821), .Y(n44394) );
  NOR2X1 U54843 ( .A(n44421), .B(net272625), .Y(net214961) );
  NOR2X1 U54844 ( .A(n44416), .B(net272620), .Y(net214970) );
  NAND2X1 U54845 ( .A(n19251), .B(n19252), .Y(n36582) );
  AOI221XL U54846 ( .A0(n37530), .A1(data[17]), .B0(n37182), .B1(data[9]),
        .C0(n19253), .Y(n19252) );
  AOI222XL U54847 ( .A0(n19247), .A1(n50164), .B0(n19249), .B1(n50163), .C0(
        n42733), .C1(data[1]), .Y(n19251) );
  OAI22XL U54848 ( .A0(n49530), .A1(n50131), .B0(n34497), .B1(n42454), .Y(
        n19253) );
  NAND2X1 U54849 ( .A(n19255), .B(n19256), .Y(n36583) );
  AOI221XL U54850 ( .A0(n37530), .A1(data[18]), .B0(n37182), .B1(data[10]),
        .C0(n19257), .Y(n19256) );
  AOI222XL U54851 ( .A0(n19247), .A1(n50162), .B0(n19249), .B1(n50161), .C0(
        n42734), .C1(data[2]), .Y(n19255) );
  OAI22XL U54852 ( .A0(n49529), .A1(n50131), .B0(n34496), .B1(n42454), .Y(
        n19257) );
  NAND2X1 U54853 ( .A(n19259), .B(n19260), .Y(n36584) );
  AOI221XL U54854 ( .A0(n37530), .A1(data[19]), .B0(n37182), .B1(data[11]),
        .C0(n19261), .Y(n19260) );
  AOI222XL U54855 ( .A0(n19247), .A1(n50160), .B0(n19249), .B1(n50159), .C0(
        n42734), .C1(data[3]), .Y(n19259) );
  OAI22XL U54856 ( .A0(n49528), .A1(n50131), .B0(n34495), .B1(n42454), .Y(
        n19261) );
  NAND2X1 U54857 ( .A(n19263), .B(n19264), .Y(n36585) );
  AOI221XL U54858 ( .A0(n37530), .A1(data[20]), .B0(n37182), .B1(data[12]),
        .C0(n19265), .Y(n19264) );
  AOI222XL U54859 ( .A0(n19247), .A1(n50158), .B0(n19249), .B1(n50157), .C0(
        n42733), .C1(data[4]), .Y(n19263) );
  OAI22XL U54860 ( .A0(n49527), .A1(n50131), .B0(n34494), .B1(n50114), .Y(
        n19265) );
  NAND2X1 U54861 ( .A(n19267), .B(n19268), .Y(n36586) );
  AOI221XL U54862 ( .A0(n37530), .A1(data[21]), .B0(n37182), .B1(data[13]),
        .C0(n19269), .Y(n19268) );
  AOI222XL U54863 ( .A0(n19247), .A1(n50156), .B0(n19249), .B1(n50155), .C0(
        n42734), .C1(data[5]), .Y(n19267) );
  OAI22XL U54864 ( .A0(n49526), .A1(n50131), .B0(n34493), .B1(n50114), .Y(
        n19269) );
  NAND2X1 U54865 ( .A(n19271), .B(n19272), .Y(n36587) );
  AOI221XL U54866 ( .A0(n37530), .A1(data[22]), .B0(n37182), .B1(data[14]),
        .C0(n19273), .Y(n19272) );
  AOI222XL U54867 ( .A0(n19247), .A1(n50154), .B0(n19249), .B1(n50153), .C0(
        n42733), .C1(data[6]), .Y(n19271) );
  OAI22XL U54868 ( .A0(n49525), .A1(n50131), .B0(n34492), .B1(n50114), .Y(
        n19273) );
  NAND2X1 U54869 ( .A(n19275), .B(n19276), .Y(n36588) );
  AOI221XL U54870 ( .A0(n37530), .A1(data[23]), .B0(n37182), .B1(data[15]),
        .C0(n19277), .Y(n19276) );
  AOI222XL U54871 ( .A0(n19247), .A1(n50152), .B0(n19249), .B1(n50151), .C0(
        n42734), .C1(data[7]), .Y(n19275) );
  OAI22XL U54872 ( .A0(n49524), .A1(n50131), .B0(n34491), .B1(n50114), .Y(
        n19277) );
  NAND2X1 U54873 ( .A(n19240), .B(n19241), .Y(n36581) );
  AOI221XL U54874 ( .A0(data[16]), .A1(n37530), .B0(n37182), .B1(data[8]),
        .C0(n19243), .Y(n19241) );
  AOI222XL U54875 ( .A0(n19247), .A1(n50150), .B0(n19249), .B1(n49557), .C0(
        n42733), .C1(data[0]), .Y(n19240) );
  OAI22XL U54876 ( .A0(n49531), .A1(n50131), .B0(n34498), .B1(n42454), .Y(
        n19243) );
  OAI21XL U54877 ( .A0(n9652), .A1(net266151), .B0(n50113), .Y(n34507) );
  CLKINVX1 U54878 ( .A(n9754), .Y(n50113) );
  CLKBUFX3 U54879 ( .A(n32871), .Y(n41998) );
  CLKBUFX3 U54880 ( .A(n32863), .Y(n41999) );
  CLKBUFX3 U54881 ( .A(n32855), .Y(n42000) );
  CLKBUFX3 U54882 ( .A(n32847), .Y(n42001) );
  CLKBUFX3 U54883 ( .A(n32839), .Y(n42002) );
  CLKBUFX3 U54884 ( .A(n32831), .Y(n42003) );
  CLKBUFX3 U54885 ( .A(n32823), .Y(n42004) );
  CLKBUFX3 U54886 ( .A(n32815), .Y(n42005) );
  CLKBUFX3 U54887 ( .A(n32807), .Y(n42006) );
  CLKBUFX3 U54888 ( .A(n32799), .Y(n42007) );
  CLKBUFX3 U54889 ( .A(n32791), .Y(n42008) );
  CLKBUFX3 U54890 ( .A(n32783), .Y(n42009) );
  CLKBUFX3 U54891 ( .A(n32775), .Y(n42010) );
  CLKBUFX3 U54892 ( .A(n32767), .Y(n42011) );
  CLKBUFX3 U54893 ( .A(n32759), .Y(n42012) );
  CLKBUFX3 U54894 ( .A(n32751), .Y(n42013) );
  CLKBUFX3 U54895 ( .A(n32743), .Y(n42014) );
  CLKBUFX3 U54896 ( .A(n32735), .Y(n42015) );
  CLKBUFX3 U54897 ( .A(n32727), .Y(n42016) );
  CLKBUFX3 U54898 ( .A(n32719), .Y(n42017) );
  CLKBUFX3 U54899 ( .A(n32711), .Y(n42018) );
  CLKBUFX3 U54900 ( .A(n32703), .Y(n42019) );
  CLKBUFX3 U54901 ( .A(n32695), .Y(n42020) );
  CLKBUFX3 U54902 ( .A(n32687), .Y(n42021) );
  CLKBUFX3 U54903 ( .A(n32679), .Y(n42022) );
  CLKBUFX3 U54904 ( .A(n32671), .Y(n42023) );
  CLKBUFX3 U54905 ( .A(n32663), .Y(n42024) );
  CLKBUFX3 U54906 ( .A(n32655), .Y(n42025) );
  CLKBUFX3 U54907 ( .A(n32647), .Y(n42026) );
  CLKBUFX3 U54908 ( .A(n32639), .Y(n42027) );
  CLKBUFX3 U54909 ( .A(n32631), .Y(n42028) );
  CLKBUFX3 U54910 ( .A(n32623), .Y(n42029) );
  CLKBUFX3 U54911 ( .A(n32615), .Y(n42030) );
  CLKBUFX3 U54912 ( .A(n32607), .Y(n42031) );
  CLKBUFX3 U54913 ( .A(n32599), .Y(n42032) );
  CLKBUFX3 U54914 ( .A(n32591), .Y(n42033) );
  CLKBUFX3 U54915 ( .A(n32583), .Y(n42034) );
  CLKBUFX3 U54916 ( .A(n32575), .Y(n42035) );
  CLKBUFX3 U54917 ( .A(n32567), .Y(n42036) );
  CLKBUFX3 U54918 ( .A(n32559), .Y(n42037) );
  CLKBUFX3 U54919 ( .A(n32551), .Y(n42038) );
  CLKBUFX3 U54920 ( .A(n32543), .Y(n42039) );
  CLKBUFX3 U54921 ( .A(n32535), .Y(n42040) );
  CLKBUFX3 U54922 ( .A(n32527), .Y(n42041) );
  CLKBUFX3 U54923 ( .A(n32519), .Y(n42042) );
  CLKBUFX3 U54924 ( .A(n32511), .Y(n42043) );
  CLKBUFX3 U54925 ( .A(n32503), .Y(n42044) );
  CLKBUFX3 U54926 ( .A(n32495), .Y(n42045) );
  CLKBUFX3 U54927 ( .A(n32487), .Y(n42046) );
  CLKBUFX3 U54928 ( .A(n32479), .Y(n42047) );
  CLKBUFX3 U54929 ( .A(n32471), .Y(n42048) );
  CLKBUFX3 U54930 ( .A(n32463), .Y(n42049) );
  CLKBUFX3 U54931 ( .A(n32455), .Y(n42050) );
  CLKBUFX3 U54932 ( .A(n32439), .Y(n42052) );
  CLKBUFX3 U54933 ( .A(n32447), .Y(n42051) );
  CLKBUFX3 U54934 ( .A(n32431), .Y(n42053) );
  CLKBUFX3 U54935 ( .A(n32423), .Y(n42054) );
  CLKBUFX3 U54936 ( .A(n32415), .Y(n42055) );
  CLKBUFX3 U54937 ( .A(n32867), .Y(n42257) );
  CLKBUFX3 U54938 ( .A(n32859), .Y(n42258) );
  CLKBUFX3 U54939 ( .A(n32851), .Y(n42259) );
  CLKBUFX3 U54940 ( .A(n32843), .Y(n42260) );
  CLKBUFX3 U54941 ( .A(n32835), .Y(n42261) );
  CLKBUFX3 U54942 ( .A(n32827), .Y(n42262) );
  CLKBUFX3 U54943 ( .A(n32819), .Y(n42263) );
  CLKBUFX3 U54944 ( .A(n32811), .Y(n42264) );
  CLKBUFX3 U54945 ( .A(n32803), .Y(n42265) );
  CLKBUFX3 U54946 ( .A(n32795), .Y(n42266) );
  CLKBUFX3 U54947 ( .A(n32787), .Y(n42267) );
  CLKBUFX3 U54948 ( .A(n32779), .Y(n42268) );
  CLKBUFX3 U54949 ( .A(n32771), .Y(n42269) );
  CLKBUFX3 U54950 ( .A(n32763), .Y(n42270) );
  CLKBUFX3 U54951 ( .A(n32755), .Y(n42271) );
  CLKBUFX3 U54952 ( .A(n32747), .Y(n42272) );
  CLKBUFX3 U54953 ( .A(n32739), .Y(n42273) );
  CLKBUFX3 U54954 ( .A(n32731), .Y(n42274) );
  CLKBUFX3 U54955 ( .A(n32723), .Y(n42275) );
  CLKBUFX3 U54956 ( .A(n32715), .Y(n42276) );
  CLKBUFX3 U54957 ( .A(n32707), .Y(n42277) );
  CLKBUFX3 U54958 ( .A(n32699), .Y(n42278) );
  CLKBUFX3 U54959 ( .A(n32691), .Y(n42279) );
  CLKBUFX3 U54960 ( .A(n32683), .Y(n42280) );
  CLKBUFX3 U54961 ( .A(n32675), .Y(n42281) );
  CLKBUFX3 U54962 ( .A(n32667), .Y(n42282) );
  CLKBUFX3 U54963 ( .A(n32659), .Y(n42283) );
  CLKBUFX3 U54964 ( .A(n32651), .Y(n42284) );
  CLKBUFX3 U54965 ( .A(n32643), .Y(n42285) );
  CLKBUFX3 U54966 ( .A(n32635), .Y(n42286) );
  CLKBUFX3 U54967 ( .A(n32627), .Y(n42287) );
  CLKBUFX3 U54968 ( .A(n32619), .Y(n42288) );
  CLKBUFX3 U54969 ( .A(n32611), .Y(n42289) );
  CLKBUFX3 U54970 ( .A(n32603), .Y(n42290) );
  CLKBUFX3 U54971 ( .A(n32595), .Y(n42291) );
  CLKBUFX3 U54972 ( .A(n32587), .Y(n42292) );
  CLKBUFX3 U54973 ( .A(n32579), .Y(n42293) );
  CLKBUFX3 U54974 ( .A(n32571), .Y(n42294) );
  CLKBUFX3 U54975 ( .A(n32563), .Y(n42295) );
  CLKBUFX3 U54976 ( .A(n32555), .Y(n42296) );
  CLKBUFX3 U54977 ( .A(n32547), .Y(n42297) );
  CLKBUFX3 U54978 ( .A(n32539), .Y(n42298) );
  CLKBUFX3 U54979 ( .A(n32531), .Y(n42299) );
  CLKBUFX3 U54980 ( .A(n32523), .Y(n42300) );
  CLKBUFX3 U54981 ( .A(n32515), .Y(n42301) );
  CLKBUFX3 U54982 ( .A(n32507), .Y(n42302) );
  CLKBUFX3 U54983 ( .A(n32499), .Y(n42303) );
  CLKBUFX3 U54984 ( .A(n32491), .Y(n42304) );
  CLKBUFX3 U54985 ( .A(n32483), .Y(n42305) );
  CLKBUFX3 U54986 ( .A(n32475), .Y(n42306) );
  CLKBUFX3 U54987 ( .A(n32467), .Y(n42307) );
  CLKBUFX3 U54988 ( .A(n32459), .Y(n42308) );
  CLKBUFX3 U54989 ( .A(n32451), .Y(n42309) );
  CLKBUFX3 U54990 ( .A(n32435), .Y(n42311) );
  CLKBUFX3 U54991 ( .A(n32443), .Y(n42310) );
  CLKBUFX3 U54992 ( .A(n32427), .Y(n42312) );
  CLKBUFX3 U54993 ( .A(n32419), .Y(n42313) );
  CLKBUFX3 U54994 ( .A(n32411), .Y(n42314) );
  CLKBUFX3 U54995 ( .A(n32407), .Y(n42056) );
  CLKBUFX3 U54996 ( .A(n32403), .Y(n42315) );
  OR4X1 U54997 ( .A(n19370), .B(n19371), .C(n19372), .D(n19373), .Y(n36604) );
  OAI22XL U54998 ( .A0(n49540), .A1(n42731), .B0(n49548), .B1(n37183), .Y(
        n19373) );
  OAI222XL U54999 ( .A0(n49532), .A1(n37525), .B0(n36767), .B1(n19343), .C0(
        n49524), .C1(n19344), .Y(n19372) );
  OAI22XL U55000 ( .A0(n34483), .A1(n43038), .B0(n34475), .B1(n42454), .Y(
        n19370) );
  OR4X1 U55001 ( .A(n19366), .B(n19367), .C(n19368), .D(n19369), .Y(n36603) );
  OAI22XL U55002 ( .A0(n49541), .A1(n42731), .B0(n49549), .B1(n37183), .Y(
        n19369) );
  OAI222XL U55003 ( .A0(n49533), .A1(n37525), .B0(n36735), .B1(n19343), .C0(
        n49525), .C1(n19344), .Y(n19368) );
  OAI22XL U55004 ( .A0(n34484), .A1(n43038), .B0(n34476), .B1(n42454), .Y(
        n19366) );
  OR4X1 U55005 ( .A(n19362), .B(n19363), .C(n19364), .D(n19365), .Y(n36602) );
  OAI22XL U55006 ( .A0(n49542), .A1(n19292), .B0(n49550), .B1(n37183), .Y(
        n19365) );
  OAI222XL U55007 ( .A0(n49534), .A1(n42732), .B0(n42496), .B1(n19343), .C0(
        n49526), .C1(n19344), .Y(n19364) );
  OAI22XL U55008 ( .A0(n34485), .A1(n43038), .B0(n34477), .B1(n42454), .Y(
        n19362) );
  OR4X1 U55009 ( .A(n19358), .B(n19359), .C(n19360), .D(n19361), .Y(n36601) );
  OAI22XL U55010 ( .A0(n49543), .A1(n19292), .B0(n49551), .B1(n37183), .Y(
        n19361) );
  OAI222XL U55011 ( .A0(n49535), .A1(n42732), .B0(n36746), .B1(n19343), .C0(
        n49527), .C1(n19344), .Y(n19360) );
  OAI22XL U55012 ( .A0(n34486), .A1(n43038), .B0(n34478), .B1(n42453), .Y(
        n19358) );
  OR4X1 U55013 ( .A(n19354), .B(n19355), .C(n19356), .D(n19357), .Y(n36600) );
  OAI22XL U55014 ( .A0(n49544), .A1(n42731), .B0(n49552), .B1(n37183), .Y(
        n19357) );
  OAI222XL U55015 ( .A0(n49536), .A1(n42732), .B0(n36718), .B1(n19343), .C0(
        n49528), .C1(n19344), .Y(n19356) );
  OAI22XL U55016 ( .A0(n34487), .A1(n43038), .B0(n34479), .B1(n42452), .Y(
        n19354) );
  OR4X1 U55017 ( .A(n19350), .B(n19351), .C(n19352), .D(n19353), .Y(n36599) );
  OAI22XL U55018 ( .A0(n49545), .A1(n42731), .B0(n49553), .B1(n37183), .Y(
        n19353) );
  OAI222XL U55019 ( .A0(n49537), .A1(n42732), .B0(n36792), .B1(n19343), .C0(
        n49529), .C1(n19344), .Y(n19352) );
  OAI22XL U55020 ( .A0(n34488), .A1(n43038), .B0(n34480), .B1(n42453), .Y(
        n19350) );
  OR4X1 U55021 ( .A(n19346), .B(n19347), .C(n19348), .D(n19349), .Y(n36598) );
  OAI22XL U55022 ( .A0(n49546), .A1(n42731), .B0(n49554), .B1(n37183), .Y(
        n19349) );
  OAI222XL U55023 ( .A0(n49538), .A1(n42732), .B0(n36761), .B1(n19343), .C0(
        n49530), .C1(n19344), .Y(n19348) );
  OAI22XL U55024 ( .A0(n34489), .A1(n43038), .B0(n34481), .B1(n42452), .Y(
        n19346) );
  OR4X1 U55025 ( .A(n19338), .B(n19339), .C(n19340), .D(n19341), .Y(n36597) );
  OAI22XL U55026 ( .A0(n49547), .A1(n42731), .B0(n49555), .B1(n37183), .Y(
        n19341) );
  OAI222XL U55027 ( .A0(n49539), .A1(n42732), .B0(n42473), .B1(n19343), .C0(
        n49531), .C1(n19344), .Y(n19340) );
  OAI22XL U55028 ( .A0(n34490), .A1(n43038), .B0(n34482), .B1(n42453), .Y(
        n19338) );
  OR4X1 U55029 ( .A(n19445), .B(n19446), .C(n19447), .D(n19448), .Y(n36620) );
  OAI222XL U55030 ( .A0(n49524), .A1(n19417), .B0(n42584), .B1(n50128), .C0(
        n49532), .C1(n19419), .Y(n19447) );
  OAI22XL U55031 ( .A0(n36766), .A1(n43038), .B0(n36785), .B1(n42454), .Y(
        n19448) );
  OAI22XL U55032 ( .A0(n34491), .A1(n43042), .B0(n34475), .B1(n42450), .Y(
        n19446) );
  OR4X1 U55033 ( .A(n19441), .B(n19442), .C(n19443), .D(n19444), .Y(n36619) );
  OAI222XL U55034 ( .A0(n49525), .A1(n19417), .B0(n42569), .B1(n50128), .C0(
        n49533), .C1(n19419), .Y(n19443) );
  OAI22XL U55035 ( .A0(n36733), .A1(n43038), .B0(n36843), .B1(n42454), .Y(
        n19444) );
  OAI22XL U55036 ( .A0(n34492), .A1(n43042), .B0(n34476), .B1(n42450), .Y(
        n19442) );
  OR4X1 U55037 ( .A(n19437), .B(n19438), .C(n19439), .D(n19440), .Y(n36618) );
  OAI222XL U55038 ( .A0(n49526), .A1(n19417), .B0(n41323), .B1(n50128), .C0(
        n49534), .C1(n19419), .Y(n19439) );
  OAI22XL U55039 ( .A0(n42479), .A1(n43039), .B0(n36817), .B1(n42454), .Y(
        n19440) );
  OAI22XL U55040 ( .A0(n34493), .A1(n43042), .B0(n34477), .B1(n42451), .Y(
        n19438) );
  OR4X1 U55041 ( .A(n19433), .B(n19434), .C(n19435), .D(n19436), .Y(n36617) );
  OAI222XL U55042 ( .A0(n49527), .A1(n19417), .B0(n36825), .B1(n50128), .C0(
        n49535), .C1(n19419), .Y(n19435) );
  OAI22XL U55043 ( .A0(n36742), .A1(n43039), .B0(n41300), .B1(n42454), .Y(
        n19436) );
  OAI22XL U55044 ( .A0(n34494), .A1(n43042), .B0(n34478), .B1(n42451), .Y(
        n19434) );
  OR4X1 U55045 ( .A(n19429), .B(n19430), .C(n19431), .D(n19432), .Y(n36616) );
  OAI222XL U55046 ( .A0(n49528), .A1(n19417), .B0(n42554), .B1(n50128), .C0(
        n49536), .C1(n19419), .Y(n19431) );
  OAI22XL U55047 ( .A0(n36720), .A1(n43038), .B0(n41328), .B1(n42454), .Y(
        n19432) );
  OAI22XL U55048 ( .A0(n34495), .A1(n43042), .B0(n34479), .B1(n42451), .Y(
        n19430) );
  OR4X1 U55049 ( .A(n19425), .B(n19426), .C(n19427), .D(n19428), .Y(n36615) );
  OAI222XL U55050 ( .A0(n49529), .A1(n19417), .B0(n42544), .B1(n50128), .C0(
        n49537), .C1(n19419), .Y(n19427) );
  OAI22XL U55051 ( .A0(n36791), .A1(n43039), .B0(n41290), .B1(n42454), .Y(
        n19428) );
  OAI22XL U55052 ( .A0(n34496), .A1(n43042), .B0(n34480), .B1(n42451), .Y(
        n19426) );
  OR4X1 U55053 ( .A(n19421), .B(n19422), .C(n19423), .D(n19424), .Y(n36614) );
  OAI222XL U55054 ( .A0(n49530), .A1(n19417), .B0(n42517), .B1(n50128), .C0(
        n49538), .C1(n19419), .Y(n19423) );
  OAI22XL U55055 ( .A0(n36759), .A1(n43039), .B0(n41316), .B1(n42454), .Y(
        n19424) );
  OAI22XL U55056 ( .A0(n34497), .A1(n43042), .B0(n34481), .B1(n42451), .Y(
        n19422) );
  OR4X1 U55057 ( .A(n19413), .B(n19414), .C(n19415), .D(n19416), .Y(n36613) );
  OAI222XL U55058 ( .A0(n49531), .A1(n19417), .B0(n42508), .B1(n50128), .C0(
        n49539), .C1(n19419), .Y(n19415) );
  OAI22XL U55059 ( .A0(n42464), .A1(n43038), .B0(n36853), .B1(n42454), .Y(
        n19416) );
  OAI22XL U55060 ( .A0(n34498), .A1(n43042), .B0(n34482), .B1(n42451), .Y(
        n19414) );
  OR4X1 U55061 ( .A(n19483), .B(n19484), .C(n19485), .D(n19486), .Y(n36628) );
  OAI222XL U55062 ( .A0(n49524), .A1(n19456), .B0(n34443), .B1(n19457), .C0(
        n42584), .C1(n42453), .Y(n19485) );
  OAI22XL U55063 ( .A0(n49532), .A1(n42730), .B0(n36779), .B1(n43039), .Y(
        n19486) );
  OAI22XL U55064 ( .A0(n34483), .A1(n43041), .B0(n36771), .B1(n42451), .Y(
        n19484) );
  OR4X1 U55065 ( .A(n19479), .B(n19480), .C(n19481), .D(n19482), .Y(n36627) );
  OAI222XL U55066 ( .A0(n49525), .A1(n19456), .B0(n36907), .B1(n19457), .C0(
        n42569), .C1(n42452), .Y(n19481) );
  OAI22XL U55067 ( .A0(n49533), .A1(n42730), .B0(n36840), .B1(n43040), .Y(
        n19482) );
  OAI22XL U55068 ( .A0(n34484), .A1(n43041), .B0(n36736), .B1(n42451), .Y(
        n19480) );
  OR4X1 U55069 ( .A(n19475), .B(n19476), .C(n19477), .D(n19478), .Y(n36626) );
  OAI222XL U55070 ( .A0(n49526), .A1(n19456), .B0(n42663), .B1(n19457), .C0(
        n36801), .C1(n42453), .Y(n19477) );
  OAI22XL U55071 ( .A0(n49534), .A1(n42730), .B0(n36810), .B1(n43040), .Y(
        n19478) );
  OAI22XL U55072 ( .A0(n34485), .A1(n43041), .B0(n42479), .B1(n42450), .Y(
        n19476) );
  OR4X1 U55073 ( .A(n19471), .B(n19472), .C(n19473), .D(n19474), .Y(n36625) );
  OAI222XL U55074 ( .A0(n49527), .A1(n19456), .B0(n42644), .B1(n19457), .C0(
        n36827), .C1(n42452), .Y(n19473) );
  OAI22XL U55075 ( .A0(n49535), .A1(n42730), .B0(n41302), .B1(n43040), .Y(
        n19474) );
  OAI22XL U55076 ( .A0(n34486), .A1(n43041), .B0(n36747), .B1(n42450), .Y(
        n19472) );
  OR4X1 U55077 ( .A(n19467), .B(n19468), .C(n19469), .D(n19470), .Y(n36624) );
  OAI222XL U55078 ( .A0(n49528), .A1(n19456), .B0(n42633), .B1(n19457), .C0(
        n42554), .C1(n42452), .Y(n19469) );
  OAI22XL U55079 ( .A0(n49536), .A1(n42730), .B0(n41330), .B1(n43040), .Y(
        n19470) );
  OAI22XL U55080 ( .A0(n34487), .A1(n43041), .B0(n36714), .B1(n42450), .Y(
        n19468) );
  OR4X1 U55081 ( .A(n19463), .B(n19464), .C(n19465), .D(n19466), .Y(n36623) );
  OAI222XL U55082 ( .A0(n49529), .A1(n19456), .B0(n42620), .B1(n19457), .C0(
        n42544), .C1(n42453), .Y(n19465) );
  OAI22XL U55083 ( .A0(n49537), .A1(n42730), .B0(n41292), .B1(n43040), .Y(
        n19466) );
  OAI22XL U55084 ( .A0(n34488), .A1(n43042), .B0(n36795), .B1(n42451), .Y(
        n19464) );
  OR4X1 U55085 ( .A(n19459), .B(n19460), .C(n19461), .D(n19462), .Y(n36622) );
  OAI222XL U55086 ( .A0(n49530), .A1(n19456), .B0(n42609), .B1(n19457), .C0(
        n42517), .C1(n42452), .Y(n19461) );
  OAI22XL U55087 ( .A0(n49538), .A1(n42730), .B0(n41316), .B1(n43040), .Y(
        n19462) );
  OAI22XL U55088 ( .A0(n34489), .A1(n43042), .B0(n36757), .B1(n42451), .Y(
        n19460) );
  OR4X1 U55089 ( .A(n19452), .B(n19453), .C(n19454), .D(n19455), .Y(n36621) );
  OAI222XL U55090 ( .A0(n49531), .A1(n19456), .B0(n42592), .B1(n19457), .C0(
        n42508), .C1(n42453), .Y(n19454) );
  OAI22XL U55091 ( .A0(n49539), .A1(n42730), .B0(n36858), .B1(n43040), .Y(
        n19455) );
  OAI22XL U55092 ( .A0(n34490), .A1(n43042), .B0(n42463), .B1(n42450), .Y(
        n19453) );
  OR4X1 U55093 ( .A(n19498), .B(n19499), .C(n19500), .D(n19501), .Y(n36631) );
  OAI222XL U55094 ( .A0(n49545), .A1(n41797), .B0(n49529), .B1(n42729), .C0(
        n49537), .C1(n42728), .Y(n19500) );
  OAI22XL U55095 ( .A0(n36868), .A1(n42452), .B0(n40039), .B1(n19492), .Y(
        n19501) );
  OAI22XL U55096 ( .A0(n34480), .A1(n43041), .B0(n41291), .B1(n42450), .Y(
        n19499) );
  OR4X1 U55097 ( .A(n19494), .B(n19495), .C(n19496), .D(n19497), .Y(n36630) );
  OAI222XL U55098 ( .A0(n49546), .A1(n41797), .B0(n49530), .B1(n42729), .C0(
        n49538), .C1(n42728), .Y(n19496) );
  OAI22XL U55099 ( .A0(n42600), .A1(n42452), .B0(n36893), .B1(n19492), .Y(
        n19497) );
  OAI22XL U55100 ( .A0(n34481), .A1(n43041), .B0(n41310), .B1(n42451), .Y(
        n19495) );
  OR4X1 U55101 ( .A(n19488), .B(n19489), .C(n19490), .D(n19491), .Y(n36629) );
  OAI222XL U55102 ( .A0(n49547), .A1(n41797), .B0(n49531), .B1(n42729), .C0(
        n49539), .C1(n42728), .Y(n19490) );
  OAI22XL U55103 ( .A0(n42591), .A1(n42453), .B0(net219442), .B1(n19492), .Y(
        n19491) );
  OAI22XL U55104 ( .A0(n34482), .A1(n43041), .B0(n36854), .B1(n42450), .Y(
        n19489) );
  OR4X1 U55105 ( .A(n19407), .B(n19408), .C(n19409), .D(n19410), .Y(n36612) );
  OAI222XL U55106 ( .A0(n49540), .A1(n37183), .B0(n49524), .B1(n37525), .C0(
        n49532), .C1(n42731), .Y(n19409) );
  OAI22XL U55107 ( .A0(n36772), .A1(n42453), .B0(n36784), .B1(n19381), .Y(
        n19410) );
  OAI22XL U55108 ( .A0(n34499), .A1(n43042), .B0(n34483), .B1(n42451), .Y(
        n19408) );
  OR4X1 U55109 ( .A(n19403), .B(n19404), .C(n19405), .D(n19406), .Y(n36611) );
  OAI222XL U55110 ( .A0(n49541), .A1(n37183), .B0(n49525), .B1(n42732), .C0(
        n49533), .C1(n42731), .Y(n19405) );
  OAI22XL U55111 ( .A0(n36733), .A1(n42453), .B0(n36845), .B1(n19381), .Y(
        n19406) );
  OAI22XL U55112 ( .A0(n34500), .A1(n43042), .B0(n34484), .B1(n42451), .Y(
        n19404) );
  OR4X1 U55113 ( .A(n19399), .B(n19400), .C(n19401), .D(n19402), .Y(n36610) );
  OAI222XL U55114 ( .A0(n49542), .A1(n37183), .B0(n49526), .B1(n37525), .C0(
        n49534), .C1(n42731), .Y(n19401) );
  OAI22XL U55115 ( .A0(n42479), .A1(n42453), .B0(n36816), .B1(n19381), .Y(
        n19402) );
  OAI22XL U55116 ( .A0(n34501), .A1(n43042), .B0(n34485), .B1(n42451), .Y(
        n19400) );
  OR4X1 U55117 ( .A(n19395), .B(n19396), .C(n19397), .D(n19398), .Y(n36609) );
  OAI222XL U55118 ( .A0(n49543), .A1(n37183), .B0(n49527), .B1(n42732), .C0(
        n49535), .C1(n42731), .Y(n19397) );
  OAI22XL U55119 ( .A0(n36743), .A1(n42453), .B0(n41305), .B1(n19381), .Y(
        n19398) );
  OAI22XL U55120 ( .A0(n34502), .A1(n43042), .B0(n34486), .B1(n42451), .Y(
        n19396) );
  OR4X1 U55121 ( .A(n19391), .B(n19392), .C(n19393), .D(n19394), .Y(n36608) );
  OAI222XL U55122 ( .A0(n49544), .A1(n37183), .B0(n49528), .B1(n42732), .C0(
        n49536), .C1(n42731), .Y(n19393) );
  OAI22XL U55123 ( .A0(n36715), .A1(n42453), .B0(n41327), .B1(n19381), .Y(
        n19394) );
  OAI22XL U55124 ( .A0(n34503), .A1(n43042), .B0(n34487), .B1(n42451), .Y(
        n19392) );
  OR4X1 U55125 ( .A(n19387), .B(n19388), .C(n19389), .D(n19390), .Y(n36607) );
  OAI222XL U55126 ( .A0(n49545), .A1(n37183), .B0(n49529), .B1(n42732), .C0(
        n49537), .C1(n19292), .Y(n19389) );
  OAI22XL U55127 ( .A0(n36797), .A1(n42453), .B0(n41294), .B1(n19381), .Y(
        n19390) );
  OAI22XL U55128 ( .A0(n34504), .A1(n43042), .B0(n34488), .B1(n42451), .Y(
        n19388) );
  OR4X1 U55129 ( .A(n19383), .B(n19384), .C(n19385), .D(n19386), .Y(n36606) );
  OAI222XL U55130 ( .A0(n49546), .A1(n37183), .B0(n49530), .B1(n42732), .C0(
        n49538), .C1(n42731), .Y(n19385) );
  OAI22XL U55131 ( .A0(n36760), .A1(n42453), .B0(n41317), .B1(n19381), .Y(
        n19386) );
  OAI22XL U55132 ( .A0(n34505), .A1(n43042), .B0(n34489), .B1(n42451), .Y(
        n19384) );
  OR4X1 U55133 ( .A(n19377), .B(n19378), .C(n19379), .D(n19380), .Y(n36605) );
  OAI222XL U55134 ( .A0(n49547), .A1(n37183), .B0(n49531), .B1(n42732), .C0(
        n49539), .C1(n42731), .Y(n19379) );
  OAI22XL U55135 ( .A0(n42460), .A1(n42453), .B0(n36857), .B1(n19381), .Y(
        n19380) );
  OAI22XL U55136 ( .A0(n34506), .A1(n43042), .B0(n34490), .B1(n42451), .Y(
        n19378) );
  OR4X1 U55137 ( .A(n19518), .B(n19519), .C(n19520), .D(n19521), .Y(n36636) );
  OAI222XL U55138 ( .A0(n49540), .A1(n41797), .B0(n49524), .B1(n42729), .C0(
        n49532), .C1(n42728), .Y(n19520) );
  OAI22XL U55139 ( .A0(n36903), .A1(n42452), .B0(n42723), .B1(n19492), .Y(
        n19521) );
  OAI22XL U55140 ( .A0(n34475), .A1(n43041), .B0(n36780), .B1(n42451), .Y(
        n19519) );
  OR4X1 U55141 ( .A(n19293), .B(n19294), .C(n19295), .D(n19296), .Y(n36590) );
  OAI22XL U55142 ( .A0(n49530), .A1(n50130), .B0(n49538), .B1(n50140), .Y(
        n19296) );
  OAI22XL U55143 ( .A0(n49546), .A1(n42732), .B0(n34481), .B1(n19290), .Y(
        n19295) );
  OAI22XL U55144 ( .A0(n49554), .A1(n42731), .B0(n34505), .B1(n37241), .Y(
        n19294) );
  OR4X1 U55145 ( .A(n19299), .B(n19300), .C(n19301), .D(n19302), .Y(n36591) );
  OAI22XL U55146 ( .A0(n49529), .A1(n50130), .B0(n49537), .B1(n50140), .Y(
        n19302) );
  OAI22XL U55147 ( .A0(n49545), .A1(n42732), .B0(n34480), .B1(n19290), .Y(
        n19301) );
  OAI22XL U55148 ( .A0(n49553), .A1(n42731), .B0(n34504), .B1(n37241), .Y(
        n19300) );
  OR4X1 U55149 ( .A(n19305), .B(n19306), .C(n19307), .D(n19308), .Y(n36592) );
  OAI22XL U55150 ( .A0(n49528), .A1(n50130), .B0(n49536), .B1(n50140), .Y(
        n19308) );
  OAI22XL U55151 ( .A0(n49544), .A1(n42732), .B0(n34479), .B1(n19290), .Y(
        n19307) );
  OAI22XL U55152 ( .A0(n49552), .A1(n42731), .B0(n34503), .B1(n37241), .Y(
        n19306) );
  OR4X1 U55153 ( .A(n19311), .B(n19312), .C(n19313), .D(n19314), .Y(n36593) );
  OAI22XL U55154 ( .A0(n49527), .A1(n50130), .B0(n49535), .B1(n50140), .Y(
        n19314) );
  OAI22XL U55155 ( .A0(n49543), .A1(n42732), .B0(n34478), .B1(n19290), .Y(
        n19313) );
  OAI22XL U55156 ( .A0(n49551), .A1(n42731), .B0(n34502), .B1(n37241), .Y(
        n19312) );
  OR4X1 U55157 ( .A(n19317), .B(n19318), .C(n19319), .D(n19320), .Y(n36594) );
  OAI22XL U55158 ( .A0(n49526), .A1(n50130), .B0(n49534), .B1(n50140), .Y(
        n19320) );
  OAI22XL U55159 ( .A0(n49542), .A1(n42732), .B0(n34477), .B1(n19290), .Y(
        n19319) );
  OAI22XL U55160 ( .A0(n49550), .A1(n42731), .B0(n34501), .B1(n37241), .Y(
        n19318) );
  OR4X1 U55161 ( .A(n19323), .B(n19324), .C(n19325), .D(n19326), .Y(n36595) );
  OAI22XL U55162 ( .A0(n49525), .A1(n50130), .B0(n49533), .B1(n50140), .Y(
        n19326) );
  OAI22XL U55163 ( .A0(n49541), .A1(n42732), .B0(n34476), .B1(n19290), .Y(
        n19325) );
  OAI22XL U55164 ( .A0(n49549), .A1(n42731), .B0(n34500), .B1(n37241), .Y(
        n19324) );
  OR4X1 U55165 ( .A(n19329), .B(n19330), .C(n19331), .D(n19332), .Y(n36596) );
  OAI22XL U55166 ( .A0(n49524), .A1(n50130), .B0(n49532), .B1(n50140), .Y(
        n19332) );
  OAI22XL U55167 ( .A0(n49540), .A1(n42732), .B0(n34475), .B1(n19290), .Y(
        n19331) );
  OAI22XL U55168 ( .A0(n49548), .A1(n42731), .B0(n34499), .B1(n37241), .Y(
        n19330) );
  OR4X1 U55169 ( .A(n19284), .B(n19285), .C(n19286), .D(n19287), .Y(n36589) );
  OAI22XL U55170 ( .A0(n49531), .A1(n50130), .B0(n50140), .B1(n49539), .Y(
        n19287) );
  OAI22XL U55171 ( .A0(n49547), .A1(n42732), .B0(n34482), .B1(n19290), .Y(
        n19286) );
  OAI22XL U55172 ( .A0(n49555), .A1(n42731), .B0(n34506), .B1(n37241), .Y(
        n19285) );
  NAND2X1 U55173 ( .A(n32399), .B(n42316), .Y(n9734) );
  AO22X1 U55174 ( .A0(N23551), .A1(out_valid), .B0(enc_num[0]), .B1(n41791),
        .Y(n32394) );
  AO22X1 U55175 ( .A0(N23560), .A1(out_valid), .B0(enc_num[9]), .B1(n41791),
        .Y(n32385) );
  AO22X1 U55176 ( .A0(N23559), .A1(out_valid), .B0(enc_num[8]), .B1(n41791),
        .Y(n32386) );
  AO22X1 U55177 ( .A0(N23558), .A1(out_valid), .B0(enc_num[7]), .B1(n41791),
        .Y(n32387) );
  AO22X1 U55178 ( .A0(N23557), .A1(out_valid), .B0(enc_num[6]), .B1(n41791),
        .Y(n32388) );
  AO22X1 U55179 ( .A0(N23556), .A1(out_valid), .B0(enc_num[5]), .B1(n41791),
        .Y(n32389) );
  AO22X1 U55180 ( .A0(N23555), .A1(out_valid), .B0(enc_num[4]), .B1(n41791),
        .Y(n32390) );
  AO22X1 U55181 ( .A0(N23554), .A1(out_valid), .B0(enc_num[3]), .B1(n41791),
        .Y(n32391) );
  AO22X1 U55182 ( .A0(N23553), .A1(out_valid), .B0(enc_num[2]), .B1(n41791),
        .Y(n32392) );
  AO22X1 U55183 ( .A0(N23552), .A1(out_valid), .B0(enc_num[1]), .B1(n41791),
        .Y(n32393) );
  CLKBUFX3 U55184 ( .A(n32400), .Y(n42316) );
  NOR2X2 U55185 ( .A(n32399), .B(n42316), .Y(n9715) );
  OAI221XL U55186 ( .A0(n34505), .A1(n19181), .B0(n19182), .B1(n49530), .C0(
        n19199), .Y(n36572) );
  AOI222XL U55187 ( .A0(data[9]), .A1(n19185), .B0(data[1]), .B1(n19186), .C0(
        data[17]), .C1(n19187), .Y(n19199) );
  OAI221XL U55188 ( .A0(n34504), .A1(n19181), .B0(n19182), .B1(n49529), .C0(
        n19197), .Y(n36571) );
  AOI222XL U55189 ( .A0(data[10]), .A1(n19185), .B0(data[2]), .B1(n19186),
        .C0(data[18]), .C1(n19187), .Y(n19197) );
  OAI221XL U55190 ( .A0(n34503), .A1(n19181), .B0(n19182), .B1(n49528), .C0(
        n19195), .Y(n36570) );
  AOI222XL U55191 ( .A0(data[11]), .A1(n19185), .B0(data[3]), .B1(n19186),
        .C0(data[19]), .C1(n19187), .Y(n19195) );
  OAI221XL U55192 ( .A0(n34502), .A1(n19181), .B0(n19182), .B1(n49527), .C0(
        n19193), .Y(n36569) );
  AOI222XL U55193 ( .A0(data[12]), .A1(n19185), .B0(data[4]), .B1(n19186),
        .C0(data[20]), .C1(n19187), .Y(n19193) );
  OAI221XL U55194 ( .A0(n34501), .A1(n19181), .B0(n19182), .B1(n49526), .C0(
        n19191), .Y(n36568) );
  AOI222XL U55195 ( .A0(data[13]), .A1(n19185), .B0(data[5]), .B1(n19186),
        .C0(data[21]), .C1(n19187), .Y(n19191) );
  OAI221XL U55196 ( .A0(n34500), .A1(n19181), .B0(n19182), .B1(n49525), .C0(
        n19189), .Y(n36567) );
  AOI222XL U55197 ( .A0(data[14]), .A1(n19185), .B0(data[6]), .B1(n19186),
        .C0(data[22]), .C1(n19187), .Y(n19189) );
  OAI221XL U55198 ( .A0(n34499), .A1(n19181), .B0(n19182), .B1(n49524), .C0(
        n19184), .Y(n36566) );
  AOI222XL U55199 ( .A0(data[15]), .A1(n19185), .B0(data[7]), .B1(n19186),
        .C0(data[23]), .C1(n19187), .Y(n19184) );
  OAI221XL U55200 ( .A0(n34506), .A1(n19181), .B0(n19182), .B1(n49531), .C0(
        n32367), .Y(n36637) );
  AOI222XL U55201 ( .A0(data[8]), .A1(n19185), .B0(data[0]), .B1(n19186), .C0(
        data[16]), .C1(n19187), .Y(n32367) );
  INVX3 U55202 ( .A(data[25]), .Y(n49530) );
  INVX3 U55203 ( .A(data[26]), .Y(n49529) );
  INVX3 U55204 ( .A(data[27]), .Y(n49528) );
  INVX3 U55205 ( .A(data[28]), .Y(n49527) );
  INVX3 U55206 ( .A(data[29]), .Y(n49526) );
  INVX3 U55207 ( .A(data[30]), .Y(n49525) );
  INVX3 U55208 ( .A(data[31]), .Y(n49524) );
  INVX3 U55209 ( .A(data[24]), .Y(n49531) );
  INVX3 U55210 ( .A(data[9]), .Y(n49546) );
  INVX3 U55211 ( .A(data[10]), .Y(n49545) );
  INVX3 U55212 ( .A(data[11]), .Y(n49544) );
  INVX3 U55213 ( .A(data[12]), .Y(n49543) );
  INVX3 U55214 ( .A(data[13]), .Y(n49542) );
  INVX3 U55215 ( .A(data[14]), .Y(n49541) );
  INVX3 U55216 ( .A(data[15]), .Y(n49540) );
  OAI211X1 U55217 ( .A0(n50130), .A1(n49547), .B0(n19202), .C0(n19203), .Y(
        n36573) );
  AOI222XL U55218 ( .A0(n41736), .A1(n49557), .B0(data[0]), .B1(n37182), .C0(
        data[16]), .C1(n37520), .Y(n19203) );
  AOI2BB2X1 U55219 ( .B0(data[24]), .B1(n19207), .A0N(n34498), .A1N(n19208),
        .Y(n19202) );
  INVX3 U55220 ( .A(data[8]), .Y(n49547) );
  OAI211X1 U55221 ( .A0(n9679), .A1(n9680), .B0(n9681), .C0(n9682), .Y(
        nxt_state[1]) );
  OAI21XL U55222 ( .A0(n50134), .A1(n50146), .B0(n9689), .Y(n9681) );
  AOI2BB2X1 U55223 ( .B0(n9690), .B1(n50143), .A0N(n49556), .A1N(n50149), .Y(
        n9680) );
  NOR3X1 U55224 ( .A(n50147), .B(n32397), .C(n9734), .Y(n32369) );
  NAND2X1 U55225 ( .A(n9651), .B(data_valid), .Y(n9690) );
  OAI21XL U55226 ( .A0(n32398), .A1(n50141), .B0(n32397), .Y(n9683) );
  OAI211X1 U55227 ( .A0(n49546), .A1(n50130), .B0(n19210), .C0(n19211), .Y(
        n36574) );
  AOI222XL U55228 ( .A0(n41736), .A1(n50163), .B0(n37182), .B1(data[1]), .C0(
        n37520), .C1(data[17]), .Y(n19211) );
  AOI2BB2X1 U55229 ( .B0(n19207), .B1(data[25]), .A0N(n34497), .A1N(n19208),
        .Y(n19210) );
  OAI211X1 U55230 ( .A0(n49545), .A1(n50130), .B0(n19214), .C0(n19215), .Y(
        n36575) );
  AOI222XL U55231 ( .A0(n41736), .A1(n50161), .B0(n37182), .B1(data[2]), .C0(
        n37520), .C1(data[18]), .Y(n19215) );
  AOI2BB2X1 U55232 ( .B0(n19207), .B1(data[26]), .A0N(n34496), .A1N(n19208),
        .Y(n19214) );
  OAI211X1 U55233 ( .A0(n49544), .A1(n50130), .B0(n19218), .C0(n19219), .Y(
        n36576) );
  AOI222XL U55234 ( .A0(n41736), .A1(n50159), .B0(n37182), .B1(data[3]), .C0(
        n37520), .C1(data[19]), .Y(n19219) );
  AOI2BB2X1 U55235 ( .B0(n19207), .B1(data[27]), .A0N(n34495), .A1N(n19208),
        .Y(n19218) );
  OAI211X1 U55236 ( .A0(n49543), .A1(n50130), .B0(n19222), .C0(n19223), .Y(
        n36577) );
  AOI222XL U55237 ( .A0(n41736), .A1(n50157), .B0(n37182), .B1(data[4]), .C0(
        n37520), .C1(data[20]), .Y(n19223) );
  AOI2BB2X1 U55238 ( .B0(n19207), .B1(data[28]), .A0N(n34494), .A1N(n19208),
        .Y(n19222) );
  OAI211X1 U55239 ( .A0(n49542), .A1(n50130), .B0(n19226), .C0(n19227), .Y(
        n36578) );
  AOI222XL U55240 ( .A0(n41736), .A1(n50155), .B0(n37182), .B1(data[5]), .C0(
        n37520), .C1(data[21]), .Y(n19227) );
  AOI2BB2X1 U55241 ( .B0(n19207), .B1(data[29]), .A0N(n34493), .A1N(n19208),
        .Y(n19226) );
  OAI211X1 U55242 ( .A0(n49541), .A1(n50130), .B0(n19230), .C0(n19231), .Y(
        n36579) );
  AOI222XL U55243 ( .A0(n41736), .A1(n50153), .B0(n37182), .B1(data[6]), .C0(
        n37520), .C1(data[22]), .Y(n19231) );
  AOI2BB2X1 U55244 ( .B0(n19207), .B1(data[30]), .A0N(n34492), .A1N(n19208),
        .Y(n19230) );
  OAI211X1 U55245 ( .A0(n49540), .A1(n50130), .B0(n19234), .C0(n19235), .Y(
        n36580) );
  AOI222XL U55246 ( .A0(n41736), .A1(n50151), .B0(n37182), .B1(data[7]), .C0(
        n37520), .C1(data[23]), .Y(n19235) );
  AOI2BB2X1 U55247 ( .B0(n19207), .B1(data[31]), .A0N(n34491), .A1N(n19208),
        .Y(n19234) );
  CLKINVX1 U55248 ( .A(drop_done), .Y(n49556) );
  NOR3X1 U55249 ( .A(net209923), .B(net256309), .C(net210441), .Y(n47808) );
  NAND2X1 U55250 ( .A(n48305), .B(n47727), .Y(n47728) );
  OAI21XL U55251 ( .A0(n48306), .A1(net209615), .B0(n48305), .Y(n48308) );
  NAND2BX1 U55252 ( .AN(net210554), .B(net210553), .Y(n47799) );
  NAND4XL U55253 ( .A(net213675), .B(n45528), .C(n41752), .D(net210477), .Y(
        n47840) );
  AOI211XL U55254 ( .A0(net209307), .A1(net209308), .B0(n48451), .C0(net209310), .Y(n48452) );
  NOR2X4 U55255 ( .A(n45512), .B(net209604), .Y(net213700) );
  OAI211XL U55256 ( .A0(net209315), .A1(net209316), .B0(net209308), .C0(
        net209317), .Y(n48453) );
  OAI21XL U55257 ( .A0(net209634), .A1(net209635), .B0(net209636), .Y(n48298)
         );
  INVX2 U55258 ( .A(net209902), .Y(net209901) );
  OAI21XL U55259 ( .A0(net209342), .A1(net209343), .B0(net209344), .Y(n48434)
         );
  AOI21XL U55260 ( .A0(n48434), .A1(net209313), .B0(n48433), .Y(n48459) );
  NAND3BXL U55261 ( .AN(net210442), .B(net210443), .C(net209900), .Y(n47809)
         );
  AOI21XL U55262 ( .A0(n48144), .A1(n48143), .B0(n48142), .Y(n48155) );
  CLKINVX2 U55263 ( .A(n43010), .Y(n42736) );
  CLKINVX2 U55264 ( .A(n43010), .Y(n42739) );
  CLKINVX2 U55265 ( .A(n43009), .Y(n42740) );
  CLKINVX2 U55266 ( .A(n43020), .Y(n42741) );
  CLKINVX2 U55267 ( .A(n43017), .Y(n42742) );
  CLKINVX2 U55268 ( .A(n43017), .Y(n42743) );
  CLKINVX2 U55269 ( .A(n43017), .Y(n42744) );
  CLKINVX2 U55270 ( .A(n43017), .Y(n42745) );
  CLKINVX2 U55271 ( .A(n43017), .Y(n42746) );
  CLKINVX2 U55272 ( .A(n43017), .Y(n42747) );
  CLKINVX2 U55273 ( .A(n43017), .Y(n42748) );
  CLKINVX2 U55274 ( .A(n43017), .Y(n42749) );
  CLKINVX2 U55275 ( .A(n43017), .Y(n42751) );
  CLKINVX2 U55276 ( .A(n43017), .Y(n42752) );
  CLKINVX2 U55277 ( .A(n43017), .Y(n42754) );
  CLKINVX2 U55278 ( .A(n43017), .Y(n42755) );
  CLKINVX2 U55279 ( .A(n43017), .Y(n42756) );
  CLKINVX2 U55280 ( .A(n43018), .Y(n42757) );
  CLKINVX2 U55281 ( .A(n43018), .Y(n42758) );
  CLKINVX2 U55282 ( .A(n43018), .Y(n42759) );
  CLKINVX2 U55283 ( .A(n43018), .Y(n42760) );
  CLKINVX2 U55284 ( .A(n43018), .Y(n42761) );
  CLKINVX2 U55285 ( .A(n43018), .Y(n42762) );
  CLKINVX2 U55286 ( .A(n43018), .Y(n42764) );
  CLKINVX2 U55287 ( .A(n43018), .Y(n42765) );
  CLKINVX2 U55288 ( .A(n43018), .Y(n42766) );
  CLKINVX2 U55289 ( .A(n43018), .Y(n42767) );
  CLKINVX2 U55290 ( .A(n43018), .Y(n42768) );
  CLKINVX2 U55291 ( .A(n43018), .Y(n42770) );
  CLKINVX2 U55292 ( .A(n43018), .Y(n42771) );
  CLKINVX2 U55293 ( .A(n43018), .Y(n42772) );
  CLKINVX2 U55294 ( .A(n43018), .Y(n42773) );
  CLKINVX2 U55295 ( .A(n43018), .Y(n42774) );
  CLKINVX2 U55296 ( .A(n43019), .Y(n42776) );
  CLKINVX2 U55297 ( .A(n43019), .Y(n42777) );
  CLKINVX2 U55298 ( .A(n43019), .Y(n42778) );
  CLKINVX2 U55299 ( .A(n43019), .Y(n42780) );
  CLKINVX2 U55300 ( .A(n43019), .Y(n42781) );
  CLKINVX2 U55301 ( .A(n43019), .Y(n42782) );
  CLKINVX2 U55302 ( .A(n43019), .Y(n42783) );
  CLKINVX2 U55303 ( .A(n43019), .Y(n42785) );
  CLKINVX2 U55304 ( .A(n43019), .Y(n42786) );
  CLKINVX2 U55305 ( .A(n43019), .Y(n42787) );
  CLKINVX2 U55306 ( .A(n43019), .Y(n42788) );
  CLKINVX2 U55307 ( .A(n43019), .Y(n42789) );
  CLKINVX2 U55308 ( .A(n43019), .Y(n42790) );
  CLKINVX2 U55309 ( .A(n43019), .Y(n42791) );
  CLKINVX2 U55310 ( .A(n43019), .Y(n42792) );
  CLKINVX2 U55311 ( .A(n43020), .Y(n42793) );
  CLKINVX2 U55312 ( .A(n43020), .Y(n42794) );
  CLKINVX2 U55313 ( .A(n43020), .Y(n42795) );
  CLKINVX2 U55314 ( .A(n43020), .Y(n42796) );
  CLKINVX2 U55315 ( .A(n43020), .Y(n42797) );
  CLKINVX2 U55316 ( .A(n43020), .Y(n42798) );
  CLKINVX2 U55317 ( .A(n43020), .Y(n42799) );
  CLKINVX2 U55318 ( .A(n43020), .Y(n42800) );
  CLKINVX2 U55319 ( .A(n43020), .Y(n42801) );
  CLKINVX2 U55320 ( .A(n43020), .Y(n42802) );
  CLKINVX2 U55321 ( .A(n43020), .Y(n42803) );
  CLKINVX2 U55322 ( .A(n43020), .Y(n42804) );
  CLKINVX2 U55323 ( .A(n43020), .Y(n42806) );
  CLKINVX2 U55324 ( .A(n43020), .Y(n42807) );
  CLKINVX2 U55325 ( .A(n43020), .Y(n42808) );
  CLKINVX2 U55326 ( .A(n43020), .Y(n42809) );
  CLKINVX2 U55327 ( .A(n43021), .Y(n42812) );
  CLKINVX2 U55328 ( .A(n43021), .Y(n42813) );
  CLKINVX2 U55329 ( .A(n43021), .Y(n42814) );
  CLKINVX2 U55330 ( .A(n43021), .Y(n42815) );
  CLKINVX2 U55331 ( .A(n43021), .Y(n42816) );
  CLKINVX2 U55332 ( .A(n43021), .Y(n42817) );
  CLKINVX2 U55333 ( .A(n43021), .Y(n42818) );
  CLKINVX2 U55334 ( .A(n43021), .Y(n42819) );
  CLKINVX2 U55335 ( .A(n43021), .Y(n42820) );
  CLKINVX2 U55336 ( .A(n43021), .Y(n42821) );
  CLKINVX2 U55337 ( .A(n43021), .Y(n42822) );
  CLKINVX2 U55338 ( .A(n43021), .Y(n42823) );
  CLKINVX2 U55339 ( .A(n43021), .Y(n42824) );
  CLKINVX2 U55340 ( .A(n43021), .Y(n42825) );
  CLKINVX2 U55341 ( .A(n43021), .Y(n42826) );
  CLKINVX2 U55342 ( .A(n43021), .Y(n42827) );
  CLKINVX2 U55343 ( .A(n43022), .Y(n42828) );
  CLKINVX2 U55344 ( .A(n43022), .Y(n42829) );
  CLKINVX2 U55345 ( .A(n43022), .Y(n42830) );
  CLKINVX2 U55346 ( .A(n43022), .Y(n42831) );
  CLKINVX2 U55347 ( .A(n43022), .Y(n42832) );
  CLKINVX2 U55348 ( .A(n43022), .Y(n42833) );
  CLKINVX2 U55349 ( .A(n43022), .Y(n42834) );
  CLKINVX2 U55350 ( .A(n43022), .Y(n42835) );
  CLKINVX2 U55351 ( .A(n43022), .Y(n42836) );
  CLKINVX2 U55352 ( .A(n43022), .Y(n42837) );
  CLKINVX2 U55353 ( .A(n43022), .Y(n42838) );
  CLKINVX2 U55354 ( .A(n43022), .Y(n42839) );
  CLKINVX2 U55355 ( .A(n43022), .Y(n42840) );
  CLKINVX2 U55356 ( .A(n43022), .Y(n42841) );
  CLKINVX2 U55357 ( .A(n43022), .Y(n42842) );
  CLKINVX2 U55358 ( .A(n43022), .Y(n42843) );
  CLKINVX2 U55359 ( .A(n43022), .Y(n42844) );
  CLKINVX2 U55360 ( .A(n43023), .Y(n42847) );
  CLKINVX2 U55361 ( .A(n43023), .Y(n42848) );
  CLKINVX2 U55362 ( .A(n43023), .Y(n42849) );
  CLKINVX2 U55363 ( .A(n43023), .Y(n42850) );
  CLKINVX2 U55364 ( .A(n43023), .Y(n42851) );
  CLKINVX2 U55365 ( .A(n43023), .Y(n42852) );
  CLKINVX2 U55366 ( .A(n43023), .Y(n42853) );
  CLKINVX2 U55367 ( .A(n43023), .Y(n42854) );
  CLKINVX2 U55368 ( .A(n43023), .Y(n42855) );
  CLKINVX2 U55369 ( .A(n43023), .Y(n42856) );
  CLKINVX2 U55370 ( .A(n43023), .Y(n42857) );
  CLKINVX2 U55371 ( .A(n43023), .Y(n42858) );
  CLKINVX2 U55372 ( .A(n43023), .Y(n42859) );
  CLKINVX2 U55373 ( .A(n43023), .Y(n42862) );
  CLKINVX2 U55374 ( .A(n43023), .Y(n42863) );
  CLKINVX2 U55375 ( .A(n43032), .Y(n42864) );
  CLKINVX2 U55376 ( .A(n43009), .Y(n42865) );
  CLKINVX2 U55377 ( .A(n43013), .Y(n42866) );
  CLKINVX2 U55378 ( .A(n43010), .Y(n42867) );
  CLKINVX2 U55379 ( .A(n43010), .Y(n42868) );
  CLKINVX2 U55380 ( .A(n43010), .Y(n42869) );
  CLKINVX2 U55381 ( .A(n43010), .Y(n42870) );
  CLKINVX2 U55382 ( .A(n43010), .Y(n42871) );
  CLKINVX2 U55383 ( .A(n43010), .Y(n42872) );
  CLKINVX2 U55384 ( .A(n43010), .Y(n42873) );
  CLKINVX2 U55385 ( .A(n43010), .Y(n42874) );
  CLKINVX2 U55386 ( .A(n43010), .Y(n42875) );
  CLKINVX2 U55387 ( .A(n43010), .Y(n42876) );
  CLKINVX2 U55388 ( .A(n43010), .Y(n42877) );
  CLKINVX2 U55389 ( .A(n43010), .Y(n42878) );
  CLKINVX2 U55390 ( .A(n43010), .Y(n42879) );
  CLKINVX2 U55391 ( .A(n43010), .Y(n42880) );
  CLKINVX2 U55392 ( .A(n43011), .Y(n42881) );
  CLKINVX2 U55393 ( .A(n43011), .Y(n42882) );
  CLKINVX2 U55394 ( .A(n43011), .Y(n42883) );
  CLKINVX2 U55395 ( .A(n43011), .Y(n42884) );
  CLKINVX2 U55396 ( .A(n43011), .Y(n42885) );
  CLKINVX2 U55397 ( .A(n43011), .Y(n42886) );
  CLKINVX2 U55398 ( .A(n43011), .Y(n42887) );
  CLKINVX2 U55399 ( .A(n43011), .Y(n42888) );
  CLKINVX2 U55400 ( .A(n43011), .Y(n42889) );
  CLKINVX2 U55401 ( .A(n43011), .Y(n42890) );
  CLKINVX2 U55402 ( .A(n43011), .Y(n42891) );
  CLKINVX2 U55403 ( .A(n43011), .Y(n42892) );
  CLKINVX2 U55404 ( .A(n43011), .Y(n42893) );
  CLKINVX2 U55405 ( .A(n43011), .Y(n42894) );
  CLKINVX2 U55406 ( .A(n43011), .Y(n42895) );
  CLKINVX2 U55407 ( .A(n43011), .Y(n42896) );
  CLKINVX2 U55408 ( .A(n43011), .Y(n42897) );
  CLKINVX2 U55409 ( .A(n43011), .Y(n42898) );
  CLKINVX2 U55410 ( .A(n43012), .Y(n42899) );
  CLKINVX2 U55411 ( .A(n43012), .Y(n42900) );
  CLKINVX2 U55412 ( .A(n43012), .Y(n42901) );
  CLKINVX2 U55413 ( .A(n43012), .Y(n42902) );
  CLKINVX2 U55414 ( .A(n43012), .Y(n42903) );
  CLKINVX2 U55415 ( .A(n43012), .Y(n42904) );
  CLKINVX2 U55416 ( .A(n43012), .Y(n42905) );
  CLKINVX2 U55417 ( .A(n43012), .Y(n42906) );
  CLKINVX2 U55418 ( .A(n43012), .Y(n42907) );
  CLKINVX2 U55419 ( .A(n43012), .Y(n42908) );
  CLKINVX2 U55420 ( .A(n43012), .Y(n42910) );
  CLKINVX2 U55421 ( .A(n43012), .Y(n42911) );
  CLKINVX2 U55422 ( .A(n43012), .Y(n42912) );
  CLKINVX2 U55423 ( .A(n43012), .Y(n42913) );
  CLKINVX2 U55424 ( .A(n43012), .Y(n42914) );
  CLKINVX2 U55425 ( .A(n43012), .Y(n42915) );
  CLKINVX2 U55426 ( .A(n43012), .Y(n42916) );
  CLKINVX2 U55427 ( .A(n43013), .Y(n42917) );
  CLKINVX2 U55428 ( .A(n43013), .Y(n42918) );
  CLKINVX2 U55429 ( .A(n43013), .Y(n42919) );
  CLKINVX2 U55430 ( .A(n43013), .Y(n42920) );
  CLKINVX2 U55431 ( .A(n43013), .Y(n42921) );
  CLKINVX2 U55432 ( .A(n43013), .Y(n42922) );
  CLKINVX2 U55433 ( .A(n43013), .Y(n42923) );
  CLKINVX2 U55434 ( .A(n43013), .Y(n42924) );
  CLKINVX2 U55435 ( .A(n43013), .Y(n42925) );
  CLKINVX2 U55436 ( .A(n43013), .Y(n42926) );
  CLKINVX2 U55437 ( .A(n43013), .Y(n42927) );
  CLKINVX2 U55438 ( .A(n43013), .Y(n42928) );
  CLKINVX2 U55439 ( .A(n43013), .Y(n42929) );
  CLKINVX2 U55440 ( .A(n43013), .Y(n42930) );
  CLKINVX2 U55441 ( .A(n43013), .Y(n42931) );
  CLKINVX2 U55442 ( .A(n43013), .Y(n42932) );
  CLKINVX2 U55443 ( .A(n43013), .Y(n42933) );
  CLKINVX2 U55444 ( .A(n43014), .Y(n42934) );
  CLKINVX2 U55445 ( .A(n43014), .Y(n42935) );
  CLKINVX2 U55446 ( .A(n43014), .Y(n42936) );
  CLKINVX2 U55447 ( .A(n43014), .Y(n42937) );
  CLKINVX2 U55448 ( .A(n43014), .Y(n42938) );
  CLKINVX2 U55449 ( .A(n43014), .Y(n42939) );
  CLKINVX2 U55450 ( .A(n43014), .Y(n42940) );
  CLKINVX2 U55451 ( .A(n43014), .Y(n42941) );
  CLKINVX2 U55452 ( .A(n43014), .Y(n42942) );
  CLKINVX2 U55453 ( .A(n43014), .Y(n42943) );
  CLKINVX2 U55454 ( .A(n43014), .Y(n42944) );
  CLKINVX2 U55455 ( .A(n43014), .Y(n42945) );
  CLKINVX2 U55456 ( .A(n43014), .Y(n42946) );
  CLKINVX2 U55457 ( .A(n43014), .Y(n42947) );
  CLKINVX2 U55458 ( .A(n43014), .Y(n42948) );
  CLKINVX2 U55459 ( .A(n43014), .Y(n42949) );
  CLKINVX2 U55460 ( .A(n43015), .Y(n42952) );
  CLKINVX2 U55461 ( .A(n43015), .Y(n42953) );
  CLKINVX2 U55462 ( .A(n43015), .Y(n42954) );
  CLKINVX2 U55463 ( .A(n43015), .Y(n42955) );
  CLKINVX2 U55464 ( .A(n43015), .Y(n42958) );
  CLKINVX2 U55465 ( .A(n43015), .Y(n42959) );
  CLKINVX2 U55466 ( .A(n43015), .Y(n42960) );
  CLKINVX2 U55467 ( .A(n43015), .Y(n42961) );
  CLKINVX2 U55468 ( .A(n43015), .Y(n42962) );
  CLKINVX2 U55469 ( .A(n43015), .Y(n42963) );
  CLKINVX2 U55470 ( .A(n43015), .Y(n42964) );
  CLKINVX2 U55471 ( .A(n43015), .Y(n42965) );
  CLKINVX2 U55472 ( .A(n43015), .Y(n42966) );
  CLKINVX2 U55473 ( .A(n43015), .Y(n42967) );
  CLKINVX2 U55474 ( .A(n43015), .Y(n42968) );
  CLKINVX2 U55475 ( .A(n43015), .Y(n42969) );
  CLKINVX2 U55476 ( .A(n43016), .Y(n42970) );
  CLKINVX2 U55477 ( .A(n43016), .Y(n42971) );
  CLKINVX2 U55478 ( .A(n43016), .Y(n42972) );
  CLKINVX2 U55479 ( .A(n43016), .Y(n42973) );
  CLKINVX2 U55480 ( .A(n43016), .Y(n42974) );
  CLKINVX2 U55481 ( .A(n43016), .Y(n42975) );
  CLKINVX2 U55482 ( .A(n43016), .Y(n42976) );
  CLKINVX2 U55483 ( .A(n43016), .Y(n42977) );
  CLKINVX2 U55484 ( .A(n43016), .Y(n42978) );
  CLKINVX2 U55485 ( .A(n43016), .Y(n42979) );
  CLKINVX2 U55486 ( .A(n43016), .Y(n42980) );
  CLKINVX2 U55487 ( .A(n43016), .Y(n42981) );
  CLKINVX2 U55488 ( .A(n43016), .Y(n42982) );
  CLKINVX2 U55489 ( .A(n43016), .Y(n42983) );
  CLKINVX2 U55490 ( .A(n43016), .Y(n42984) );
  CLKINVX2 U55491 ( .A(n43016), .Y(n42985) );
  CLKINVX2 U55492 ( .A(n43016), .Y(n42986) );
  CLKINVX2 U55493 ( .A(n43016), .Y(n42987) );
  CLKINVX2 U55494 ( .A(n43017), .Y(n42988) );
  CLKINVX2 U55495 ( .A(n43017), .Y(n42989) );
  CLKINVX2 U55496 ( .A(n43017), .Y(n42990) );
  OAI21X4 U55497 ( .A0(n47783), .A1(net210548), .B0(n41764), .Y(n47784) );
  AOI21X4 U55498 ( .A0(n41763), .A1(n47784), .B0(net210544), .Y(n47787) );
  CLKINVX3 U55499 ( .A(n48133), .Y(n48134) );
endmodule

module CHIP(
  clk,
  reset,
  data,
  data_valid,
  drop_done,
  busy,
  codeword,
  enc_num,
  out_valid,
  finish
);

input         clk;
input         reset;
input  [31:0] data;
input         data_valid;
input         drop_done;
output        busy;
output [10:0] codeword;
output [11:0] enc_num;
output        out_valid;
output        finish;


wire          clk_i;
wire          reset_i;
wire   [31:0] data_i;
wire          data_valid_i;
wire          drop_done_i;
wire          busy_i;
wire   [10:0] codeword_i;
wire   [11:0] enc_num_i;
wire          out_valid_i;
wire          finish_i;


LZSS LZSS(  .clk(clk_i), .reset(reset_i), .data(data_i), .data_valid(data_valid_i), .drop_done(drop_done_i),
  .busy(busy_i), .codeword(codeword_i), .enc_num(enc_num_i),
  .out_valid(out_valid_i), .finish(finish_i)          );



PDIDGZ    ipad_clk( .PAD(clk),      .C(clk_i)  );
PDIDGZ    ipad_rst( .PAD(reset),      .C(reset_i)  );
PDIDGZ    ipad_val( .PAD(data_valid), .C(data_valid_i)  );
PDIDGZ    ipad_don( .PAD(drop_done),  .C(drop_done_i)  );
PDIDGZ    ipad_dat00( .PAD(data[0 ]), .C(data_i[0 ])  );
PDIDGZ    ipad_dat01( .PAD(data[1 ]), .C(data_i[1 ])  );
PDIDGZ    ipad_dat02( .PAD(data[2 ]), .C(data_i[2 ])  );
PDIDGZ    ipad_dat03( .PAD(data[3 ]), .C(data_i[3 ])  );
PDIDGZ    ipad_dat04( .PAD(data[4 ]), .C(data_i[4 ])  );
PDIDGZ    ipad_dat05( .PAD(data[5 ]), .C(data_i[5 ])  );
PDIDGZ    ipad_dat06( .PAD(data[6 ]), .C(data_i[6 ])  );
PDIDGZ    ipad_dat07( .PAD(data[7 ]), .C(data_i[7 ])  );
PDIDGZ    ipad_dat08( .PAD(data[8 ]), .C(data_i[8 ])  );
PDIDGZ    ipad_dat09( .PAD(data[9 ]), .C(data_i[9 ])  );
PDIDGZ    ipad_dat10( .PAD(data[10]), .C(data_i[10])  );
PDIDGZ    ipad_dat11( .PAD(data[11]), .C(data_i[11])  );
PDIDGZ    ipad_dat12( .PAD(data[12]), .C(data_i[12])  );
PDIDGZ    ipad_dat13( .PAD(data[13]), .C(data_i[13])  );
PDIDGZ    ipad_dat14( .PAD(data[14]), .C(data_i[14])  );
PDIDGZ    ipad_dat15( .PAD(data[15]), .C(data_i[15])  );
PDIDGZ    ipad_dat16( .PAD(data[16]), .C(data_i[16])  );
PDIDGZ    ipad_dat17( .PAD(data[17]), .C(data_i[17])  );
PDIDGZ    ipad_dat18( .PAD(data[18]), .C(data_i[18])  );
PDIDGZ    ipad_dat19( .PAD(data[19]), .C(data_i[19])  );
PDIDGZ    ipad_dat20( .PAD(data[20]), .C(data_i[20])  );
PDIDGZ    ipad_dat21( .PAD(data[21]), .C(data_i[21])  );
PDIDGZ    ipad_dat22( .PAD(data[22]), .C(data_i[22])  );
PDIDGZ    ipad_dat23( .PAD(data[23]), .C(data_i[23])  );
PDIDGZ    ipad_dat24( .PAD(data[24]), .C(data_i[24])  );
PDIDGZ    ipad_dat25( .PAD(data[25]), .C(data_i[25])  );
PDIDGZ    ipad_dat26( .PAD(data[26]), .C(data_i[26])  );
PDIDGZ    ipad_dat27( .PAD(data[27]), .C(data_i[27])  );
PDIDGZ    ipad_dat28( .PAD(data[28]), .C(data_i[28])  );
PDIDGZ    ipad_dat29( .PAD(data[29]), .C(data_i[29])  );
PDIDGZ    ipad_dat30( .PAD(data[30]), .C(data_i[30])  );
PDIDGZ    ipad_dat31( .PAD(data[31]), .C(data_i[31])  );


PDO12CDG  opad_busy( .PAD(busy)       ,.I(busy_i)   );
PDO12CDG  opad_outv( .PAD(out_valid)    ,.I(out_valid_i)    );
PDO12CDG  opad_done( .PAD(finish)     ,.I(finish_i)   );
PDO12CDG  opad_cw00( .PAD(codeword[ 0 ]) ,.I(codeword_i[ 0 ]) );
PDO12CDG  opad_cw01( .PAD(codeword[ 1 ]) ,.I(codeword_i[ 1 ]) );
PDO12CDG  opad_cw02( .PAD(codeword[ 2 ]) ,.I(codeword_i[ 2 ]) );
PDO12CDG  opad_cw03( .PAD(codeword[ 3 ]) ,.I(codeword_i[ 3 ]) );
PDO12CDG  opad_cw04( .PAD(codeword[ 4 ]) ,.I(codeword_i[ 4 ]) );
PDO12CDG  opad_cw05( .PAD(codeword[ 5 ]) ,.I(codeword_i[ 5 ]) );
PDO12CDG  opad_cw06( .PAD(codeword[ 6 ]) ,.I(codeword_i[ 6 ]) );
PDO12CDG  opad_cw07( .PAD(codeword[ 7 ]) ,.I(codeword_i[ 7 ]) );
PDO12CDG  opad_cw08( .PAD(codeword[ 8 ]) ,.I(codeword_i[ 8 ]) );
PDO12CDG  opad_cw09( .PAD(codeword[ 9 ]) ,.I(codeword_i[ 9 ]) );
PDO12CDG  opad_cw10( .PAD(codeword[10]) ,.I(codeword_i[10]) );

PDO12CDG  opad_en00( .PAD(enc_num[ 0 ])  ,.I(enc_num_i[ 0 ]) );
PDO12CDG  opad_en01( .PAD(enc_num[ 1 ])  ,.I(enc_num_i[ 1 ]) );
PDO12CDG  opad_en02( .PAD(enc_num[ 2 ])  ,.I(enc_num_i[ 2 ]) );
PDO12CDG  opad_en03( .PAD(enc_num[ 3 ])  ,.I(enc_num_i[ 3 ]) );
PDO12CDG  opad_en04( .PAD(enc_num[ 4 ])  ,.I(enc_num_i[ 4 ]) );
PDO12CDG  opad_en05( .PAD(enc_num[ 5 ])  ,.I(enc_num_i[ 5 ]) );
PDO12CDG  opad_en06( .PAD(enc_num[ 6 ])  ,.I(enc_num_i[ 6 ]) );
PDO12CDG  opad_en07( .PAD(enc_num[ 7 ])  ,.I(enc_num_i[ 7 ]) );
PDO12CDG  opad_en08( .PAD(enc_num[ 8 ])  ,.I(enc_num_i[ 8 ]) );
PDO12CDG  opad_en09( .PAD(enc_num[ 9 ])  ,.I(enc_num_i[ 9 ]) );
PDO12CDG  opad_en10( .PAD(enc_num[10])  ,.I(enc_num_i[10]) );
PDO12CDG  opad_en11( .PAD(enc_num[11])  ,.I(enc_num_i[11]) );

endmodule
