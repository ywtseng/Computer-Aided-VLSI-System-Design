
module FAS_DW01_add_0 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2;
  wire   [31:2] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  CLKINVX1 U2 ( .A(A[0]), .Y(n2) );
  XNOR2X1 U3 ( .A(B[0]), .B(n2), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_1 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_;
  wire   n1;
  wire   [35:4] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  XOR3XL U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[2]), .B(A_2_), .Y(n1) );
  XOR2X1 U2 ( .A(B[2]), .B(A_2_), .Y(SUM[2]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
  BUFX2 U4 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module FAS_DW01_add_2 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_3 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_;
  wire   n1;
  wire   [35:4] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[2]), .B(A_2_), .Y(n1) );
  XOR2X1 U2 ( .A(B[2]), .B(A_2_), .Y(SUM[2]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
  BUFX2 U4 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module FAS_DW01_add_4 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_5 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_6 ( A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, 
        A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, 
        A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, 
        A_2_, A_1_, B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, 
        B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, 
        B_2_, B_1_, B_0_, SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, 
        SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, 
        SUM_0_ );
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_,
         B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_,
         B_0_;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_,
         SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_,
         SUM_2_, SUM_1_, SUM_0_;
  wire   n1;
  wire   [31:3] carry;

  ADDFXL U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFXL U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFXL U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFXL U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  ADDFXL U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFXL U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFXL U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  ADDFXL U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFXL U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFXL U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(n1), .CO(carry[3]), .S(SUM_2_) );
  XOR3X1 U1_31 ( .A(A_31_), .B(B_31_), .C(carry[31]), .Y(SUM_31_) );
  AND2X2 U1 ( .A(B_1_), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B_1_), .B(A_1_), .Y(SUM_1_) );
  BUFX2 U3 ( .A(B_0_), .Y(SUM_0_) );
endmodule


module FAS_DW01_add_7 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_addsub_2 ( A, B, ADD_SUB, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input ADD_SUB;
  wire   carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_,
         carry_2_, carry_1_;
  wire   [15:0] B_AS;

  XOR3X1 U1_15 ( .A(A[15]), .B(B_AS[15]), .C(carry_15_), .Y(SUM[15]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B_AS[1]), .CI(carry_1_), .CO(carry_2_), .S(SUM[1]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B_AS[14]), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B_AS[13]), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B_AS[12]), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B_AS[11]), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B_AS[10]), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B_AS[9]), .CI(carry_9_), .CO(carry_10_), .S(
        SUM[9]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B_AS[8]), .CI(carry_8_), .CO(carry_9_), .S(SUM[8]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B_AS[7]), .CI(carry_7_), .CO(carry_8_), .S(SUM[7]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B_AS[6]), .CI(carry_6_), .CO(carry_7_), .S(SUM[6]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B_AS[5]), .CI(carry_5_), .CO(carry_6_), .S(SUM[5]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B_AS[4]), .CI(carry_4_), .CO(carry_5_), .S(SUM[4]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B_AS[3]), .CI(carry_3_), .CO(carry_4_), .S(SUM[3]) );
  ADDFXL U1_2 ( .A(A[2]), .B(B_AS[2]), .CI(carry_2_), .CO(carry_3_), .S(SUM[2]) );
  ADDFXL U1_0 ( .A(A[0]), .B(B_AS[0]), .CI(ADD_SUB), .CO(carry_1_), .S(SUM[0])
         );
  XOR2X1 U1 ( .A(B[9]), .B(ADD_SUB), .Y(B_AS[9]) );
  XOR2X1 U2 ( .A(B[8]), .B(ADD_SUB), .Y(B_AS[8]) );
  XOR2X1 U3 ( .A(B[7]), .B(ADD_SUB), .Y(B_AS[7]) );
  XOR2X1 U4 ( .A(B[6]), .B(ADD_SUB), .Y(B_AS[6]) );
  XOR2X1 U5 ( .A(B[5]), .B(ADD_SUB), .Y(B_AS[5]) );
  XOR2X1 U6 ( .A(B[4]), .B(ADD_SUB), .Y(B_AS[4]) );
  XOR2X1 U7 ( .A(B[3]), .B(ADD_SUB), .Y(B_AS[3]) );
  XOR2X1 U8 ( .A(B[2]), .B(ADD_SUB), .Y(B_AS[2]) );
  XOR2X1 U9 ( .A(B[1]), .B(ADD_SUB), .Y(B_AS[1]) );
  XOR2X1 U10 ( .A(B[15]), .B(ADD_SUB), .Y(B_AS[15]) );
  XOR2X1 U11 ( .A(B[14]), .B(ADD_SUB), .Y(B_AS[14]) );
  XOR2X1 U12 ( .A(B[13]), .B(ADD_SUB), .Y(B_AS[13]) );
  XOR2X1 U13 ( .A(B[12]), .B(ADD_SUB), .Y(B_AS[12]) );
  XOR2X1 U14 ( .A(B[11]), .B(ADD_SUB), .Y(B_AS[11]) );
  XOR2X1 U15 ( .A(B[10]), .B(ADD_SUB), .Y(B_AS[10]) );
  XOR2X1 U16 ( .A(B[0]), .B(ADD_SUB), .Y(B_AS[0]) );
endmodule


module FAS_DW01_add_8 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_9 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_10 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_11 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_12 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_13 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_14 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_15 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_sub_0 ( A, B, DIFF );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  ADDFXL U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_31 ( .A(A[31]), .B(n2), .C(carry[31]), .Y(DIFF[31]) );
  CLKINVX1 U1 ( .A(B[0]), .Y(n33) );
  CLKINVX1 U2 ( .A(B[31]), .Y(n2) );
  XNOR2X1 U3 ( .A(n33), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U4 ( .A(A[0]), .Y(n1) );
  NAND2X1 U5 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U6 ( .A(B[1]), .Y(n32) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n31) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n30) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n29) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n28) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n27) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n26) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n25) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n24) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n23) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n22) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n21) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n20) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n19) );
  CLKINVX1 U20 ( .A(B[15]), .Y(n18) );
  CLKINVX1 U21 ( .A(B[16]), .Y(n17) );
  CLKINVX1 U22 ( .A(B[17]), .Y(n16) );
  CLKINVX1 U23 ( .A(B[18]), .Y(n15) );
  CLKINVX1 U24 ( .A(B[19]), .Y(n14) );
  CLKINVX1 U25 ( .A(B[20]), .Y(n13) );
  CLKINVX1 U26 ( .A(B[21]), .Y(n12) );
  CLKINVX1 U27 ( .A(B[22]), .Y(n11) );
  CLKINVX1 U28 ( .A(B[23]), .Y(n10) );
  CLKINVX1 U29 ( .A(B[24]), .Y(n9) );
  CLKINVX1 U30 ( .A(B[25]), .Y(n8) );
  CLKINVX1 U31 ( .A(B[26]), .Y(n7) );
  CLKINVX1 U32 ( .A(B[27]), .Y(n6) );
  CLKINVX1 U33 ( .A(B[28]), .Y(n5) );
  CLKINVX1 U34 ( .A(B[29]), .Y(n4) );
  CLKINVX1 U35 ( .A(B[30]), .Y(n3) );
endmodule


module FAS_DW01_sub_1 ( A, B, DIFF );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  XOR3X1 U2_31 ( .A(A[31]), .B(n2), .C(carry[31]), .Y(DIFF[31]) );
  ADDFXL U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  CLKINVX1 U1 ( .A(B[0]), .Y(n33) );
  XNOR2X1 U2 ( .A(n33), .B(A[0]), .Y(DIFF[0]) );
  NAND2X1 U3 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n32) );
  CLKINVX1 U5 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U6 ( .A(B[2]), .Y(n31) );
  CLKINVX1 U7 ( .A(B[3]), .Y(n30) );
  CLKINVX1 U8 ( .A(B[4]), .Y(n29) );
  CLKINVX1 U9 ( .A(B[5]), .Y(n28) );
  CLKINVX1 U10 ( .A(B[6]), .Y(n27) );
  CLKINVX1 U11 ( .A(B[7]), .Y(n26) );
  CLKINVX1 U12 ( .A(B[8]), .Y(n25) );
  CLKINVX1 U13 ( .A(B[9]), .Y(n24) );
  CLKINVX1 U14 ( .A(B[10]), .Y(n23) );
  CLKINVX1 U15 ( .A(B[11]), .Y(n22) );
  CLKINVX1 U16 ( .A(B[12]), .Y(n21) );
  CLKINVX1 U17 ( .A(B[13]), .Y(n20) );
  CLKINVX1 U18 ( .A(B[14]), .Y(n19) );
  CLKINVX1 U19 ( .A(B[15]), .Y(n18) );
  CLKINVX1 U20 ( .A(B[16]), .Y(n17) );
  CLKINVX1 U21 ( .A(B[17]), .Y(n16) );
  CLKINVX1 U22 ( .A(B[18]), .Y(n15) );
  CLKINVX1 U23 ( .A(B[19]), .Y(n14) );
  CLKINVX1 U24 ( .A(B[20]), .Y(n13) );
  CLKINVX1 U25 ( .A(B[21]), .Y(n12) );
  CLKINVX1 U26 ( .A(B[22]), .Y(n11) );
  CLKINVX1 U27 ( .A(B[23]), .Y(n10) );
  CLKINVX1 U28 ( .A(B[24]), .Y(n9) );
  CLKINVX1 U29 ( .A(B[25]), .Y(n8) );
  CLKINVX1 U30 ( .A(B[26]), .Y(n7) );
  CLKINVX1 U31 ( .A(B[27]), .Y(n6) );
  CLKINVX1 U32 ( .A(B[28]), .Y(n5) );
  CLKINVX1 U33 ( .A(B[29]), .Y(n4) );
  CLKINVX1 U34 ( .A(B[30]), .Y(n3) );
  CLKINVX1 U35 ( .A(B[31]), .Y(n2) );
endmodule


module FAS_DW01_addsub_3 ( A, B, SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, 
        SUM_26_, SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, 
        SUM_18_, SUM_17_, SUM_16_ );
  input [31:0] A;
  input [31:0] B;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;
  wire   [31:16] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM_31_) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  OAI2BB1X1 U1 ( .A0N(n1), .A1N(A[15]), .B0(n2), .Y(carry[16]) );
  OAI21XL U2 ( .A0(A[15]), .A1(n1), .B0(B[15]), .Y(n2) );
  OAI2BB1X1 U3 ( .A0N(n3), .A1N(A[14]), .B0(n4), .Y(n1) );
  OAI21XL U4 ( .A0(A[14]), .A1(n3), .B0(B[14]), .Y(n4) );
  OAI2BB1X1 U5 ( .A0N(n5), .A1N(A[13]), .B0(n6), .Y(n3) );
  OAI21XL U6 ( .A0(A[13]), .A1(n5), .B0(B[13]), .Y(n6) );
  OAI2BB1X1 U7 ( .A0N(n7), .A1N(A[12]), .B0(n8), .Y(n5) );
  OAI21XL U8 ( .A0(A[12]), .A1(n7), .B0(B[12]), .Y(n8) );
  OAI2BB1X1 U9 ( .A0N(n9), .A1N(A[11]), .B0(n10), .Y(n7) );
  OAI21XL U10 ( .A0(A[11]), .A1(n9), .B0(B[11]), .Y(n10) );
  OAI2BB1X1 U11 ( .A0N(n11), .A1N(A[10]), .B0(n12), .Y(n9) );
  OAI21XL U12 ( .A0(A[10]), .A1(n11), .B0(B[10]), .Y(n12) );
  OAI2BB1X1 U13 ( .A0N(n13), .A1N(A[9]), .B0(n14), .Y(n11) );
  OAI21XL U14 ( .A0(A[9]), .A1(n13), .B0(B[9]), .Y(n14) );
  OAI2BB1X1 U15 ( .A0N(n15), .A1N(A[8]), .B0(n16), .Y(n13) );
  OAI21XL U16 ( .A0(A[8]), .A1(n15), .B0(B[8]), .Y(n16) );
  OAI2BB1X1 U17 ( .A0N(n17), .A1N(A[7]), .B0(n18), .Y(n15) );
  OAI21XL U18 ( .A0(A[7]), .A1(n17), .B0(B[7]), .Y(n18) );
  OAI2BB1X1 U19 ( .A0N(n19), .A1N(A[6]), .B0(n20), .Y(n17) );
  OAI21XL U20 ( .A0(A[6]), .A1(n19), .B0(B[6]), .Y(n20) );
  OAI2BB1X1 U21 ( .A0N(n21), .A1N(A[5]), .B0(n22), .Y(n19) );
  OAI21XL U22 ( .A0(A[5]), .A1(n21), .B0(B[5]), .Y(n22) );
  OAI2BB1X1 U23 ( .A0N(n23), .A1N(A[4]), .B0(n24), .Y(n21) );
  OAI21XL U24 ( .A0(A[4]), .A1(n23), .B0(B[4]), .Y(n24) );
  OAI2BB1X1 U25 ( .A0N(n25), .A1N(A[3]), .B0(n26), .Y(n23) );
  OAI21XL U26 ( .A0(A[3]), .A1(n25), .B0(B[3]), .Y(n26) );
  OAI2BB1X1 U27 ( .A0N(n27), .A1N(A[2]), .B0(n28), .Y(n25) );
  OAI21XL U28 ( .A0(A[2]), .A1(n27), .B0(B[2]), .Y(n28) );
  OAI2BB1X1 U29 ( .A0N(A[1]), .A1N(B[1]), .B0(n29), .Y(n27) );
  OAI211X1 U30 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n29) );
endmodule


module FAS_DW01_add_16 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_17 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_18 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_;
  wire   n1;
  wire   [35:4] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[2]), .B(A_2_), .Y(n1) );
  XOR2X1 U2 ( .A(B[2]), .B(A_2_), .Y(SUM[2]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
  BUFX2 U4 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module FAS_DW01_add_19 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_20 ( A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, 
        A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, 
        A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, 
        A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, B_35_, B_34_, B_33_, 
        B_32_, B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, 
        B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, 
        B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, 
        B_1_, SUM_35_, SUM_34_, SUM_33_, SUM_32_, SUM_31_, SUM_30_, SUM_29_, 
        SUM_28_, SUM_27_, SUM_26_, SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, 
        SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, 
        SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, 
        SUM_4_, SUM_3_, SUM_2_, SUM_1_ );
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_, B_35_, B_34_, B_33_, B_32_, B_31_,
         B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_, B_21_,
         B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_,
         B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_;
  output SUM_35_, SUM_34_, SUM_33_, SUM_32_, SUM_31_, SUM_30_, SUM_29_,
         SUM_28_, SUM_27_, SUM_26_, SUM_25_, SUM_24_, SUM_23_, SUM_22_,
         SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B_34_), .CI(carry[34]), .CO(carry[35]), .S(
        SUM_34_) );
  ADDFXL U1_33 ( .A(A_33_), .B(B_33_), .CI(carry[33]), .CO(carry[34]), .S(
        SUM_33_) );
  ADDFXL U1_32 ( .A(A_32_), .B(B_32_), .CI(carry[32]), .CO(carry[33]), .S(
        SUM_32_) );
  ADDFXL U1_31 ( .A(A_31_), .B(B_31_), .CI(carry[31]), .CO(carry[32]), .S(
        SUM_31_) );
  ADDFXL U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFXL U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFXL U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFXL U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  ADDFXL U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFXL U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFXL U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  ADDFXL U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFXL U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFXL U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(n1), .CO(carry[3]), .S(SUM_2_) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B_35_), .C(carry[35]), .Y(SUM_35_) );
  AND2X2 U1 ( .A(B_1_), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B_1_), .B(A_1_), .Y(SUM_1_) );
endmodule


module FAS_DW01_add_21 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_;
  wire   n1;
  wire   [35:4] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[2]), .B(A_2_), .Y(n1) );
  XOR2X1 U2 ( .A(B[2]), .B(A_2_), .Y(SUM[2]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
  BUFX2 U4 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module FAS_DW01_add_22 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_;
  wire   n1;
  wire   [35:4] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[2]), .B(A_2_), .Y(n1) );
  XOR2X1 U2 ( .A(B[2]), .B(A_2_), .Y(SUM[2]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
  BUFX2 U4 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module FAS_DW01_add_23 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_;
  wire   n1;
  wire   [35:4] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[2]), .B(A_2_), .Y(n1) );
  XOR2X1 U2 ( .A(B[2]), .B(A_2_), .Y(SUM[2]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
  BUFX2 U4 ( .A(B[1]), .Y(SUM[1]) );
endmodule


module FAS_DW01_add_24 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_25 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_26 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_27 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_sub_2 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n4), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n5), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n6), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n7), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n8), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n9), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n10), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n11), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n13), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n14), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n16), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n17), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n3), .C(carry[15]), .Y(DIFF[15]) );
  CLKINVX1 U1 ( .A(B[15]), .Y(n3) );
  CLKINVX1 U2 ( .A(B[0]), .Y(n2) );
  XNOR2X1 U3 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U4 ( .A(A[0]), .Y(n1) );
  NAND2X1 U5 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U6 ( .A(B[1]), .Y(n17) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n16) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n15) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n14) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n13) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n12) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n11) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n10) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n9) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n8) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n7) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n6) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n5) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n4) );
endmodule


module FAS_DW01_add_28 ( A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, 
        A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, 
        A_3_, A_2_, A_1_, B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, 
        B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        B_3_, B_2_, B_1_, SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, 
        SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_ );
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_,
         B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [31:16] carry;

  ADDFXL U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFXL U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFXL U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFXL U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  ADDFXL U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFXL U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFXL U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  ADDFXL U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFXL U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFXL U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  XOR3X1 U1_31 ( .A(A_31_), .B(B_31_), .C(carry[31]), .Y(SUM_31_) );
  AND2X2 U1 ( .A(A_1_), .B(B_1_), .Y(n1) );
  OAI2BB1X1 U2 ( .A0N(n2), .A1N(A_15_), .B0(n3), .Y(carry[16]) );
  OAI21XL U3 ( .A0(A_15_), .A1(n2), .B0(B_15_), .Y(n3) );
  OAI2BB1X1 U4 ( .A0N(n4), .A1N(A_14_), .B0(n5), .Y(n2) );
  OAI21XL U5 ( .A0(A_14_), .A1(n4), .B0(B_14_), .Y(n5) );
  OAI2BB1X1 U6 ( .A0N(n6), .A1N(A_13_), .B0(n7), .Y(n4) );
  OAI21XL U7 ( .A0(A_13_), .A1(n6), .B0(B_13_), .Y(n7) );
  OAI2BB1X1 U8 ( .A0N(n8), .A1N(A_12_), .B0(n9), .Y(n6) );
  OAI21XL U9 ( .A0(A_12_), .A1(n8), .B0(B_12_), .Y(n9) );
  OAI2BB1X1 U10 ( .A0N(n10), .A1N(A_11_), .B0(n11), .Y(n8) );
  OAI21XL U11 ( .A0(A_11_), .A1(n10), .B0(B_11_), .Y(n11) );
  OAI2BB1X1 U12 ( .A0N(n12), .A1N(A_10_), .B0(n13), .Y(n10) );
  OAI21XL U13 ( .A0(A_10_), .A1(n12), .B0(B_10_), .Y(n13) );
  OAI2BB1X1 U14 ( .A0N(n14), .A1N(A_9_), .B0(n15), .Y(n12) );
  OAI21XL U15 ( .A0(A_9_), .A1(n14), .B0(B_9_), .Y(n15) );
  OAI2BB1X1 U16 ( .A0N(n16), .A1N(A_8_), .B0(n17), .Y(n14) );
  OAI21XL U17 ( .A0(A_8_), .A1(n16), .B0(B_8_), .Y(n17) );
  OAI2BB1X1 U18 ( .A0N(n18), .A1N(A_7_), .B0(n19), .Y(n16) );
  OAI21XL U19 ( .A0(A_7_), .A1(n18), .B0(B_7_), .Y(n19) );
  OAI2BB1X1 U20 ( .A0N(n20), .A1N(A_6_), .B0(n21), .Y(n18) );
  OAI21XL U21 ( .A0(A_6_), .A1(n20), .B0(B_6_), .Y(n21) );
  OAI2BB1X1 U22 ( .A0N(n22), .A1N(A_5_), .B0(n23), .Y(n20) );
  OAI21XL U23 ( .A0(A_5_), .A1(n22), .B0(B_5_), .Y(n23) );
  OAI2BB1X1 U24 ( .A0N(n24), .A1N(A_4_), .B0(n25), .Y(n22) );
  OAI21XL U25 ( .A0(A_4_), .A1(n24), .B0(B_4_), .Y(n25) );
  OAI2BB1X1 U26 ( .A0N(n26), .A1N(A_3_), .B0(n27), .Y(n24) );
  OAI21XL U27 ( .A0(A_3_), .A1(n26), .B0(B_3_), .Y(n27) );
  OAI2BB1X1 U28 ( .A0N(n1), .A1N(A_2_), .B0(n28), .Y(n26) );
  OAI21XL U29 ( .A0(A_2_), .A1(n1), .B0(B_2_), .Y(n28) );
endmodule


module FAS_DW01_add_29 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_30 ( A, B, SUM );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  wire   n1;
  wire   [35:2] carry;

  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_35 ( .A(A[35]), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_sub_3 ( A, B, DIFF );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  ADDFXL U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_31 ( .A(A[31]), .B(n2), .C(carry[31]), .Y(DIFF[31]) );
  CLKINVX1 U1 ( .A(B[0]), .Y(n33) );
  CLKINVX1 U2 ( .A(B[31]), .Y(n2) );
  XNOR2X1 U3 ( .A(n33), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U4 ( .A(A[0]), .Y(n1) );
  NAND2X1 U5 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U6 ( .A(B[1]), .Y(n32) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n31) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n30) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n29) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n28) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n27) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n26) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n25) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n24) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n23) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n22) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n21) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n20) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n19) );
  CLKINVX1 U20 ( .A(B[15]), .Y(n18) );
  CLKINVX1 U21 ( .A(B[16]), .Y(n17) );
  CLKINVX1 U22 ( .A(B[17]), .Y(n16) );
  CLKINVX1 U23 ( .A(B[18]), .Y(n15) );
  CLKINVX1 U24 ( .A(B[19]), .Y(n14) );
  CLKINVX1 U25 ( .A(B[20]), .Y(n13) );
  CLKINVX1 U26 ( .A(B[21]), .Y(n12) );
  CLKINVX1 U27 ( .A(B[22]), .Y(n11) );
  CLKINVX1 U28 ( .A(B[23]), .Y(n10) );
  CLKINVX1 U29 ( .A(B[24]), .Y(n9) );
  CLKINVX1 U30 ( .A(B[25]), .Y(n8) );
  CLKINVX1 U31 ( .A(B[26]), .Y(n7) );
  CLKINVX1 U32 ( .A(B[27]), .Y(n6) );
  CLKINVX1 U33 ( .A(B[28]), .Y(n5) );
  CLKINVX1 U34 ( .A(B[29]), .Y(n4) );
  CLKINVX1 U35 ( .A(B[30]), .Y(n3) );
endmodule


module FAS_DW01_sub_4 ( A, B, DIFF );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  ADDFXL U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_31 ( .A(A[31]), .B(n2), .C(carry[31]), .Y(DIFF[31]) );
  CLKINVX1 U1 ( .A(B[0]), .Y(n33) );
  CLKINVX1 U2 ( .A(B[31]), .Y(n2) );
  XNOR2X1 U3 ( .A(n33), .B(A[0]), .Y(DIFF[0]) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n32) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n31) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n30) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n29) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n28) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n27) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n26) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n25) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n24) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n23) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n22) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n21) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n20) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n19) );
  CLKINVX1 U20 ( .A(B[15]), .Y(n18) );
  CLKINVX1 U21 ( .A(B[16]), .Y(n17) );
  CLKINVX1 U22 ( .A(B[17]), .Y(n16) );
  CLKINVX1 U23 ( .A(B[18]), .Y(n15) );
  CLKINVX1 U24 ( .A(B[19]), .Y(n14) );
  CLKINVX1 U25 ( .A(B[20]), .Y(n13) );
  CLKINVX1 U26 ( .A(B[21]), .Y(n12) );
  CLKINVX1 U27 ( .A(B[22]), .Y(n11) );
  CLKINVX1 U28 ( .A(B[23]), .Y(n10) );
  CLKINVX1 U29 ( .A(B[24]), .Y(n9) );
  CLKINVX1 U30 ( .A(B[25]), .Y(n8) );
  CLKINVX1 U31 ( .A(B[26]), .Y(n7) );
  CLKINVX1 U32 ( .A(B[27]), .Y(n6) );
  CLKINVX1 U33 ( .A(B[28]), .Y(n5) );
  CLKINVX1 U34 ( .A(B[29]), .Y(n4) );
  CLKINVX1 U35 ( .A(B[30]), .Y(n3) );
endmodule


module FAS_DW01_add_31 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1;
  wire   [31:2] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_32 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1;
  wire   [31:2] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_33 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1;
  wire   [31:2] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_sub_5 ( A, B, DIFF );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [31:1] carry;

  XOR3X1 U2_31 ( .A(A[31]), .B(n2), .C(carry[31]), .Y(DIFF[31]) );
  ADDFXL U2_3 ( .A(A[3]), .B(n30), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n32), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n27), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n28), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n29), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n31), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_30 ( .A(A[30]), .B(n3), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n4), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n5), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n6), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n7), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n8), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n9), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n10), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n11), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n18), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n19), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n20), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n22), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n23), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n24), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n25), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n26), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_21 ( .A(A[21]), .B(n12), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n13), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n14), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n15), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  CLKINVX1 U1 ( .A(B[16]), .Y(n17) );
  CLKINVX1 U2 ( .A(B[17]), .Y(n16) );
  CLKINVX1 U3 ( .A(B[18]), .Y(n15) );
  CLKINVX1 U4 ( .A(B[19]), .Y(n14) );
  CLKINVX1 U5 ( .A(B[20]), .Y(n13) );
  CLKINVX1 U6 ( .A(B[21]), .Y(n12) );
  CLKINVX1 U7 ( .A(B[7]), .Y(n26) );
  CLKINVX1 U8 ( .A(B[8]), .Y(n25) );
  CLKINVX1 U9 ( .A(B[9]), .Y(n24) );
  CLKINVX1 U10 ( .A(B[10]), .Y(n23) );
  CLKINVX1 U11 ( .A(B[11]), .Y(n22) );
  CLKINVX1 U12 ( .A(B[12]), .Y(n21) );
  CLKINVX1 U13 ( .A(B[13]), .Y(n20) );
  CLKINVX1 U14 ( .A(B[14]), .Y(n19) );
  CLKINVX1 U15 ( .A(B[15]), .Y(n18) );
  CLKINVX1 U16 ( .A(B[22]), .Y(n11) );
  CLKINVX1 U17 ( .A(B[23]), .Y(n10) );
  CLKINVX1 U18 ( .A(B[24]), .Y(n9) );
  CLKINVX1 U19 ( .A(B[25]), .Y(n8) );
  CLKINVX1 U20 ( .A(B[26]), .Y(n7) );
  CLKINVX1 U21 ( .A(B[27]), .Y(n6) );
  CLKINVX1 U22 ( .A(B[28]), .Y(n5) );
  CLKINVX1 U23 ( .A(B[29]), .Y(n4) );
  CLKINVX1 U24 ( .A(B[30]), .Y(n3) );
  XNOR2X1 U25 ( .A(n33), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U26 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U27 ( .A(B[2]), .Y(n31) );
  CLKINVX1 U28 ( .A(B[4]), .Y(n29) );
  CLKINVX1 U29 ( .A(B[5]), .Y(n28) );
  CLKINVX1 U30 ( .A(B[6]), .Y(n27) );
  CLKINVX1 U31 ( .A(B[0]), .Y(n33) );
  NAND2X1 U32 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U33 ( .A(B[1]), .Y(n32) );
  CLKINVX1 U34 ( .A(B[3]), .Y(n30) );
  CLKINVX1 U35 ( .A(B[31]), .Y(n2) );
endmodule


module FAS_DW01_sub_6 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  CLKINVX1 U1 ( .A(B[0]), .Y(n17) );
  XNOR2X1 U2 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  NAND2X1 U3 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n16) );
  CLKINVX1 U5 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U6 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U7 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U8 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U9 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U10 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U11 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U12 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U13 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U14 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U15 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U16 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U17 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[14]), .Y(n3) );
  CLKINVX1 U19 ( .A(B[15]), .Y(n2) );
endmodule


module FAS_DW01_add_34 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_35 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_36 ( B, SUM, A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, 
        A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, 
        A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [35:0] B;
  output [35:0] SUM;
  input A_35_, A_34_, A_33_, A_32_, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_,
         A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_,
         A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_,
         A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n1;
  wire   [35:3] carry;

  ADDFXL U1_34 ( .A(A_34_), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_33 ( .A(A_33_), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_32 ( .A(A_32_), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_31 ( .A(A_31_), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_35 ( .A(A_35_), .B(B[35]), .C(carry[35]), .Y(SUM[35]) );
  AND2X2 U1 ( .A(B[1]), .B(A_1_), .Y(n1) );
  XOR2X1 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  BUFX2 U3 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module FAS_DW01_add_37 ( SUM, A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, 
        A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, 
        A_3_, A_2_, A_0_, B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, 
        B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, 
        B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, 
        B_3_, B_2_, B_0_ );
  output [31:0] SUM;
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_0_,
         B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_0_;
  wire   n1;
  wire   [31:4] carry;

  XOR3X1 U1_31 ( .A(A_31_), .B(B_31_), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  AND2X2 U1 ( .A(B_2_), .B(A_2_), .Y(n1) );
  XOR2X1 U2 ( .A(B_2_), .B(A_2_), .Y(SUM[2]) );
  XOR2X1 U3 ( .A(B_0_), .B(A_0_), .Y(SUM[0]) );
  AND2X2 U4 ( .A(B_0_), .B(A_0_), .Y(SUM[1]) );
endmodule


module FAS_DW_mult_tc_22 ( a, product_31_, product_30_, product_29_, 
        product_28_, product_27_, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_, product_14_, 
        product_13_, product_12_, product_11_, product_10_, product_9_, 
        product_8_, product_7_, product_6_, product_5_, product_4_, product_3_, 
        product_2_, product_0_ );
  input [15:0] a;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_0_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328;

  CLKINVX1 U1 ( .A(n1), .Y(product_31_) );
  ADDFXL U2 ( .A(n179), .B(a[15]), .CI(n2), .CO(n1), .S(product_30_) );
  ADDFXL U3 ( .A(n30), .B(n180), .CI(n3), .CO(n2), .S(product_29_) );
  ADDFXL U4 ( .A(n32), .B(n31), .CI(n4), .CO(n3), .S(product_28_) );
  ADDFXL U5 ( .A(n35), .B(n33), .CI(n5), .CO(n4), .S(product_27_) );
  ADDFXL U6 ( .A(n38), .B(n36), .CI(n6), .CO(n5), .S(product_26_) );
  ADDFXL U7 ( .A(n41), .B(n39), .CI(n7), .CO(n6), .S(product_25_) );
  ADDFXL U8 ( .A(n42), .B(n46), .CI(n8), .CO(n7), .S(product_24_) );
  ADDFXL U9 ( .A(n51), .B(n47), .CI(n9), .CO(n8), .S(product_23_) );
  ADDFXL U10 ( .A(n52), .B(n57), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U11 ( .A(n58), .B(n63), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U12 ( .A(n64), .B(n71), .CI(n12), .CO(n11), .S(product_20_) );
  ADDFXL U13 ( .A(n79), .B(n72), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFXL U14 ( .A(n80), .B(n88), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFXL U15 ( .A(n89), .B(n97), .CI(n15), .CO(n14), .S(product_17_) );
  ADDFXL U16 ( .A(n98), .B(n108), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFXL U17 ( .A(n109), .B(n118), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFXL U18 ( .A(n119), .B(n128), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFXL U19 ( .A(n129), .B(n136), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFXL U20 ( .A(n137), .B(n144), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFXL U21 ( .A(n145), .B(n151), .CI(n21), .CO(n20), .S(product_11_) );
  ADDFXL U22 ( .A(n152), .B(n158), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFXL U23 ( .A(n159), .B(n163), .CI(n23), .CO(n22), .S(product_9_) );
  ADDFXL U24 ( .A(n164), .B(n167), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFXL U25 ( .A(n168), .B(n171), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFXL U26 ( .A(n172), .B(n174), .CI(n26), .CO(n25), .S(product_6_) );
  ADDFXL U27 ( .A(n176), .B(n177), .CI(n27), .CO(n26), .S(product_5_) );
  ADDFXL U28 ( .A(n178), .B(n295), .CI(n28), .CO(n27), .S(product_4_) );
  ADDHXL U29 ( .A(n297), .B(n29), .CO(n28), .S(product_3_) );
  ADDHXL U30 ( .A(a[1]), .B(n298), .CO(n29), .S(product_2_) );
  ADDFXL U31 ( .A(n194), .B(a[14]), .CI(n181), .CO(n30), .S(n31) );
  ADDFXL U32 ( .A(n182), .B(n195), .CI(n34), .CO(n32), .S(n33) );
  CMPR42X1 U33 ( .A(a[13]), .B(n196), .C(n208), .D(n183), .ICI(n37), .S(n36), 
        .ICO(n34), .CO(n35) );
  CMPR42X1 U34 ( .A(n209), .B(n197), .C(n184), .D(n43), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U35 ( .A(n221), .B(n210), .C(n44), .D(n48), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFXL U36 ( .A(n198), .B(a[12]), .CI(n185), .CO(n43), .S(n44) );
  CMPR42X1 U37 ( .A(n199), .B(n53), .C(n49), .D(n54), .ICI(n50), .S(n47), 
        .ICO(n45), .CO(n46) );
  ADDFXL U38 ( .A(n211), .B(n222), .CI(n186), .CO(n48), .S(n49) );
  CMPR42X1 U39 ( .A(n223), .B(n212), .C(n60), .D(n55), .ICI(n56), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U40 ( .A(a[11]), .B(n200), .C(n233), .D(n187), .ICI(n59), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U41 ( .A(n201), .B(n68), .C(n66), .D(n61), .ICI(n62), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U42 ( .A(n213), .B(n234), .C(n224), .D(n188), .ICI(n65), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U43 ( .A(n69), .B(n76), .C(n74), .D(n67), .ICI(n70), .S(n64), .ICO(
        n62), .CO(n63) );
  CMPR42X1 U44 ( .A(n225), .B(n244), .C(n235), .D(n214), .ICI(n73), .S(n67), 
        .ICO(n65), .CO(n66) );
  ADDFXL U45 ( .A(n202), .B(a[10]), .CI(n189), .CO(n68), .S(n69) );
  CMPR42X1 U46 ( .A(n77), .B(n85), .C(n82), .D(n75), .ICI(n78), .S(n72), .ICO(
        n70), .CO(n71) );
  CMPR42X1 U47 ( .A(n236), .B(n215), .C(n226), .D(n84), .ICI(n81), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFXL U48 ( .A(n203), .B(n245), .CI(n190), .CO(n76), .S(n77) );
  CMPR42X1 U49 ( .A(n94), .B(n91), .C(n86), .D(n83), .ICI(n87), .S(n80), .ICO(
        n78), .CO(n79) );
  CMPR42X1 U50 ( .A(n227), .B(n246), .C(n237), .D(n216), .ICI(n90), .S(n83), 
        .ICO(n81), .CO(n82) );
  CMPR42X1 U51 ( .A(a[9]), .B(n204), .C(n254), .D(n191), .ICI(n93), .S(n86), 
        .ICO(n84), .CO(n85) );
  CMPR42X1 U52 ( .A(n103), .B(n100), .C(n92), .D(n95), .ICI(n96), .S(n89), 
        .ICO(n87), .CO(n88) );
  CMPR42X1 U53 ( .A(n228), .B(n247), .C(n238), .D(n217), .ICI(n99), .S(n92), 
        .ICO(n90), .CO(n91) );
  CMPR42X1 U54 ( .A(n255), .B(n205), .C(n192), .D(n105), .ICI(n102), .S(n95), 
        .ICO(n93), .CO(n94) );
  CMPR42X1 U55 ( .A(n113), .B(n111), .C(n101), .D(n104), .ICI(n107), .S(n98), 
        .ICO(n96), .CO(n97) );
  CMPR42X1 U56 ( .A(n248), .B(n218), .C(n229), .D(n239), .ICI(n115), .S(n101), 
        .ICO(n99), .CO(n100) );
  CMPR42X1 U57 ( .A(n256), .B(n206), .C(n193), .D(n106), .ICI(n110), .S(n104), 
        .ICO(n102), .CO(n103) );
  XNOR2X1 U58 ( .A(n263), .B(a[8]), .Y(n106) );
  OR2X1 U59 ( .A(n263), .B(a[8]), .Y(n105) );
  CMPR42X1 U60 ( .A(n123), .B(n114), .C(n121), .D(n112), .ICI(n117), .S(n109), 
        .ICO(n107), .CO(n108) );
  CMPR42X1 U61 ( .A(n257), .B(n230), .C(n249), .D(n116), .ICI(n120), .S(n112), 
        .ICO(n110), .CO(n111) );
  ADDFXL U62 ( .A(n264), .B(n240), .CI(n125), .CO(n113), .S(n114) );
  ADDHXL U63 ( .A(n219), .B(n207), .CO(n115), .S(n116) );
  CMPR42X1 U64 ( .A(n250), .B(n124), .C(n131), .D(n122), .ICI(n127), .S(n119), 
        .ICO(n117), .CO(n118) );
  CMPR42X1 U65 ( .A(n265), .B(n241), .C(n258), .D(n133), .ICI(n130), .S(n122), 
        .ICO(n120), .CO(n121) );
  ADDFXL U66 ( .A(n231), .B(n271), .CI(n126), .CO(n123), .S(n124) );
  ADDHXL U67 ( .A(a[7]), .B(n220), .CO(n125), .S(n126) );
  CMPR42X1 U68 ( .A(n251), .B(n134), .C(n139), .D(n132), .ICI(n135), .S(n129), 
        .ICO(n127), .CO(n128) );
  CMPR42X1 U69 ( .A(n259), .B(n272), .C(n266), .D(n141), .ICI(n138), .S(n132), 
        .ICO(n130), .CO(n131) );
  ADDHXL U70 ( .A(n242), .B(n232), .CO(n133), .S(n134) );
  CMPR42X1 U71 ( .A(n267), .B(n260), .C(n146), .D(n143), .ICI(n140), .S(n137), 
        .ICO(n135), .CO(n136) );
  CMPR42X1 U72 ( .A(n278), .B(n252), .C(n273), .D(n148), .ICI(n142), .S(n140), 
        .ICO(n138), .CO(n139) );
  ADDHXL U73 ( .A(a[6]), .B(n243), .CO(n141), .S(n142) );
  CMPR42X1 U74 ( .A(n279), .B(n149), .C(n150), .D(n153), .ICI(n147), .S(n145), 
        .ICO(n143), .CO(n144) );
  ADDFXL U75 ( .A(n274), .B(n268), .CI(n155), .CO(n146), .S(n147) );
  ADDHXL U76 ( .A(n261), .B(n253), .CO(n148), .S(n149) );
  CMPR42X1 U77 ( .A(n280), .B(n275), .C(n160), .D(n157), .ICI(n154), .S(n152), 
        .ICO(n150), .CO(n151) );
  ADDFXL U78 ( .A(n269), .B(n284), .CI(n156), .CO(n153), .S(n154) );
  ADDHXL U79 ( .A(a[5]), .B(n262), .CO(n155), .S(n156) );
  CMPR42X1 U80 ( .A(n285), .B(n281), .C(n165), .D(n161), .ICI(n162), .S(n159), 
        .ICO(n157), .CO(n158) );
  ADDHXL U81 ( .A(n276), .B(n270), .CO(n160), .S(n161) );
  CMPR42X1 U82 ( .A(n289), .B(n282), .C(n286), .D(n169), .ICI(n166), .S(n164), 
        .ICO(n162), .CO(n163) );
  ADDHXL U83 ( .A(a[4]), .B(n277), .CO(n165), .S(n166) );
  ADDFXL U84 ( .A(n173), .B(n287), .CI(n170), .CO(n167), .S(n168) );
  ADDHXL U85 ( .A(n290), .B(n283), .CO(n169), .S(n170) );
  ADDFXL U86 ( .A(n291), .B(n293), .CI(n175), .CO(n171), .S(n172) );
  ADDHXL U87 ( .A(a[3]), .B(n288), .CO(n173), .S(n174) );
  ADDHXL U88 ( .A(n294), .B(n292), .CO(n175), .S(n176) );
  ADDHXL U89 ( .A(a[2]), .B(n296), .CO(n177), .S(n178) );
  OR2X1 U90 ( .A(n315), .B(n314), .Y(n179) );
  OR2X1 U91 ( .A(n316), .B(n314), .Y(n180) );
  OR2X1 U92 ( .A(n317), .B(n314), .Y(n181) );
  OR2X1 U93 ( .A(n318), .B(n314), .Y(n182) );
  OR2X1 U94 ( .A(n319), .B(n314), .Y(n183) );
  OR2X1 U95 ( .A(n320), .B(n314), .Y(n184) );
  OR2X1 U96 ( .A(n321), .B(n314), .Y(n185) );
  OR2X1 U97 ( .A(n322), .B(n314), .Y(n186) );
  OR2X1 U98 ( .A(n323), .B(n314), .Y(n187) );
  OR2X1 U99 ( .A(n324), .B(n314), .Y(n188) );
  OR2X1 U100 ( .A(n325), .B(n314), .Y(n189) );
  OR2X1 U101 ( .A(n326), .B(n314), .Y(n190) );
  OR2X1 U102 ( .A(n327), .B(n314), .Y(n191) );
  OR2X1 U103 ( .A(n328), .B(n314), .Y(n192) );
  OR2X1 U104 ( .A(n313), .B(n314), .Y(n193) );
  NOR2X1 U105 ( .A(n316), .B(n315), .Y(n194) );
  NOR2X1 U106 ( .A(n317), .B(n315), .Y(n195) );
  NOR2X1 U107 ( .A(n318), .B(n315), .Y(n196) );
  NOR2X1 U108 ( .A(n319), .B(n315), .Y(n197) );
  NOR2X1 U109 ( .A(n320), .B(n315), .Y(n198) );
  NOR2X1 U110 ( .A(n321), .B(n315), .Y(n199) );
  NOR2X1 U111 ( .A(n322), .B(n315), .Y(n200) );
  NOR2X1 U112 ( .A(n323), .B(n315), .Y(n201) );
  NOR2X1 U113 ( .A(n324), .B(n315), .Y(n202) );
  NOR2X1 U114 ( .A(n325), .B(n315), .Y(n203) );
  NOR2X1 U115 ( .A(n326), .B(n315), .Y(n204) );
  NOR2X1 U116 ( .A(n327), .B(n315), .Y(n205) );
  NOR2X1 U117 ( .A(n328), .B(n315), .Y(n206) );
  NOR2X1 U118 ( .A(n313), .B(n315), .Y(n207) );
  NOR2X1 U119 ( .A(n317), .B(n316), .Y(n208) );
  NOR2X1 U120 ( .A(n318), .B(n316), .Y(n209) );
  NOR2X1 U121 ( .A(n319), .B(n316), .Y(n210) );
  NOR2X1 U122 ( .A(n320), .B(n316), .Y(n211) );
  NOR2X1 U123 ( .A(n321), .B(n316), .Y(n212) );
  NOR2X1 U124 ( .A(n322), .B(n316), .Y(n213) );
  NOR2X1 U125 ( .A(n323), .B(n316), .Y(n214) );
  NOR2X1 U126 ( .A(n324), .B(n316), .Y(n215) );
  NOR2X1 U127 ( .A(n325), .B(n316), .Y(n216) );
  NOR2X1 U128 ( .A(n326), .B(n316), .Y(n217) );
  NOR2X1 U129 ( .A(n327), .B(n316), .Y(n218) );
  NOR2X1 U130 ( .A(n328), .B(n316), .Y(n219) );
  NOR2X1 U131 ( .A(n313), .B(n316), .Y(n220) );
  NOR2X1 U132 ( .A(n318), .B(n317), .Y(n221) );
  NOR2X1 U133 ( .A(n319), .B(n317), .Y(n222) );
  NOR2X1 U134 ( .A(n320), .B(n317), .Y(n223) );
  NOR2X1 U135 ( .A(n321), .B(n317), .Y(n224) );
  NOR2X1 U136 ( .A(n322), .B(n317), .Y(n225) );
  NOR2X1 U137 ( .A(n323), .B(n317), .Y(n226) );
  NOR2X1 U138 ( .A(n324), .B(n317), .Y(n227) );
  NOR2X1 U139 ( .A(n325), .B(n317), .Y(n228) );
  NOR2X1 U140 ( .A(n326), .B(n317), .Y(n229) );
  NOR2X1 U141 ( .A(n327), .B(n317), .Y(n230) );
  NOR2X1 U142 ( .A(n328), .B(n317), .Y(n231) );
  NOR2X1 U143 ( .A(n313), .B(n317), .Y(n232) );
  NOR2X1 U144 ( .A(n319), .B(n318), .Y(n233) );
  NOR2X1 U145 ( .A(n320), .B(n318), .Y(n234) );
  NOR2X1 U146 ( .A(n321), .B(n318), .Y(n235) );
  NOR2X1 U147 ( .A(n322), .B(n318), .Y(n236) );
  NOR2X1 U148 ( .A(n323), .B(n318), .Y(n237) );
  NOR2X1 U149 ( .A(n324), .B(n318), .Y(n238) );
  NOR2X1 U150 ( .A(n325), .B(n318), .Y(n239) );
  NOR2X1 U151 ( .A(n326), .B(n318), .Y(n240) );
  NOR2X1 U152 ( .A(n327), .B(n318), .Y(n241) );
  NOR2X1 U153 ( .A(n328), .B(n318), .Y(n242) );
  NOR2X1 U154 ( .A(n313), .B(n318), .Y(n243) );
  NOR2X1 U155 ( .A(n320), .B(n319), .Y(n244) );
  NOR2X1 U156 ( .A(n321), .B(n319), .Y(n245) );
  NOR2X1 U157 ( .A(n322), .B(n319), .Y(n246) );
  NOR2X1 U158 ( .A(n323), .B(n319), .Y(n247) );
  NOR2X1 U159 ( .A(n324), .B(n319), .Y(n248) );
  NOR2X1 U160 ( .A(n325), .B(n319), .Y(n249) );
  NOR2X1 U161 ( .A(n326), .B(n319), .Y(n250) );
  NOR2X1 U162 ( .A(n327), .B(n319), .Y(n251) );
  NOR2X1 U163 ( .A(n328), .B(n319), .Y(n252) );
  NOR2X1 U164 ( .A(n313), .B(n319), .Y(n253) );
  NOR2X1 U165 ( .A(n321), .B(n320), .Y(n254) );
  NOR2X1 U166 ( .A(n322), .B(n320), .Y(n255) );
  NOR2X1 U167 ( .A(n323), .B(n320), .Y(n256) );
  NOR2X1 U168 ( .A(n324), .B(n320), .Y(n257) );
  NOR2X1 U169 ( .A(n325), .B(n320), .Y(n258) );
  NOR2X1 U170 ( .A(n326), .B(n320), .Y(n259) );
  NOR2X1 U171 ( .A(n327), .B(n320), .Y(n260) );
  NOR2X1 U172 ( .A(n328), .B(n320), .Y(n261) );
  NOR2X1 U173 ( .A(n313), .B(n320), .Y(n262) );
  NOR2X1 U174 ( .A(n322), .B(n321), .Y(n263) );
  NOR2X1 U175 ( .A(n323), .B(n321), .Y(n264) );
  NOR2X1 U176 ( .A(n324), .B(n321), .Y(n265) );
  NOR2X1 U177 ( .A(n325), .B(n321), .Y(n266) );
  NOR2X1 U178 ( .A(n326), .B(n321), .Y(n267) );
  NOR2X1 U179 ( .A(n327), .B(n321), .Y(n268) );
  NOR2X1 U180 ( .A(n328), .B(n321), .Y(n269) );
  NOR2X1 U181 ( .A(n313), .B(n321), .Y(n270) );
  NOR2X1 U182 ( .A(n323), .B(n322), .Y(n271) );
  NOR2X1 U183 ( .A(n324), .B(n322), .Y(n272) );
  NOR2X1 U184 ( .A(n325), .B(n322), .Y(n273) );
  NOR2X1 U185 ( .A(n326), .B(n322), .Y(n274) );
  NOR2X1 U186 ( .A(n327), .B(n322), .Y(n275) );
  NOR2X1 U187 ( .A(n328), .B(n322), .Y(n276) );
  NOR2X1 U188 ( .A(n313), .B(n322), .Y(n277) );
  NOR2X1 U189 ( .A(n324), .B(n323), .Y(n278) );
  NOR2X1 U190 ( .A(n325), .B(n323), .Y(n279) );
  NOR2X1 U191 ( .A(n326), .B(n323), .Y(n280) );
  NOR2X1 U192 ( .A(n327), .B(n323), .Y(n281) );
  NOR2X1 U193 ( .A(n328), .B(n323), .Y(n282) );
  NOR2X1 U194 ( .A(n313), .B(n323), .Y(n283) );
  NOR2X1 U195 ( .A(n325), .B(n324), .Y(n284) );
  NOR2X1 U196 ( .A(n326), .B(n324), .Y(n285) );
  NOR2X1 U197 ( .A(n327), .B(n324), .Y(n286) );
  NOR2X1 U198 ( .A(n328), .B(n324), .Y(n287) );
  NOR2X1 U199 ( .A(n313), .B(n324), .Y(n288) );
  NOR2X1 U200 ( .A(n326), .B(n325), .Y(n289) );
  NOR2X1 U201 ( .A(n327), .B(n325), .Y(n290) );
  NOR2X1 U202 ( .A(n328), .B(n325), .Y(n291) );
  NOR2X1 U203 ( .A(n313), .B(n325), .Y(n292) );
  NOR2X1 U204 ( .A(n327), .B(n326), .Y(n293) );
  NOR2X1 U205 ( .A(n328), .B(n326), .Y(n294) );
  NOR2X1 U206 ( .A(n313), .B(n326), .Y(n295) );
  NOR2X1 U207 ( .A(n328), .B(n327), .Y(n296) );
  NOR2X1 U208 ( .A(n313), .B(n327), .Y(n297) );
  NOR2X1 U209 ( .A(n313), .B(n328), .Y(n298) );
  CLKINVX1 U243 ( .A(a[0]), .Y(n313) );
  CLKINVX1 U244 ( .A(a[1]), .Y(n328) );
  CLKINVX1 U245 ( .A(a[2]), .Y(n327) );
  CLKINVX1 U246 ( .A(a[3]), .Y(n326) );
  CLKINVX1 U247 ( .A(a[4]), .Y(n325) );
  CLKINVX1 U248 ( .A(a[5]), .Y(n324) );
  CLKINVX1 U249 ( .A(a[6]), .Y(n323) );
  CLKINVX1 U250 ( .A(a[7]), .Y(n322) );
  CLKINVX1 U251 ( .A(a[8]), .Y(n321) );
  CLKINVX1 U252 ( .A(a[9]), .Y(n320) );
  CLKINVX1 U253 ( .A(a[10]), .Y(n319) );
  CLKINVX1 U254 ( .A(a[11]), .Y(n318) );
  CLKINVX1 U255 ( .A(a[12]), .Y(n317) );
  CLKINVX1 U256 ( .A(a[13]), .Y(n316) );
  CLKINVX1 U257 ( .A(a[14]), .Y(n315) );
  CLKBUFX3 U258 ( .A(a[0]), .Y(product_0_) );
  CLKINVX1 U259 ( .A(a[15]), .Y(n314) );
endmodule


module FAS_DW_mult_tc_23 ( a, product_31_, product_30_, product_29_, 
        product_28_, product_27_, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_, product_14_, 
        product_13_, product_12_, product_11_, product_10_, product_9_, 
        product_8_, product_7_, product_6_, product_5_, product_4_, product_3_, 
        product_2_, product_0_ );
  input [15:0] a;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_0_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328;

  CLKINVX1 U1 ( .A(n1), .Y(product_31_) );
  ADDFXL U2 ( .A(n179), .B(a[15]), .CI(n2), .CO(n1), .S(product_30_) );
  ADDFXL U3 ( .A(n30), .B(n180), .CI(n3), .CO(n2), .S(product_29_) );
  ADDFXL U4 ( .A(n32), .B(n31), .CI(n4), .CO(n3), .S(product_28_) );
  ADDFXL U5 ( .A(n35), .B(n33), .CI(n5), .CO(n4), .S(product_27_) );
  ADDFXL U6 ( .A(n38), .B(n36), .CI(n6), .CO(n5), .S(product_26_) );
  ADDFXL U7 ( .A(n41), .B(n39), .CI(n7), .CO(n6), .S(product_25_) );
  ADDFXL U8 ( .A(n42), .B(n46), .CI(n8), .CO(n7), .S(product_24_) );
  ADDFXL U9 ( .A(n51), .B(n47), .CI(n9), .CO(n8), .S(product_23_) );
  ADDFXL U10 ( .A(n52), .B(n57), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U11 ( .A(n58), .B(n63), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U12 ( .A(n64), .B(n71), .CI(n12), .CO(n11), .S(product_20_) );
  ADDFXL U13 ( .A(n79), .B(n72), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFXL U14 ( .A(n80), .B(n88), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFXL U15 ( .A(n89), .B(n97), .CI(n15), .CO(n14), .S(product_17_) );
  ADDFXL U16 ( .A(n98), .B(n108), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFXL U17 ( .A(n109), .B(n118), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFXL U18 ( .A(n119), .B(n128), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFXL U19 ( .A(n129), .B(n136), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFXL U20 ( .A(n137), .B(n144), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFXL U21 ( .A(n145), .B(n151), .CI(n21), .CO(n20), .S(product_11_) );
  ADDFXL U22 ( .A(n152), .B(n158), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFXL U23 ( .A(n159), .B(n163), .CI(n23), .CO(n22), .S(product_9_) );
  ADDFXL U24 ( .A(n164), .B(n167), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFXL U25 ( .A(n168), .B(n171), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFXL U26 ( .A(n172), .B(n174), .CI(n26), .CO(n25), .S(product_6_) );
  ADDFXL U27 ( .A(n176), .B(n177), .CI(n27), .CO(n26), .S(product_5_) );
  ADDFXL U28 ( .A(n178), .B(n295), .CI(n28), .CO(n27), .S(product_4_) );
  ADDHXL U29 ( .A(n297), .B(n29), .CO(n28), .S(product_3_) );
  ADDHXL U30 ( .A(a[1]), .B(n298), .CO(n29), .S(product_2_) );
  ADDFXL U31 ( .A(n194), .B(a[14]), .CI(n181), .CO(n30), .S(n31) );
  ADDFXL U32 ( .A(n182), .B(n195), .CI(n34), .CO(n32), .S(n33) );
  CMPR42X1 U33 ( .A(a[13]), .B(n196), .C(n208), .D(n183), .ICI(n37), .S(n36), 
        .ICO(n34), .CO(n35) );
  CMPR42X1 U34 ( .A(n209), .B(n197), .C(n184), .D(n43), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U35 ( .A(n221), .B(n210), .C(n44), .D(n48), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFXL U36 ( .A(n198), .B(a[12]), .CI(n185), .CO(n43), .S(n44) );
  CMPR42X1 U37 ( .A(n199), .B(n53), .C(n49), .D(n54), .ICI(n50), .S(n47), 
        .ICO(n45), .CO(n46) );
  ADDFXL U38 ( .A(n211), .B(n222), .CI(n186), .CO(n48), .S(n49) );
  CMPR42X1 U39 ( .A(n223), .B(n212), .C(n60), .D(n55), .ICI(n56), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U40 ( .A(a[11]), .B(n200), .C(n233), .D(n187), .ICI(n59), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U41 ( .A(n201), .B(n68), .C(n66), .D(n61), .ICI(n62), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U42 ( .A(n213), .B(n234), .C(n224), .D(n188), .ICI(n65), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U43 ( .A(n69), .B(n76), .C(n74), .D(n67), .ICI(n70), .S(n64), .ICO(
        n62), .CO(n63) );
  CMPR42X1 U44 ( .A(n225), .B(n244), .C(n235), .D(n214), .ICI(n73), .S(n67), 
        .ICO(n65), .CO(n66) );
  ADDFXL U45 ( .A(n202), .B(a[10]), .CI(n189), .CO(n68), .S(n69) );
  CMPR42X1 U46 ( .A(n77), .B(n85), .C(n82), .D(n75), .ICI(n78), .S(n72), .ICO(
        n70), .CO(n71) );
  CMPR42X1 U47 ( .A(n236), .B(n215), .C(n226), .D(n84), .ICI(n81), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFXL U48 ( .A(n203), .B(n245), .CI(n190), .CO(n76), .S(n77) );
  CMPR42X1 U49 ( .A(n94), .B(n91), .C(n86), .D(n83), .ICI(n87), .S(n80), .ICO(
        n78), .CO(n79) );
  CMPR42X1 U50 ( .A(n227), .B(n246), .C(n237), .D(n216), .ICI(n90), .S(n83), 
        .ICO(n81), .CO(n82) );
  CMPR42X1 U51 ( .A(a[9]), .B(n204), .C(n254), .D(n191), .ICI(n93), .S(n86), 
        .ICO(n84), .CO(n85) );
  CMPR42X1 U52 ( .A(n103), .B(n100), .C(n92), .D(n95), .ICI(n96), .S(n89), 
        .ICO(n87), .CO(n88) );
  CMPR42X1 U53 ( .A(n228), .B(n247), .C(n238), .D(n217), .ICI(n99), .S(n92), 
        .ICO(n90), .CO(n91) );
  CMPR42X1 U54 ( .A(n255), .B(n205), .C(n192), .D(n105), .ICI(n102), .S(n95), 
        .ICO(n93), .CO(n94) );
  CMPR42X1 U55 ( .A(n113), .B(n111), .C(n101), .D(n104), .ICI(n107), .S(n98), 
        .ICO(n96), .CO(n97) );
  CMPR42X1 U56 ( .A(n248), .B(n218), .C(n229), .D(n239), .ICI(n115), .S(n101), 
        .ICO(n99), .CO(n100) );
  CMPR42X1 U57 ( .A(n256), .B(n206), .C(n193), .D(n106), .ICI(n110), .S(n104), 
        .ICO(n102), .CO(n103) );
  XNOR2X1 U58 ( .A(n263), .B(a[8]), .Y(n106) );
  OR2X1 U59 ( .A(n263), .B(a[8]), .Y(n105) );
  CMPR42X1 U60 ( .A(n123), .B(n114), .C(n121), .D(n112), .ICI(n117), .S(n109), 
        .ICO(n107), .CO(n108) );
  CMPR42X1 U61 ( .A(n257), .B(n230), .C(n249), .D(n116), .ICI(n120), .S(n112), 
        .ICO(n110), .CO(n111) );
  ADDFXL U62 ( .A(n264), .B(n240), .CI(n125), .CO(n113), .S(n114) );
  ADDHXL U63 ( .A(n219), .B(n207), .CO(n115), .S(n116) );
  CMPR42X1 U64 ( .A(n250), .B(n124), .C(n131), .D(n122), .ICI(n127), .S(n119), 
        .ICO(n117), .CO(n118) );
  CMPR42X1 U65 ( .A(n265), .B(n241), .C(n258), .D(n133), .ICI(n130), .S(n122), 
        .ICO(n120), .CO(n121) );
  ADDFXL U66 ( .A(n231), .B(n271), .CI(n126), .CO(n123), .S(n124) );
  ADDHXL U67 ( .A(a[7]), .B(n220), .CO(n125), .S(n126) );
  CMPR42X1 U68 ( .A(n251), .B(n134), .C(n139), .D(n132), .ICI(n135), .S(n129), 
        .ICO(n127), .CO(n128) );
  CMPR42X1 U69 ( .A(n259), .B(n272), .C(n266), .D(n141), .ICI(n138), .S(n132), 
        .ICO(n130), .CO(n131) );
  ADDHXL U70 ( .A(n242), .B(n232), .CO(n133), .S(n134) );
  CMPR42X1 U71 ( .A(n267), .B(n260), .C(n146), .D(n143), .ICI(n140), .S(n137), 
        .ICO(n135), .CO(n136) );
  CMPR42X1 U72 ( .A(n278), .B(n252), .C(n273), .D(n148), .ICI(n142), .S(n140), 
        .ICO(n138), .CO(n139) );
  ADDHXL U73 ( .A(a[6]), .B(n243), .CO(n141), .S(n142) );
  CMPR42X1 U74 ( .A(n279), .B(n149), .C(n150), .D(n153), .ICI(n147), .S(n145), 
        .ICO(n143), .CO(n144) );
  ADDFXL U75 ( .A(n274), .B(n268), .CI(n155), .CO(n146), .S(n147) );
  ADDHXL U76 ( .A(n261), .B(n253), .CO(n148), .S(n149) );
  CMPR42X1 U77 ( .A(n280), .B(n275), .C(n160), .D(n157), .ICI(n154), .S(n152), 
        .ICO(n150), .CO(n151) );
  ADDFXL U78 ( .A(n269), .B(n284), .CI(n156), .CO(n153), .S(n154) );
  ADDHXL U79 ( .A(a[5]), .B(n262), .CO(n155), .S(n156) );
  CMPR42X1 U80 ( .A(n285), .B(n281), .C(n165), .D(n161), .ICI(n162), .S(n159), 
        .ICO(n157), .CO(n158) );
  ADDHXL U81 ( .A(n276), .B(n270), .CO(n160), .S(n161) );
  CMPR42X1 U82 ( .A(n289), .B(n282), .C(n286), .D(n169), .ICI(n166), .S(n164), 
        .ICO(n162), .CO(n163) );
  ADDHXL U83 ( .A(a[4]), .B(n277), .CO(n165), .S(n166) );
  ADDFXL U84 ( .A(n173), .B(n287), .CI(n170), .CO(n167), .S(n168) );
  ADDHXL U85 ( .A(n290), .B(n283), .CO(n169), .S(n170) );
  ADDFXL U86 ( .A(n291), .B(n293), .CI(n175), .CO(n171), .S(n172) );
  ADDHXL U87 ( .A(a[3]), .B(n288), .CO(n173), .S(n174) );
  ADDHXL U88 ( .A(n294), .B(n292), .CO(n175), .S(n176) );
  ADDHXL U89 ( .A(a[2]), .B(n296), .CO(n177), .S(n178) );
  OR2X1 U90 ( .A(n315), .B(n314), .Y(n179) );
  OR2X1 U91 ( .A(n316), .B(n314), .Y(n180) );
  OR2X1 U92 ( .A(n317), .B(n314), .Y(n181) );
  OR2X1 U93 ( .A(n318), .B(n314), .Y(n182) );
  OR2X1 U94 ( .A(n319), .B(n314), .Y(n183) );
  OR2X1 U95 ( .A(n320), .B(n314), .Y(n184) );
  OR2X1 U96 ( .A(n321), .B(n314), .Y(n185) );
  OR2X1 U97 ( .A(n322), .B(n314), .Y(n186) );
  OR2X1 U98 ( .A(n323), .B(n314), .Y(n187) );
  OR2X1 U99 ( .A(n324), .B(n314), .Y(n188) );
  OR2X1 U100 ( .A(n325), .B(n314), .Y(n189) );
  OR2X1 U101 ( .A(n326), .B(n314), .Y(n190) );
  OR2X1 U102 ( .A(n327), .B(n314), .Y(n191) );
  OR2X1 U103 ( .A(n328), .B(n314), .Y(n192) );
  OR2X1 U104 ( .A(n313), .B(n314), .Y(n193) );
  NOR2X1 U105 ( .A(n316), .B(n315), .Y(n194) );
  NOR2X1 U106 ( .A(n317), .B(n315), .Y(n195) );
  NOR2X1 U107 ( .A(n318), .B(n315), .Y(n196) );
  NOR2X1 U108 ( .A(n319), .B(n315), .Y(n197) );
  NOR2X1 U109 ( .A(n320), .B(n315), .Y(n198) );
  NOR2X1 U110 ( .A(n321), .B(n315), .Y(n199) );
  NOR2X1 U111 ( .A(n322), .B(n315), .Y(n200) );
  NOR2X1 U112 ( .A(n323), .B(n315), .Y(n201) );
  NOR2X1 U113 ( .A(n324), .B(n315), .Y(n202) );
  NOR2X1 U114 ( .A(n325), .B(n315), .Y(n203) );
  NOR2X1 U115 ( .A(n326), .B(n315), .Y(n204) );
  NOR2X1 U116 ( .A(n327), .B(n315), .Y(n205) );
  NOR2X1 U117 ( .A(n328), .B(n315), .Y(n206) );
  NOR2X1 U118 ( .A(n313), .B(n315), .Y(n207) );
  NOR2X1 U119 ( .A(n317), .B(n316), .Y(n208) );
  NOR2X1 U120 ( .A(n318), .B(n316), .Y(n209) );
  NOR2X1 U121 ( .A(n319), .B(n316), .Y(n210) );
  NOR2X1 U122 ( .A(n320), .B(n316), .Y(n211) );
  NOR2X1 U123 ( .A(n321), .B(n316), .Y(n212) );
  NOR2X1 U124 ( .A(n322), .B(n316), .Y(n213) );
  NOR2X1 U125 ( .A(n323), .B(n316), .Y(n214) );
  NOR2X1 U126 ( .A(n324), .B(n316), .Y(n215) );
  NOR2X1 U127 ( .A(n325), .B(n316), .Y(n216) );
  NOR2X1 U128 ( .A(n326), .B(n316), .Y(n217) );
  NOR2X1 U129 ( .A(n327), .B(n316), .Y(n218) );
  NOR2X1 U130 ( .A(n328), .B(n316), .Y(n219) );
  NOR2X1 U131 ( .A(n313), .B(n316), .Y(n220) );
  NOR2X1 U132 ( .A(n318), .B(n317), .Y(n221) );
  NOR2X1 U133 ( .A(n319), .B(n317), .Y(n222) );
  NOR2X1 U134 ( .A(n320), .B(n317), .Y(n223) );
  NOR2X1 U135 ( .A(n321), .B(n317), .Y(n224) );
  NOR2X1 U136 ( .A(n322), .B(n317), .Y(n225) );
  NOR2X1 U137 ( .A(n323), .B(n317), .Y(n226) );
  NOR2X1 U138 ( .A(n324), .B(n317), .Y(n227) );
  NOR2X1 U139 ( .A(n325), .B(n317), .Y(n228) );
  NOR2X1 U140 ( .A(n326), .B(n317), .Y(n229) );
  NOR2X1 U141 ( .A(n327), .B(n317), .Y(n230) );
  NOR2X1 U142 ( .A(n328), .B(n317), .Y(n231) );
  NOR2X1 U143 ( .A(n313), .B(n317), .Y(n232) );
  NOR2X1 U144 ( .A(n319), .B(n318), .Y(n233) );
  NOR2X1 U145 ( .A(n320), .B(n318), .Y(n234) );
  NOR2X1 U146 ( .A(n321), .B(n318), .Y(n235) );
  NOR2X1 U147 ( .A(n322), .B(n318), .Y(n236) );
  NOR2X1 U148 ( .A(n323), .B(n318), .Y(n237) );
  NOR2X1 U149 ( .A(n324), .B(n318), .Y(n238) );
  NOR2X1 U150 ( .A(n325), .B(n318), .Y(n239) );
  NOR2X1 U151 ( .A(n326), .B(n318), .Y(n240) );
  NOR2X1 U152 ( .A(n327), .B(n318), .Y(n241) );
  NOR2X1 U153 ( .A(n328), .B(n318), .Y(n242) );
  NOR2X1 U154 ( .A(n313), .B(n318), .Y(n243) );
  NOR2X1 U155 ( .A(n320), .B(n319), .Y(n244) );
  NOR2X1 U156 ( .A(n321), .B(n319), .Y(n245) );
  NOR2X1 U157 ( .A(n322), .B(n319), .Y(n246) );
  NOR2X1 U158 ( .A(n323), .B(n319), .Y(n247) );
  NOR2X1 U159 ( .A(n324), .B(n319), .Y(n248) );
  NOR2X1 U160 ( .A(n325), .B(n319), .Y(n249) );
  NOR2X1 U161 ( .A(n326), .B(n319), .Y(n250) );
  NOR2X1 U162 ( .A(n327), .B(n319), .Y(n251) );
  NOR2X1 U163 ( .A(n328), .B(n319), .Y(n252) );
  NOR2X1 U164 ( .A(n313), .B(n319), .Y(n253) );
  NOR2X1 U165 ( .A(n321), .B(n320), .Y(n254) );
  NOR2X1 U166 ( .A(n322), .B(n320), .Y(n255) );
  NOR2X1 U167 ( .A(n323), .B(n320), .Y(n256) );
  NOR2X1 U168 ( .A(n324), .B(n320), .Y(n257) );
  NOR2X1 U169 ( .A(n325), .B(n320), .Y(n258) );
  NOR2X1 U170 ( .A(n326), .B(n320), .Y(n259) );
  NOR2X1 U171 ( .A(n327), .B(n320), .Y(n260) );
  NOR2X1 U172 ( .A(n328), .B(n320), .Y(n261) );
  NOR2X1 U173 ( .A(n313), .B(n320), .Y(n262) );
  NOR2X1 U174 ( .A(n322), .B(n321), .Y(n263) );
  NOR2X1 U175 ( .A(n323), .B(n321), .Y(n264) );
  NOR2X1 U176 ( .A(n324), .B(n321), .Y(n265) );
  NOR2X1 U177 ( .A(n325), .B(n321), .Y(n266) );
  NOR2X1 U178 ( .A(n326), .B(n321), .Y(n267) );
  NOR2X1 U179 ( .A(n327), .B(n321), .Y(n268) );
  NOR2X1 U180 ( .A(n328), .B(n321), .Y(n269) );
  NOR2X1 U181 ( .A(n313), .B(n321), .Y(n270) );
  NOR2X1 U182 ( .A(n323), .B(n322), .Y(n271) );
  NOR2X1 U183 ( .A(n324), .B(n322), .Y(n272) );
  NOR2X1 U184 ( .A(n325), .B(n322), .Y(n273) );
  NOR2X1 U185 ( .A(n326), .B(n322), .Y(n274) );
  NOR2X1 U186 ( .A(n327), .B(n322), .Y(n275) );
  NOR2X1 U187 ( .A(n328), .B(n322), .Y(n276) );
  NOR2X1 U188 ( .A(n313), .B(n322), .Y(n277) );
  NOR2X1 U189 ( .A(n324), .B(n323), .Y(n278) );
  NOR2X1 U190 ( .A(n325), .B(n323), .Y(n279) );
  NOR2X1 U191 ( .A(n326), .B(n323), .Y(n280) );
  NOR2X1 U192 ( .A(n327), .B(n323), .Y(n281) );
  NOR2X1 U193 ( .A(n328), .B(n323), .Y(n282) );
  NOR2X1 U194 ( .A(n313), .B(n323), .Y(n283) );
  NOR2X1 U195 ( .A(n325), .B(n324), .Y(n284) );
  NOR2X1 U196 ( .A(n326), .B(n324), .Y(n285) );
  NOR2X1 U197 ( .A(n327), .B(n324), .Y(n286) );
  NOR2X1 U198 ( .A(n328), .B(n324), .Y(n287) );
  NOR2X1 U199 ( .A(n313), .B(n324), .Y(n288) );
  NOR2X1 U200 ( .A(n326), .B(n325), .Y(n289) );
  NOR2X1 U201 ( .A(n327), .B(n325), .Y(n290) );
  NOR2X1 U202 ( .A(n328), .B(n325), .Y(n291) );
  NOR2X1 U203 ( .A(n313), .B(n325), .Y(n292) );
  NOR2X1 U204 ( .A(n327), .B(n326), .Y(n293) );
  NOR2X1 U205 ( .A(n328), .B(n326), .Y(n294) );
  NOR2X1 U206 ( .A(n313), .B(n326), .Y(n295) );
  NOR2X1 U207 ( .A(n328), .B(n327), .Y(n296) );
  NOR2X1 U208 ( .A(n313), .B(n327), .Y(n297) );
  NOR2X1 U209 ( .A(n313), .B(n328), .Y(n298) );
  CLKINVX1 U243 ( .A(a[0]), .Y(n313) );
  CLKINVX1 U244 ( .A(a[1]), .Y(n328) );
  CLKINVX1 U245 ( .A(a[2]), .Y(n327) );
  CLKINVX1 U246 ( .A(a[3]), .Y(n326) );
  CLKINVX1 U247 ( .A(a[4]), .Y(n325) );
  CLKINVX1 U248 ( .A(a[5]), .Y(n324) );
  CLKINVX1 U249 ( .A(a[6]), .Y(n323) );
  CLKINVX1 U250 ( .A(a[7]), .Y(n322) );
  CLKINVX1 U251 ( .A(a[8]), .Y(n321) );
  CLKINVX1 U252 ( .A(a[9]), .Y(n320) );
  CLKINVX1 U253 ( .A(a[10]), .Y(n319) );
  CLKINVX1 U254 ( .A(a[11]), .Y(n318) );
  CLKINVX1 U255 ( .A(a[12]), .Y(n317) );
  CLKINVX1 U256 ( .A(a[13]), .Y(n316) );
  CLKINVX1 U257 ( .A(a[14]), .Y(n315) );
  CLKBUFX3 U258 ( .A(a[0]), .Y(product_0_) );
  CLKINVX1 U259 ( .A(a[15]), .Y(n314) );
endmodule


module FAS_DW_mult_tc_24 ( a, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_, product_14_, 
        product_13_, product_12_, product_11_, product_10_, product_9_, 
        product_8_, product_7_, product_6_, product_5_, product_4_, product_3_, 
        product_2_, product_1_ );
  input [15:0] a;
  output product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63;

  CLKINVX1 U2 ( .A(n63), .Y(product_25_) );
  ADDFXL U4 ( .A(a[14]), .B(a[15]), .CI(n3), .CO(product_24_), .S(product_23_)
         );
  ADDFXL U5 ( .A(a[13]), .B(a[15]), .CI(n4), .CO(n3), .S(product_22_) );
  ADDFXL U6 ( .A(n23), .B(a[12]), .CI(n5), .CO(n4), .S(product_21_) );
  ADDFXL U7 ( .A(n25), .B(n24), .CI(n6), .CO(n5), .S(product_20_) );
  ADDFXL U8 ( .A(n27), .B(n26), .CI(n7), .CO(n6), .S(product_19_) );
  ADDFXL U9 ( .A(n30), .B(n28), .CI(n8), .CO(n7), .S(product_18_) );
  ADDFXL U10 ( .A(n31), .B(n33), .CI(n9), .CO(n8), .S(product_17_) );
  ADDFXL U11 ( .A(n36), .B(n34), .CI(n10), .CO(n9), .S(product_16_) );
  ADDFXL U12 ( .A(n37), .B(n39), .CI(n11), .CO(n10), .S(product_15_) );
  ADDFXL U13 ( .A(n40), .B(n42), .CI(n12), .CO(n11), .S(product_14_) );
  ADDFXL U14 ( .A(n43), .B(n45), .CI(n13), .CO(n12), .S(product_13_) );
  ADDFXL U15 ( .A(n46), .B(n48), .CI(n14), .CO(n13), .S(product_12_) );
  ADDFXL U16 ( .A(n49), .B(n51), .CI(n15), .CO(n14), .S(product_11_) );
  ADDFXL U17 ( .A(n52), .B(n53), .CI(n16), .CO(n15), .S(product_10_) );
  ADDFXL U18 ( .A(n54), .B(n57), .CI(n17), .CO(n16), .S(product_9_) );
  ADDFXL U19 ( .A(n58), .B(n59), .CI(n18), .CO(n17), .S(product_8_) );
  ADDFXL U20 ( .A(n60), .B(n61), .CI(n19), .CO(n18), .S(product_7_) );
  ADDFXL U21 ( .A(n62), .B(a[0]), .CI(n20), .CO(n19), .S(product_6_) );
  ADDFXL U22 ( .A(a[4]), .B(a[2]), .CI(n21), .CO(n20), .S(product_5_) );
  ADDFXL U23 ( .A(a[3]), .B(a[1]), .CI(n22), .CO(n21), .S(product_4_) );
  ADDHXL U24 ( .A(a[0]), .B(a[2]), .CO(n22), .S(product_3_) );
  ADDFXL U25 ( .A(a[11]), .B(a[15]), .CI(a[14]), .CO(n23), .S(n24) );
  ADDFXL U26 ( .A(a[10]), .B(a[15]), .CI(a[13]), .CO(n25), .S(n26) );
  ADDFXL U27 ( .A(a[9]), .B(a[12]), .CI(n29), .CO(n27), .S(n28) );
  CMPR42X1 U28 ( .A(a[15]), .B(a[14]), .C(a[8]), .D(a[11]), .ICI(n32), .S(n31), 
        .ICO(n29), .CO(n30) );
  CMPR42X1 U29 ( .A(a[15]), .B(a[13]), .C(a[7]), .D(a[10]), .ICI(n35), .S(n34), 
        .ICO(n32), .CO(n33) );
  CMPR42X1 U30 ( .A(a[9]), .B(a[6]), .C(a[12]), .D(a[14]), .ICI(n38), .S(n37), 
        .ICO(n35), .CO(n36) );
  CMPR42X1 U31 ( .A(a[8]), .B(a[5]), .C(a[11]), .D(a[13]), .ICI(n41), .S(n40), 
        .ICO(n38), .CO(n39) );
  CMPR42X1 U32 ( .A(a[7]), .B(a[4]), .C(a[10]), .D(a[12]), .ICI(n44), .S(n43), 
        .ICO(n41), .CO(n42) );
  CMPR42X1 U33 ( .A(a[6]), .B(a[3]), .C(a[9]), .D(a[11]), .ICI(n47), .S(n46), 
        .ICO(n44), .CO(n45) );
  CMPR42X1 U34 ( .A(a[5]), .B(a[2]), .C(a[8]), .D(a[10]), .ICI(n50), .S(n49), 
        .ICO(n47), .CO(n48) );
  CMPR42X1 U35 ( .A(a[4]), .B(a[1]), .C(a[7]), .D(a[9]), .ICI(n55), .S(n52), 
        .ICO(n50), .CO(n51) );
  ADDFXL U36 ( .A(a[6]), .B(a[8]), .CI(n56), .CO(n53), .S(n54) );
  ADDHXL U37 ( .A(a[3]), .B(a[0]), .CO(n55), .S(n56) );
  ADDFXL U38 ( .A(a[2]), .B(a[7]), .CI(a[5]), .CO(n57), .S(n58) );
  ADDFXL U39 ( .A(a[1]), .B(a[6]), .CI(a[4]), .CO(n59), .S(n60) );
  ADDHXL U40 ( .A(a[5]), .B(a[3]), .CO(n61), .S(n62) );
  CLKBUFX3 U46 ( .A(product_25_), .Y(product_26_) );
  CLKINVX1 U47 ( .A(a[15]), .Y(n63) );
  BUFX2 U48 ( .A(a[0]), .Y(product_1_) );
  BUFX2 U49 ( .A(a[1]), .Y(product_2_) );
endmodule


module FAS_DW_mult_tc_25 ( a, b_17_, b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, 
        b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input [15:0] a;
  input b_17_, b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_, b_8_,
         b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n3, n5, n7, n9, n11, n13, n15, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n697;

  XOR2X1 U51 ( .A(n52), .B(n51), .Y(product_31_) );
  XOR2X1 U52 ( .A(n83), .B(n697), .Y(n51) );
  ADDFXL U53 ( .A(n84), .B(n85), .CI(n53), .CO(n52), .S(product_30_) );
  ADDFXL U54 ( .A(n90), .B(n86), .CI(n54), .CO(n53), .S(product_29_) );
  ADDFXL U55 ( .A(n93), .B(n91), .CI(n55), .CO(n54), .S(product_28_) );
  ADDFXL U56 ( .A(n94), .B(n98), .CI(n56), .CO(n55), .S(product_27_) );
  ADDFXL U57 ( .A(n99), .B(n103), .CI(n57), .CO(n56), .S(product_26_) );
  ADDFXL U58 ( .A(n104), .B(n110), .CI(n58), .CO(n57), .S(product_25_) );
  ADDFXL U59 ( .A(n111), .B(n116), .CI(n59), .CO(n58), .S(product_24_) );
  ADDFXL U60 ( .A(n117), .B(n124), .CI(n60), .CO(n59), .S(product_23_) );
  ADDFXL U61 ( .A(n132), .B(n125), .CI(n61), .CO(n60), .S(product_22_) );
  ADDFXL U62 ( .A(n142), .B(n133), .CI(n62), .CO(n61), .S(product_21_) );
  ADDFXL U63 ( .A(n143), .B(n151), .CI(n63), .CO(n62), .S(product_20_) );
  ADDFXL U64 ( .A(n152), .B(n162), .CI(n64), .CO(n63), .S(product_19_) );
  ADDFXL U65 ( .A(n163), .B(n173), .CI(n65), .CO(n64), .S(product_18_) );
  ADDFXL U66 ( .A(n174), .B(n184), .CI(n66), .CO(n65), .S(product_17_) );
  ADDFXL U67 ( .A(n185), .B(n195), .CI(n67), .CO(n66), .S(product_16_) );
  ADDFXL U68 ( .A(n196), .B(n206), .CI(n68), .CO(n67), .S(product_15_) );
  ADDFXL U69 ( .A(n207), .B(n215), .CI(n69), .CO(n68), .S(product_14_) );
  ADDFXL U70 ( .A(n216), .B(n225), .CI(n70), .CO(n69), .S(product_13_) );
  ADDFXL U71 ( .A(n226), .B(n233), .CI(n71), .CO(n70), .S(product_12_) );
  ADDFXL U72 ( .A(n234), .B(n241), .CI(n72), .CO(n71), .S(product_11_) );
  ADDFXL U73 ( .A(n242), .B(n247), .CI(n73), .CO(n72), .S(product_10_) );
  ADDFXL U74 ( .A(n248), .B(n254), .CI(n74), .CO(n73), .S(product_9_) );
  ADDFXL U75 ( .A(n255), .B(n259), .CI(n75), .CO(n74), .S(product_8_) );
  ADDFXL U76 ( .A(n260), .B(n264), .CI(n76), .CO(n75), .S(product_7_) );
  ADDFXL U77 ( .A(n265), .B(n266), .CI(n77), .CO(n76), .S(product_6_) );
  ADDFXL U78 ( .A(n267), .B(n270), .CI(n78), .CO(n77), .S(product_5_) );
  ADDFXL U79 ( .A(n271), .B(n272), .CI(n79), .CO(n78), .S(product_4_) );
  ADDFXL U80 ( .A(n273), .B(n406), .CI(n80), .CO(n79), .S(product_3_) );
  ADDFXL U81 ( .A(n424), .B(n407), .CI(n81), .CO(n80), .S(product_2_) );
  ADDHXL U82 ( .A(n281), .B(n425), .CO(n81), .S(product_1_) );
  ADDFXL U84 ( .A(n283), .B(n87), .CI(n300), .CO(n83), .S(n84) );
  ADDFXL U85 ( .A(n88), .B(n284), .CI(n89), .CO(n85), .S(n86) );
  CLKINVX1 U86 ( .A(n87), .Y(n88) );
  CMPR42X1 U87 ( .A(n95), .B(n285), .C(n301), .D(n318), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U88 ( .A(n302), .B(n286), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CLKINVX1 U89 ( .A(n95), .Y(n96) );
  CMPR42X1 U90 ( .A(n319), .B(n303), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFXL U91 ( .A(n107), .B(n287), .CI(n335), .CO(n100), .S(n101) );
  CMPR42X1 U92 ( .A(n320), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFXL U93 ( .A(n304), .B(n288), .CI(n108), .CO(n105), .S(n106) );
  CLKINVX1 U94 ( .A(n107), .Y(n108) );
  CMPR42X1 U95 ( .A(n321), .B(n305), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U96 ( .A(n289), .B(n121), .C(n336), .D(n353), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U97 ( .A(n290), .B(n129), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U98 ( .A(n306), .B(n354), .C(n337), .D(n122), .ICI(n126), .S(n120), 
        .ICO(n118), .CO(n119) );
  CLKINVX1 U99 ( .A(n121), .Y(n122) );
  CMPR42X1 U100 ( .A(n137), .B(n130), .C(n135), .D(n128), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U101 ( .A(n307), .B(n338), .C(n322), .D(n139), .ICI(n134), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFXL U102 ( .A(n355), .B(n291), .CI(n372), .CO(n129), .S(n130) );
  CMPR42X1 U103 ( .A(n138), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U104 ( .A(n356), .B(n323), .C(n339), .D(n144), .ICI(n147), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFXL U105 ( .A(n292), .B(n308), .CI(n140), .CO(n137), .S(n138) );
  CLKINVX1 U106 ( .A(n139), .Y(n140) );
  CMPR42X1 U107 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U108 ( .A(n309), .B(n340), .C(n324), .D(n159), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U109 ( .A(n293), .B(n373), .C(n357), .D(n390), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U110 ( .A(n168), .B(n165), .C(n155), .D(n158), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U111 ( .A(n325), .B(n358), .C(n341), .D(n294), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U112 ( .A(n310), .B(n374), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CLKINVX1 U113 ( .A(n159), .Y(n160) );
  CMPR42X1 U114 ( .A(n179), .B(n176), .C(n166), .D(n169), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U115 ( .A(n295), .B(n375), .C(n342), .D(n181), .ICI(n175), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U116 ( .A(n326), .B(n391), .C(n408), .D(n171), .ICI(n178), .S(n169), 
        .ICO(n167), .CO(n168) );
  XNOR2X1 U117 ( .A(n359), .B(n311), .Y(n171) );
  OR2X1 U118 ( .A(n359), .B(n311), .Y(n170) );
  CMPR42X1 U119 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U120 ( .A(n312), .B(n360), .C(n343), .D(n182), .ICI(n186), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U121 ( .A(n327), .B(n392), .C(n376), .D(n192), .ICI(n189), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U122 ( .A(n409), .B(n296), .CO(n181), .S(n182) );
  CMPR42X1 U123 ( .A(n201), .B(n198), .C(n191), .D(n188), .ICI(n194), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U124 ( .A(n313), .B(n328), .C(n361), .D(n193), .ICI(n200), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U125 ( .A(n344), .B(n393), .C(n377), .D(n203), .ICI(n197), .S(n191), 
        .ICO(n189), .CO(n190) );
  ADDHXL U126 ( .A(n410), .B(n297), .CO(n192), .S(n193) );
  CMPR42X1 U127 ( .A(n212), .B(n209), .C(n202), .D(n199), .ICI(n205), .S(n196), 
        .ICO(n194), .CO(n195) );
  CMPR42X1 U128 ( .A(n314), .B(n329), .C(n345), .D(n211), .ICI(n204), .S(n199), 
        .ICO(n197), .CO(n198) );
  CMPR42X1 U129 ( .A(n274), .B(n298), .C(n394), .D(n362), .ICI(n208), .S(n202), 
        .ICO(n200), .CO(n201) );
  ADDHXL U130 ( .A(n411), .B(n378), .CO(n203), .S(n204) );
  CMPR42X1 U131 ( .A(n220), .B(n213), .C(n218), .D(n210), .ICI(n214), .S(n207), 
        .ICO(n205), .CO(n206) );
  CMPR42X1 U132 ( .A(n395), .B(n346), .C(n363), .D(n379), .ICI(n222), .S(n210), 
        .ICO(n208), .CO(n209) );
  CMPR42X1 U133 ( .A(n299), .B(n412), .C(n315), .D(n330), .ICI(n217), .S(n213), 
        .ICO(n211), .CO(n212) );
  CMPR42X1 U134 ( .A(n230), .B(n221), .C(n228), .D(n219), .ICI(n224), .S(n216), 
        .ICO(n214), .CO(n215) );
  CMPR42X1 U135 ( .A(n331), .B(n364), .C(n347), .D(n316), .ICI(n227), .S(n219), 
        .ICO(n217), .CO(n218) );
  ADDFXL U136 ( .A(n396), .B(n275), .CI(n223), .CO(n220), .S(n221) );
  ADDHXL U137 ( .A(n413), .B(n380), .CO(n222), .S(n223) );
  CMPR42X1 U138 ( .A(n365), .B(n235), .C(n236), .D(n229), .ICI(n232), .S(n226), 
        .ICO(n224), .CO(n225) );
  CMPR42X1 U139 ( .A(n397), .B(n348), .C(n381), .D(n238), .ICI(n231), .S(n229), 
        .ICO(n227), .CO(n228) );
  ADDFXL U140 ( .A(n414), .B(n317), .CI(n332), .CO(n230), .S(n231) );
  CMPR42X1 U141 ( .A(n366), .B(n243), .C(n244), .D(n237), .ICI(n240), .S(n234), 
        .ICO(n232), .CO(n233) );
  CMPR42X1 U142 ( .A(n276), .B(n333), .C(n398), .D(n349), .ICI(n239), .S(n237), 
        .ICO(n235), .CO(n236) );
  ADDHXL U143 ( .A(n415), .B(n382), .CO(n238), .S(n239) );
  CMPR42X1 U144 ( .A(n399), .B(n383), .C(n249), .D(n246), .ICI(n245), .S(n242), 
        .ICO(n240), .CO(n241) );
  CMPR42X1 U145 ( .A(n334), .B(n416), .C(n350), .D(n367), .ICI(n251), .S(n245), 
        .ICO(n243), .CO(n244) );
  CMPR42X1 U146 ( .A(n400), .B(n368), .C(n253), .D(n256), .ICI(n250), .S(n248), 
        .ICO(n246), .CO(n247) );
  ADDFXL U147 ( .A(n351), .B(n277), .CI(n252), .CO(n249), .S(n250) );
  ADDHXL U148 ( .A(n417), .B(n384), .CO(n251), .S(n252) );
  CMPR42X1 U149 ( .A(n401), .B(n385), .C(n261), .D(n258), .ICI(n257), .S(n255), 
        .ICO(n253), .CO(n254) );
  ADDFXL U150 ( .A(n418), .B(n352), .CI(n369), .CO(n256), .S(n257) );
  CMPR42X1 U151 ( .A(n278), .B(n370), .C(n402), .D(n263), .ICI(n262), .S(n260), 
        .ICO(n258), .CO(n259) );
  ADDHXL U152 ( .A(n419), .B(n386), .CO(n261), .S(n262) );
  CMPR42X1 U153 ( .A(n371), .B(n420), .C(n387), .D(n403), .ICI(n268), .S(n265), 
        .ICO(n263), .CO(n264) );
  ADDFXL U154 ( .A(n404), .B(n279), .CI(n269), .CO(n266), .S(n267) );
  ADDHXL U155 ( .A(n421), .B(n388), .CO(n268), .S(n269) );
  ADDFXL U156 ( .A(n422), .B(n389), .CI(n405), .CO(n270), .S(n271) );
  ADDHXL U157 ( .A(n423), .B(n280), .CO(n272), .S(n273) );
  OAI22XL U158 ( .A0(n48), .A1(n620), .B0(n32), .B1(n444), .Y(n274) );
  OAI22XL U160 ( .A0(n48), .A1(n428), .B0(n32), .B1(n427), .Y(n283) );
  OAI22XL U161 ( .A0(n48), .A1(n429), .B0(n32), .B1(n428), .Y(n284) );
  OAI22XL U162 ( .A0(n48), .A1(n430), .B0(n32), .B1(n429), .Y(n285) );
  OAI22XL U163 ( .A0(n48), .A1(n431), .B0(n32), .B1(n430), .Y(n286) );
  OAI22XL U164 ( .A0(n48), .A1(n432), .B0(n32), .B1(n431), .Y(n287) );
  OAI22XL U165 ( .A0(n48), .A1(n433), .B0(n32), .B1(n432), .Y(n288) );
  OAI22XL U166 ( .A0(n48), .A1(n434), .B0(n32), .B1(n433), .Y(n289) );
  OAI22XL U167 ( .A0(n47), .A1(n435), .B0(n31), .B1(n434), .Y(n290) );
  OAI22XL U168 ( .A0(n47), .A1(n436), .B0(n31), .B1(n435), .Y(n291) );
  OAI22XL U169 ( .A0(n47), .A1(n437), .B0(n31), .B1(n436), .Y(n292) );
  OAI22XL U170 ( .A0(n47), .A1(n438), .B0(n31), .B1(n437), .Y(n293) );
  OAI22XL U171 ( .A0(n47), .A1(n439), .B0(n31), .B1(n438), .Y(n294) );
  OAI22XL U172 ( .A0(n47), .A1(n440), .B0(n31), .B1(n439), .Y(n295) );
  OAI22XL U173 ( .A0(n47), .A1(n441), .B0(n31), .B1(n440), .Y(n296) );
  OAI22XL U174 ( .A0(n47), .A1(n442), .B0(n31), .B1(n441), .Y(n297) );
  OAI22XL U175 ( .A0(n47), .A1(n443), .B0(n31), .B1(n442), .Y(n298) );
  NOR2BX1 U176 ( .AN(n49), .B(n31), .Y(n299) );
  XNOR2X1 U177 ( .A(n15), .B(n578), .Y(n426) );
  XNOR2X1 U178 ( .A(n15), .B(n579), .Y(n427) );
  XNOR2X1 U179 ( .A(n15), .B(n580), .Y(n428) );
  XNOR2X1 U180 ( .A(n15), .B(n581), .Y(n429) );
  XNOR2X1 U181 ( .A(n15), .B(n582), .Y(n430) );
  XNOR2X1 U182 ( .A(n15), .B(n583), .Y(n431) );
  XNOR2X1 U183 ( .A(n15), .B(n584), .Y(n432) );
  XNOR2X1 U184 ( .A(n15), .B(n585), .Y(n433) );
  XNOR2X1 U185 ( .A(n15), .B(n586), .Y(n434) );
  XNOR2X1 U186 ( .A(n15), .B(n587), .Y(n435) );
  XNOR2X1 U187 ( .A(n15), .B(n588), .Y(n436) );
  XNOR2X1 U188 ( .A(n15), .B(n589), .Y(n437) );
  XNOR2X1 U189 ( .A(n15), .B(n590), .Y(n438) );
  XNOR2X1 U190 ( .A(n15), .B(n591), .Y(n439) );
  XNOR2X1 U191 ( .A(n15), .B(n592), .Y(n440) );
  XNOR2X1 U192 ( .A(n15), .B(n593), .Y(n441) );
  XNOR2X1 U193 ( .A(n15), .B(n594), .Y(n442) );
  XNOR2X1 U194 ( .A(n15), .B(n49), .Y(n443) );
  NAND2BX1 U195 ( .AN(n49), .B(n15), .Y(n444) );
  OAI22XL U196 ( .A0(n46), .A1(n621), .B0(n30), .B1(n463), .Y(n275) );
  AO21X1 U197 ( .A0(n46), .A1(n30), .B0(n445), .Y(n300) );
  OAI22XL U198 ( .A0(n46), .A1(n446), .B0(n30), .B1(n445), .Y(n87) );
  OAI22XL U199 ( .A0(n46), .A1(n447), .B0(n30), .B1(n446), .Y(n301) );
  OAI22XL U200 ( .A0(n46), .A1(n448), .B0(n30), .B1(n447), .Y(n302) );
  OAI22XL U201 ( .A0(n46), .A1(n449), .B0(n30), .B1(n448), .Y(n303) );
  OAI22XL U202 ( .A0(n46), .A1(n450), .B0(n30), .B1(n449), .Y(n304) );
  OAI22XL U203 ( .A0(n46), .A1(n451), .B0(n30), .B1(n450), .Y(n305) );
  OAI22XL U204 ( .A0(n46), .A1(n452), .B0(n30), .B1(n451), .Y(n306) );
  OAI22XL U205 ( .A0(n46), .A1(n453), .B0(n30), .B1(n452), .Y(n307) );
  OAI22XL U206 ( .A0(n45), .A1(n454), .B0(n29), .B1(n453), .Y(n308) );
  OAI22XL U207 ( .A0(n45), .A1(n455), .B0(n29), .B1(n454), .Y(n309) );
  OAI22XL U208 ( .A0(n45), .A1(n456), .B0(n29), .B1(n455), .Y(n310) );
  OAI22XL U209 ( .A0(n45), .A1(n457), .B0(n29), .B1(n456), .Y(n311) );
  OAI22XL U210 ( .A0(n45), .A1(n458), .B0(n29), .B1(n457), .Y(n312) );
  OAI22XL U211 ( .A0(n45), .A1(n459), .B0(n29), .B1(n458), .Y(n313) );
  OAI22XL U212 ( .A0(n45), .A1(n460), .B0(n29), .B1(n459), .Y(n314) );
  OAI22XL U213 ( .A0(n45), .A1(n461), .B0(n29), .B1(n460), .Y(n315) );
  OAI22XL U214 ( .A0(n45), .A1(n462), .B0(n29), .B1(n461), .Y(n316) );
  NOR2BX1 U215 ( .AN(n49), .B(n29), .Y(n317) );
  XNOR2X1 U216 ( .A(n13), .B(n578), .Y(n445) );
  XNOR2X1 U217 ( .A(n13), .B(n579), .Y(n446) );
  XNOR2X1 U218 ( .A(n13), .B(n580), .Y(n447) );
  XNOR2X1 U219 ( .A(n13), .B(n581), .Y(n448) );
  XNOR2X1 U220 ( .A(n13), .B(n582), .Y(n449) );
  XNOR2X1 U221 ( .A(n13), .B(n583), .Y(n450) );
  XNOR2X1 U222 ( .A(n13), .B(n584), .Y(n451) );
  XNOR2X1 U223 ( .A(n13), .B(n585), .Y(n452) );
  XNOR2X1 U224 ( .A(n13), .B(n586), .Y(n453) );
  XNOR2X1 U225 ( .A(n13), .B(n587), .Y(n454) );
  XNOR2X1 U226 ( .A(n13), .B(n588), .Y(n455) );
  XNOR2X1 U227 ( .A(n13), .B(n589), .Y(n456) );
  XNOR2X1 U228 ( .A(n13), .B(n590), .Y(n457) );
  XNOR2X1 U229 ( .A(n13), .B(n591), .Y(n458) );
  XNOR2X1 U230 ( .A(n13), .B(n592), .Y(n459) );
  XNOR2X1 U231 ( .A(n13), .B(n593), .Y(n460) );
  XNOR2X1 U232 ( .A(n13), .B(n594), .Y(n461) );
  XNOR2X1 U233 ( .A(n13), .B(n49), .Y(n462) );
  NAND2BX1 U234 ( .AN(n49), .B(n13), .Y(n463) );
  OAI22XL U235 ( .A0(n44), .A1(n622), .B0(n28), .B1(n482), .Y(n276) );
  AO21X1 U236 ( .A0(n44), .A1(n28), .B0(n464), .Y(n318) );
  OAI22XL U237 ( .A0(n44), .A1(n465), .B0(n28), .B1(n464), .Y(n95) );
  OAI22XL U238 ( .A0(n44), .A1(n466), .B0(n28), .B1(n465), .Y(n319) );
  OAI22XL U239 ( .A0(n44), .A1(n467), .B0(n28), .B1(n466), .Y(n320) );
  OAI22XL U240 ( .A0(n44), .A1(n468), .B0(n28), .B1(n467), .Y(n321) );
  OAI22XL U241 ( .A0(n44), .A1(n469), .B0(n28), .B1(n468), .Y(n121) );
  OAI22XL U242 ( .A0(n44), .A1(n470), .B0(n28), .B1(n469), .Y(n322) );
  OAI22XL U243 ( .A0(n44), .A1(n471), .B0(n28), .B1(n470), .Y(n323) );
  OAI22XL U244 ( .A0(n44), .A1(n472), .B0(n28), .B1(n471), .Y(n324) );
  OAI22XL U245 ( .A0(n43), .A1(n473), .B0(n27), .B1(n472), .Y(n325) );
  OAI22XL U246 ( .A0(n43), .A1(n474), .B0(n27), .B1(n473), .Y(n326) );
  OAI22XL U247 ( .A0(n43), .A1(n475), .B0(n27), .B1(n474), .Y(n327) );
  OAI22XL U248 ( .A0(n43), .A1(n476), .B0(n27), .B1(n475), .Y(n328) );
  OAI22XL U249 ( .A0(n43), .A1(n477), .B0(n27), .B1(n476), .Y(n329) );
  OAI22XL U250 ( .A0(n43), .A1(n478), .B0(n27), .B1(n477), .Y(n330) );
  OAI22XL U251 ( .A0(n43), .A1(n479), .B0(n27), .B1(n478), .Y(n331) );
  OAI22XL U252 ( .A0(n43), .A1(n480), .B0(n27), .B1(n479), .Y(n332) );
  OAI22XL U253 ( .A0(n43), .A1(n481), .B0(n27), .B1(n480), .Y(n333) );
  NOR2BX1 U254 ( .AN(n49), .B(n27), .Y(n334) );
  XNOR2X1 U255 ( .A(n11), .B(n578), .Y(n464) );
  XNOR2X1 U256 ( .A(n11), .B(n579), .Y(n465) );
  XNOR2X1 U257 ( .A(n11), .B(n580), .Y(n466) );
  XNOR2X1 U258 ( .A(n11), .B(n581), .Y(n467) );
  XNOR2X1 U259 ( .A(n11), .B(n582), .Y(n468) );
  XNOR2X1 U260 ( .A(n11), .B(n583), .Y(n469) );
  XNOR2X1 U261 ( .A(n11), .B(n584), .Y(n470) );
  XNOR2X1 U262 ( .A(n11), .B(n585), .Y(n471) );
  XNOR2X1 U263 ( .A(n11), .B(n586), .Y(n472) );
  XNOR2X1 U264 ( .A(n11), .B(n587), .Y(n473) );
  XNOR2X1 U265 ( .A(n11), .B(n588), .Y(n474) );
  XNOR2X1 U266 ( .A(n11), .B(n589), .Y(n475) );
  XNOR2X1 U267 ( .A(n11), .B(n590), .Y(n476) );
  XNOR2X1 U268 ( .A(n11), .B(n591), .Y(n477) );
  XNOR2X1 U269 ( .A(n11), .B(n592), .Y(n478) );
  XNOR2X1 U270 ( .A(n11), .B(n593), .Y(n479) );
  XNOR2X1 U271 ( .A(n11), .B(n594), .Y(n480) );
  XNOR2X1 U272 ( .A(n11), .B(n49), .Y(n481) );
  NAND2BX1 U273 ( .AN(n49), .B(n11), .Y(n482) );
  OAI22XL U274 ( .A0(n42), .A1(n623), .B0(n26), .B1(n501), .Y(n277) );
  AO21X1 U275 ( .A0(n42), .A1(n26), .B0(n483), .Y(n335) );
  OAI22XL U276 ( .A0(n42), .A1(n484), .B0(n26), .B1(n483), .Y(n107) );
  OAI22XL U277 ( .A0(n42), .A1(n485), .B0(n26), .B1(n484), .Y(n336) );
  OAI22XL U278 ( .A0(n42), .A1(n486), .B0(n26), .B1(n485), .Y(n337) );
  OAI22XL U279 ( .A0(n42), .A1(n487), .B0(n26), .B1(n486), .Y(n338) );
  OAI22XL U280 ( .A0(n42), .A1(n488), .B0(n26), .B1(n487), .Y(n339) );
  OAI22XL U281 ( .A0(n42), .A1(n489), .B0(n26), .B1(n488), .Y(n340) );
  OAI22XL U282 ( .A0(n42), .A1(n490), .B0(n26), .B1(n489), .Y(n341) );
  OAI22XL U283 ( .A0(n42), .A1(n491), .B0(n26), .B1(n490), .Y(n342) );
  OAI22XL U284 ( .A0(n41), .A1(n492), .B0(n25), .B1(n491), .Y(n343) );
  OAI22XL U285 ( .A0(n41), .A1(n493), .B0(n25), .B1(n492), .Y(n344) );
  OAI22XL U286 ( .A0(n41), .A1(n494), .B0(n25), .B1(n493), .Y(n345) );
  OAI22XL U287 ( .A0(n41), .A1(n495), .B0(n25), .B1(n494), .Y(n346) );
  OAI22XL U288 ( .A0(n41), .A1(n496), .B0(n25), .B1(n495), .Y(n347) );
  OAI22XL U289 ( .A0(n41), .A1(n497), .B0(n25), .B1(n496), .Y(n348) );
  OAI22XL U290 ( .A0(n41), .A1(n498), .B0(n25), .B1(n497), .Y(n349) );
  OAI22XL U291 ( .A0(n41), .A1(n499), .B0(n25), .B1(n498), .Y(n350) );
  OAI22XL U292 ( .A0(n41), .A1(n500), .B0(n25), .B1(n499), .Y(n351) );
  NOR2BX1 U293 ( .AN(n49), .B(n25), .Y(n352) );
  XNOR2X1 U294 ( .A(n9), .B(n578), .Y(n483) );
  XNOR2X1 U295 ( .A(n9), .B(n579), .Y(n484) );
  XNOR2X1 U296 ( .A(n9), .B(n580), .Y(n485) );
  XNOR2X1 U297 ( .A(n9), .B(n581), .Y(n486) );
  XNOR2X1 U298 ( .A(n9), .B(n582), .Y(n487) );
  XNOR2X1 U299 ( .A(n9), .B(n583), .Y(n488) );
  XNOR2X1 U300 ( .A(n9), .B(n584), .Y(n489) );
  XNOR2X1 U301 ( .A(n9), .B(n585), .Y(n490) );
  XNOR2X1 U302 ( .A(n9), .B(n586), .Y(n491) );
  XNOR2X1 U303 ( .A(n9), .B(n587), .Y(n492) );
  XNOR2X1 U304 ( .A(n9), .B(n588), .Y(n493) );
  XNOR2X1 U305 ( .A(n9), .B(n589), .Y(n494) );
  XNOR2X1 U306 ( .A(n9), .B(n590), .Y(n495) );
  XNOR2X1 U307 ( .A(n9), .B(n591), .Y(n496) );
  XNOR2X1 U308 ( .A(n9), .B(n592), .Y(n497) );
  XNOR2X1 U309 ( .A(n9), .B(n593), .Y(n498) );
  XNOR2X1 U310 ( .A(n9), .B(n594), .Y(n499) );
  XNOR2X1 U311 ( .A(n9), .B(n49), .Y(n500) );
  NAND2BX1 U312 ( .AN(n49), .B(n9), .Y(n501) );
  OAI22XL U313 ( .A0(n40), .A1(n624), .B0(n24), .B1(n520), .Y(n278) );
  AO21X1 U314 ( .A0(n40), .A1(n24), .B0(n502), .Y(n353) );
  OAI22XL U315 ( .A0(n40), .A1(n503), .B0(n24), .B1(n502), .Y(n354) );
  OAI22XL U316 ( .A0(n40), .A1(n504), .B0(n24), .B1(n503), .Y(n355) );
  OAI22XL U317 ( .A0(n40), .A1(n505), .B0(n24), .B1(n504), .Y(n356) );
  OAI22XL U318 ( .A0(n40), .A1(n506), .B0(n24), .B1(n505), .Y(n357) );
  OAI22XL U319 ( .A0(n40), .A1(n507), .B0(n24), .B1(n506), .Y(n358) );
  OAI22XL U320 ( .A0(n40), .A1(n508), .B0(n24), .B1(n507), .Y(n359) );
  OAI22XL U321 ( .A0(n40), .A1(n509), .B0(n24), .B1(n508), .Y(n360) );
  OAI22XL U322 ( .A0(n40), .A1(n510), .B0(n24), .B1(n509), .Y(n361) );
  OAI22XL U323 ( .A0(n39), .A1(n511), .B0(n23), .B1(n510), .Y(n362) );
  OAI22XL U324 ( .A0(n39), .A1(n512), .B0(n23), .B1(n511), .Y(n363) );
  OAI22XL U325 ( .A0(n39), .A1(n513), .B0(n23), .B1(n512), .Y(n364) );
  OAI22XL U326 ( .A0(n39), .A1(n514), .B0(n23), .B1(n513), .Y(n365) );
  OAI22XL U327 ( .A0(n39), .A1(n515), .B0(n23), .B1(n514), .Y(n366) );
  OAI22XL U328 ( .A0(n39), .A1(n516), .B0(n23), .B1(n515), .Y(n367) );
  OAI22XL U329 ( .A0(n39), .A1(n517), .B0(n23), .B1(n516), .Y(n368) );
  OAI22XL U330 ( .A0(n39), .A1(n518), .B0(n23), .B1(n517), .Y(n369) );
  OAI22XL U331 ( .A0(n39), .A1(n519), .B0(n23), .B1(n518), .Y(n370) );
  NOR2BX1 U332 ( .AN(n49), .B(n23), .Y(n371) );
  XNOR2X1 U333 ( .A(n7), .B(n578), .Y(n502) );
  XNOR2X1 U334 ( .A(n7), .B(n579), .Y(n503) );
  XNOR2X1 U335 ( .A(n7), .B(n580), .Y(n504) );
  XNOR2X1 U336 ( .A(n7), .B(n581), .Y(n505) );
  XNOR2X1 U337 ( .A(n7), .B(n582), .Y(n506) );
  XNOR2X1 U338 ( .A(n7), .B(n583), .Y(n507) );
  XNOR2X1 U339 ( .A(n7), .B(n584), .Y(n508) );
  XNOR2X1 U340 ( .A(n7), .B(n585), .Y(n509) );
  XNOR2X1 U341 ( .A(n7), .B(n586), .Y(n510) );
  XNOR2X1 U342 ( .A(n7), .B(n587), .Y(n511) );
  XNOR2X1 U343 ( .A(n7), .B(n588), .Y(n512) );
  XNOR2X1 U344 ( .A(n7), .B(n589), .Y(n513) );
  XNOR2X1 U345 ( .A(n7), .B(n590), .Y(n514) );
  XNOR2X1 U346 ( .A(n7), .B(n591), .Y(n515) );
  XNOR2X1 U347 ( .A(n7), .B(n592), .Y(n516) );
  XNOR2X1 U348 ( .A(n7), .B(n593), .Y(n517) );
  XNOR2X1 U349 ( .A(n7), .B(n594), .Y(n518) );
  XNOR2X1 U350 ( .A(n7), .B(n49), .Y(n519) );
  NAND2BX1 U351 ( .AN(n49), .B(n7), .Y(n520) );
  OAI22XL U352 ( .A0(n38), .A1(n625), .B0(n22), .B1(n539), .Y(n279) );
  AO21X1 U353 ( .A0(n38), .A1(n22), .B0(n521), .Y(n372) );
  OAI22XL U354 ( .A0(n38), .A1(n522), .B0(n22), .B1(n521), .Y(n139) );
  OAI22XL U355 ( .A0(n38), .A1(n523), .B0(n22), .B1(n522), .Y(n373) );
  OAI22XL U356 ( .A0(n38), .A1(n524), .B0(n22), .B1(n523), .Y(n374) );
  OAI22XL U357 ( .A0(n38), .A1(n525), .B0(n22), .B1(n524), .Y(n375) );
  OAI22XL U358 ( .A0(n38), .A1(n526), .B0(n22), .B1(n525), .Y(n376) );
  OAI22XL U359 ( .A0(n38), .A1(n527), .B0(n22), .B1(n526), .Y(n377) );
  OAI22XL U360 ( .A0(n38), .A1(n528), .B0(n22), .B1(n527), .Y(n378) );
  OAI22XL U361 ( .A0(n38), .A1(n529), .B0(n22), .B1(n528), .Y(n379) );
  OAI22XL U362 ( .A0(n37), .A1(n530), .B0(n21), .B1(n529), .Y(n380) );
  OAI22XL U363 ( .A0(n37), .A1(n531), .B0(n21), .B1(n530), .Y(n381) );
  OAI22XL U364 ( .A0(n37), .A1(n532), .B0(n21), .B1(n531), .Y(n382) );
  OAI22XL U365 ( .A0(n37), .A1(n533), .B0(n21), .B1(n532), .Y(n383) );
  OAI22XL U366 ( .A0(n37), .A1(n534), .B0(n21), .B1(n533), .Y(n384) );
  OAI22XL U367 ( .A0(n37), .A1(n535), .B0(n21), .B1(n534), .Y(n385) );
  OAI22XL U368 ( .A0(n37), .A1(n536), .B0(n21), .B1(n535), .Y(n386) );
  OAI22XL U369 ( .A0(n37), .A1(n537), .B0(n21), .B1(n536), .Y(n387) );
  OAI22XL U370 ( .A0(n37), .A1(n538), .B0(n21), .B1(n537), .Y(n388) );
  NOR2BX1 U371 ( .AN(n49), .B(n21), .Y(n389) );
  XNOR2X1 U372 ( .A(n5), .B(n578), .Y(n521) );
  XNOR2X1 U373 ( .A(n5), .B(n579), .Y(n522) );
  XNOR2X1 U374 ( .A(n5), .B(n580), .Y(n523) );
  XNOR2X1 U375 ( .A(n5), .B(n581), .Y(n524) );
  XNOR2X1 U376 ( .A(n5), .B(n582), .Y(n525) );
  XNOR2X1 U377 ( .A(n5), .B(n583), .Y(n526) );
  XNOR2X1 U378 ( .A(n5), .B(n584), .Y(n527) );
  XNOR2X1 U379 ( .A(n5), .B(n585), .Y(n528) );
  XNOR2X1 U380 ( .A(n5), .B(n586), .Y(n529) );
  XNOR2X1 U381 ( .A(n5), .B(n587), .Y(n530) );
  XNOR2X1 U382 ( .A(n5), .B(n588), .Y(n531) );
  XNOR2X1 U383 ( .A(n5), .B(n589), .Y(n532) );
  XNOR2X1 U384 ( .A(n5), .B(n590), .Y(n533) );
  XNOR2X1 U385 ( .A(n5), .B(n591), .Y(n534) );
  XNOR2X1 U386 ( .A(n5), .B(n592), .Y(n535) );
  XNOR2X1 U387 ( .A(n5), .B(n593), .Y(n536) );
  XNOR2X1 U388 ( .A(n5), .B(n594), .Y(n537) );
  XNOR2X1 U389 ( .A(n5), .B(n49), .Y(n538) );
  NAND2BX1 U390 ( .AN(n49), .B(n5), .Y(n539) );
  OAI22XL U391 ( .A0(n36), .A1(n626), .B0(n20), .B1(n558), .Y(n280) );
  AO21X1 U392 ( .A0(n36), .A1(n20), .B0(n540), .Y(n390) );
  OAI22XL U393 ( .A0(n36), .A1(n541), .B0(n20), .B1(n540), .Y(n159) );
  OAI22XL U394 ( .A0(n36), .A1(n542), .B0(n20), .B1(n541), .Y(n391) );
  OAI22XL U395 ( .A0(n36), .A1(n543), .B0(n20), .B1(n542), .Y(n392) );
  OAI22XL U396 ( .A0(n36), .A1(n544), .B0(n20), .B1(n543), .Y(n393) );
  OAI22XL U397 ( .A0(n36), .A1(n545), .B0(n20), .B1(n544), .Y(n394) );
  OAI22XL U398 ( .A0(n36), .A1(n546), .B0(n20), .B1(n545), .Y(n395) );
  OAI22XL U399 ( .A0(n36), .A1(n547), .B0(n20), .B1(n546), .Y(n396) );
  OAI22XL U400 ( .A0(n36), .A1(n548), .B0(n20), .B1(n547), .Y(n397) );
  OAI22XL U401 ( .A0(n35), .A1(n549), .B0(n19), .B1(n548), .Y(n398) );
  OAI22XL U402 ( .A0(n35), .A1(n550), .B0(n19), .B1(n549), .Y(n399) );
  OAI22XL U403 ( .A0(n35), .A1(n551), .B0(n19), .B1(n550), .Y(n400) );
  OAI22XL U404 ( .A0(n35), .A1(n552), .B0(n19), .B1(n551), .Y(n401) );
  OAI22XL U405 ( .A0(n35), .A1(n553), .B0(n19), .B1(n552), .Y(n402) );
  OAI22XL U406 ( .A0(n35), .A1(n554), .B0(n19), .B1(n553), .Y(n403) );
  OAI22XL U407 ( .A0(n35), .A1(n555), .B0(n19), .B1(n554), .Y(n404) );
  OAI22XL U408 ( .A0(n35), .A1(n556), .B0(n19), .B1(n555), .Y(n405) );
  OAI22XL U409 ( .A0(n35), .A1(n557), .B0(n19), .B1(n556), .Y(n406) );
  NOR2BX1 U410 ( .AN(n49), .B(n19), .Y(n407) );
  XNOR2X1 U411 ( .A(n3), .B(n578), .Y(n540) );
  XNOR2X1 U412 ( .A(n3), .B(n579), .Y(n541) );
  XNOR2X1 U413 ( .A(n3), .B(n580), .Y(n542) );
  XNOR2X1 U414 ( .A(n3), .B(n581), .Y(n543) );
  XNOR2X1 U415 ( .A(n3), .B(n582), .Y(n544) );
  XNOR2X1 U416 ( .A(n3), .B(n583), .Y(n545) );
  XNOR2X1 U417 ( .A(n3), .B(n584), .Y(n546) );
  XNOR2X1 U418 ( .A(n3), .B(n585), .Y(n547) );
  XNOR2X1 U419 ( .A(n3), .B(n586), .Y(n548) );
  XNOR2X1 U420 ( .A(n3), .B(n587), .Y(n549) );
  XNOR2X1 U421 ( .A(n3), .B(n588), .Y(n550) );
  XNOR2X1 U422 ( .A(n3), .B(n589), .Y(n551) );
  XNOR2X1 U423 ( .A(n3), .B(n590), .Y(n552) );
  XNOR2X1 U424 ( .A(n3), .B(n591), .Y(n553) );
  XNOR2X1 U425 ( .A(n3), .B(n592), .Y(n554) );
  XNOR2X1 U426 ( .A(n3), .B(n593), .Y(n555) );
  XNOR2X1 U427 ( .A(n3), .B(n594), .Y(n556) );
  XNOR2X1 U428 ( .A(n3), .B(n49), .Y(n557) );
  NAND2BX1 U429 ( .AN(n49), .B(n3), .Y(n558) );
  OAI22XL U430 ( .A0(n34), .A1(n627), .B0(n577), .B1(n18), .Y(n281) );
  AO21X1 U431 ( .A0(n34), .A1(n18), .B0(n559), .Y(n408) );
  OAI22XL U432 ( .A0(n34), .A1(n560), .B0(n559), .B1(n18), .Y(n409) );
  OAI22XL U433 ( .A0(n34), .A1(n561), .B0(n560), .B1(n18), .Y(n410) );
  OAI22XL U434 ( .A0(n34), .A1(n562), .B0(n561), .B1(n18), .Y(n411) );
  OAI22XL U435 ( .A0(n34), .A1(n563), .B0(n562), .B1(n18), .Y(n412) );
  OAI22XL U436 ( .A0(n34), .A1(n564), .B0(n563), .B1(n18), .Y(n413) );
  OAI22XL U437 ( .A0(n34), .A1(n565), .B0(n564), .B1(n18), .Y(n414) );
  OAI22XL U438 ( .A0(n34), .A1(n566), .B0(n565), .B1(n18), .Y(n415) );
  OAI22XL U439 ( .A0(n34), .A1(n567), .B0(n566), .B1(n18), .Y(n416) );
  OAI22XL U440 ( .A0(n33), .A1(n568), .B0(n567), .B1(n17), .Y(n417) );
  OAI22XL U441 ( .A0(n33), .A1(n569), .B0(n568), .B1(n17), .Y(n418) );
  OAI22XL U442 ( .A0(n33), .A1(n570), .B0(n569), .B1(n17), .Y(n419) );
  OAI22XL U443 ( .A0(n33), .A1(n571), .B0(n570), .B1(n17), .Y(n420) );
  OAI22XL U444 ( .A0(n33), .A1(n572), .B0(n571), .B1(n17), .Y(n421) );
  OAI22XL U445 ( .A0(n33), .A1(n573), .B0(n572), .B1(n17), .Y(n422) );
  OAI22XL U446 ( .A0(n33), .A1(n574), .B0(n573), .B1(n17), .Y(n423) );
  OAI22XL U447 ( .A0(n33), .A1(n575), .B0(n574), .B1(n17), .Y(n424) );
  OAI22XL U448 ( .A0(n33), .A1(n576), .B0(n575), .B1(n17), .Y(n425) );
  NOR2BX1 U449 ( .AN(n49), .B(n17), .Y(product_0_) );
  XNOR2X1 U450 ( .A(n1), .B(n578), .Y(n559) );
  XNOR2X1 U451 ( .A(n1), .B(n579), .Y(n560) );
  XNOR2X1 U452 ( .A(n1), .B(n580), .Y(n561) );
  XNOR2X1 U453 ( .A(n1), .B(n581), .Y(n562) );
  XNOR2X1 U454 ( .A(n1), .B(n582), .Y(n563) );
  XNOR2X1 U455 ( .A(n1), .B(n583), .Y(n564) );
  XNOR2X1 U456 ( .A(n1), .B(n584), .Y(n565) );
  XNOR2X1 U457 ( .A(n1), .B(n585), .Y(n566) );
  XNOR2X1 U458 ( .A(n1), .B(n586), .Y(n567) );
  XNOR2X1 U459 ( .A(n1), .B(n587), .Y(n568) );
  XNOR2X1 U460 ( .A(n1), .B(n588), .Y(n569) );
  XNOR2X1 U461 ( .A(n1), .B(n589), .Y(n570) );
  XNOR2X1 U462 ( .A(n1), .B(n590), .Y(n571) );
  XNOR2X1 U463 ( .A(n1), .B(n591), .Y(n572) );
  XNOR2X1 U464 ( .A(n1), .B(n592), .Y(n573) );
  XNOR2X1 U465 ( .A(n1), .B(n593), .Y(n574) );
  XNOR2X1 U466 ( .A(n1), .B(n594), .Y(n575) );
  XNOR2X1 U467 ( .A(n1), .B(n49), .Y(n576) );
  NAND2BX1 U468 ( .AN(n49), .B(n1), .Y(n577) );
  CLKINVX1 U486 ( .A(n15), .Y(n620) );
  CLKINVX1 U487 ( .A(n13), .Y(n621) );
  CLKINVX1 U488 ( .A(n11), .Y(n622) );
  CLKINVX1 U489 ( .A(n9), .Y(n623) );
  CLKINVX1 U490 ( .A(n7), .Y(n624) );
  CLKINVX1 U491 ( .A(n5), .Y(n625) );
  CLKINVX1 U492 ( .A(n3), .Y(n626) );
  CLKINVX1 U493 ( .A(n1), .Y(n627) );
  NAND2X1 U494 ( .A(n596), .B(n612), .Y(n604) );
  XOR2X1 U495 ( .A(a[14]), .B(a[15]), .Y(n596) );
  XNOR2X1 U496 ( .A(a[14]), .B(a[13]), .Y(n612) );
  NAND2X1 U497 ( .A(n597), .B(n613), .Y(n605) );
  XOR2X1 U498 ( .A(a[12]), .B(a[13]), .Y(n597) );
  XNOR2X1 U499 ( .A(a[12]), .B(a[11]), .Y(n613) );
  NAND2X1 U500 ( .A(n598), .B(n614), .Y(n606) );
  XOR2X1 U501 ( .A(a[10]), .B(a[11]), .Y(n598) );
  XNOR2X1 U502 ( .A(a[10]), .B(a[9]), .Y(n614) );
  NAND2X1 U503 ( .A(n599), .B(n615), .Y(n607) );
  XOR2X1 U504 ( .A(a[8]), .B(a[9]), .Y(n599) );
  XNOR2X1 U505 ( .A(a[8]), .B(a[7]), .Y(n615) );
  NAND2X1 U506 ( .A(n600), .B(n616), .Y(n608) );
  XOR2X1 U507 ( .A(a[6]), .B(a[7]), .Y(n600) );
  XNOR2X1 U508 ( .A(a[6]), .B(a[5]), .Y(n616) );
  NAND2X1 U509 ( .A(n601), .B(n617), .Y(n609) );
  XOR2X1 U510 ( .A(a[4]), .B(a[5]), .Y(n601) );
  XNOR2X1 U511 ( .A(a[4]), .B(a[3]), .Y(n617) );
  NAND2X1 U512 ( .A(n602), .B(n618), .Y(n610) );
  XOR2X1 U513 ( .A(a[2]), .B(a[3]), .Y(n602) );
  XNOR2X1 U514 ( .A(a[2]), .B(a[1]), .Y(n618) );
  NAND2X1 U515 ( .A(n603), .B(n619), .Y(n611) );
  XOR2X1 U516 ( .A(a[0]), .B(a[1]), .Y(n603) );
  CLKINVX1 U517 ( .A(a[0]), .Y(n619) );
  OA22X1 U520 ( .A0(n48), .A1(n427), .B0(n32), .B1(n426), .Y(n697) );
  CLKBUFX3 U521 ( .A(b_2_), .Y(n593) );
  CLKBUFX3 U522 ( .A(b_0_), .Y(n49) );
  CLKBUFX3 U523 ( .A(b_3_), .Y(n592) );
  CLKBUFX3 U524 ( .A(b_9_), .Y(n586) );
  CLKBUFX3 U525 ( .A(b_17_), .Y(n578) );
  CLKBUFX3 U526 ( .A(b_4_), .Y(n591) );
  CLKBUFX3 U527 ( .A(b_5_), .Y(n590) );
  CLKBUFX3 U528 ( .A(b_6_), .Y(n589) );
  CLKBUFX3 U529 ( .A(b_10_), .Y(n585) );
  CLKBUFX3 U530 ( .A(b_15_), .Y(n580) );
  CLKBUFX3 U531 ( .A(b_7_), .Y(n588) );
  CLKBUFX3 U532 ( .A(b_14_), .Y(n581) );
  CLKBUFX3 U533 ( .A(b_1_), .Y(n594) );
  CLKBUFX3 U534 ( .A(b_16_), .Y(n579) );
  CLKBUFX3 U535 ( .A(n618), .Y(n19) );
  CLKBUFX3 U536 ( .A(n617), .Y(n21) );
  CLKBUFX3 U537 ( .A(n616), .Y(n23) );
  CLKBUFX3 U538 ( .A(n615), .Y(n25) );
  CLKBUFX3 U539 ( .A(n614), .Y(n27) );
  CLKBUFX3 U540 ( .A(n613), .Y(n29) );
  CLKBUFX3 U541 ( .A(n612), .Y(n31) );
  CLKBUFX3 U542 ( .A(n618), .Y(n20) );
  CLKBUFX3 U543 ( .A(n617), .Y(n22) );
  CLKBUFX3 U544 ( .A(n615), .Y(n26) );
  CLKBUFX3 U545 ( .A(n616), .Y(n24) );
  CLKBUFX3 U546 ( .A(n613), .Y(n30) );
  CLKBUFX3 U547 ( .A(n614), .Y(n28) );
  CLKBUFX3 U548 ( .A(b_13_), .Y(n582) );
  CLKBUFX3 U549 ( .A(b_8_), .Y(n587) );
  CLKBUFX3 U550 ( .A(n612), .Y(n32) );
  CLKBUFX3 U551 ( .A(b_11_), .Y(n584) );
  CLKBUFX3 U552 ( .A(b_12_), .Y(n583) );
  CLKBUFX3 U553 ( .A(n610), .Y(n36) );
  CLKBUFX3 U554 ( .A(n609), .Y(n38) );
  CLKBUFX3 U555 ( .A(n607), .Y(n42) );
  CLKBUFX3 U556 ( .A(n608), .Y(n40) );
  CLKBUFX3 U557 ( .A(n605), .Y(n46) );
  CLKBUFX3 U558 ( .A(n606), .Y(n44) );
  CLKBUFX3 U559 ( .A(n611), .Y(n34) );
  CLKBUFX3 U560 ( .A(n610), .Y(n35) );
  CLKBUFX3 U561 ( .A(n609), .Y(n37) );
  CLKBUFX3 U562 ( .A(n608), .Y(n39) );
  CLKBUFX3 U563 ( .A(n607), .Y(n41) );
  CLKBUFX3 U564 ( .A(n606), .Y(n43) );
  CLKBUFX3 U565 ( .A(n605), .Y(n45) );
  CLKBUFX3 U566 ( .A(n604), .Y(n47) );
  CLKBUFX3 U567 ( .A(n604), .Y(n48) );
  CLKBUFX3 U568 ( .A(n611), .Y(n33) );
  CLKBUFX3 U569 ( .A(n619), .Y(n17) );
  CLKBUFX3 U570 ( .A(n619), .Y(n18) );
  CLKBUFX3 U571 ( .A(a[1]), .Y(n1) );
  CLKBUFX3 U572 ( .A(a[3]), .Y(n3) );
  CLKBUFX3 U573 ( .A(a[5]), .Y(n5) );
  CLKBUFX3 U574 ( .A(a[7]), .Y(n7) );
  CLKBUFX3 U575 ( .A(a[9]), .Y(n9) );
  CLKBUFX3 U576 ( .A(a[11]), .Y(n11) );
  CLKBUFX3 U577 ( .A(a[13]), .Y(n13) );
  CLKBUFX3 U578 ( .A(a[15]), .Y(n15) );
endmodule


module FAS_DW_mult_tc_26 ( a, b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, 
        b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input [15:0] a;
  input b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_, b_8_, b_7_,
         b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n3, n5, n7, n9, n11, n13, n15, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600;

  XOR2X1 U51 ( .A(n52), .B(n51), .Y(product_31_) );
  XOR2X1 U52 ( .A(n272), .B(n82), .Y(n51) );
  ADDFXL U53 ( .A(n84), .B(n83), .CI(n53), .CO(n52), .S(product_30_) );
  ADDFXL U54 ( .A(n85), .B(n86), .CI(n54), .CO(n53), .S(product_29_) );
  ADDFXL U55 ( .A(n91), .B(n87), .CI(n55), .CO(n54), .S(product_28_) );
  ADDFXL U56 ( .A(n94), .B(n92), .CI(n56), .CO(n55), .S(product_27_) );
  ADDFXL U57 ( .A(n95), .B(n99), .CI(n57), .CO(n56), .S(product_26_) );
  ADDFXL U58 ( .A(n100), .B(n104), .CI(n58), .CO(n57), .S(product_25_) );
  ADDFXL U59 ( .A(n105), .B(n111), .CI(n59), .CO(n58), .S(product_24_) );
  ADDFXL U60 ( .A(n112), .B(n117), .CI(n60), .CO(n59), .S(product_23_) );
  ADDFXL U61 ( .A(n118), .B(n125), .CI(n61), .CO(n60), .S(product_22_) );
  ADDFXL U62 ( .A(n133), .B(n126), .CI(n62), .CO(n61), .S(product_21_) );
  ADDFXL U63 ( .A(n143), .B(n134), .CI(n63), .CO(n62), .S(product_20_) );
  ADDFXL U64 ( .A(n144), .B(n152), .CI(n64), .CO(n63), .S(product_19_) );
  ADDFXL U65 ( .A(n153), .B(n163), .CI(n65), .CO(n64), .S(product_18_) );
  ADDFXL U66 ( .A(n164), .B(n174), .CI(n66), .CO(n65), .S(product_17_) );
  ADDFXL U67 ( .A(n175), .B(n185), .CI(n67), .CO(n66), .S(product_16_) );
  ADDFXL U68 ( .A(n186), .B(n196), .CI(n68), .CO(n67), .S(product_15_) );
  ADDFXL U69 ( .A(n197), .B(n205), .CI(n69), .CO(n68), .S(product_14_) );
  ADDFXL U70 ( .A(n206), .B(n215), .CI(n70), .CO(n69), .S(product_13_) );
  ADDFXL U71 ( .A(n216), .B(n223), .CI(n71), .CO(n70), .S(product_12_) );
  ADDFXL U72 ( .A(n224), .B(n231), .CI(n72), .CO(n71), .S(product_11_) );
  ADDFXL U73 ( .A(n232), .B(n237), .CI(n73), .CO(n72), .S(product_10_) );
  ADDFXL U74 ( .A(n238), .B(n244), .CI(n74), .CO(n73), .S(product_9_) );
  ADDFXL U75 ( .A(n245), .B(n249), .CI(n75), .CO(n74), .S(product_8_) );
  ADDFXL U76 ( .A(n250), .B(n254), .CI(n76), .CO(n75), .S(product_7_) );
  ADDFXL U77 ( .A(n255), .B(n256), .CI(n77), .CO(n76), .S(product_6_) );
  ADDFXL U78 ( .A(n257), .B(n260), .CI(n78), .CO(n77), .S(product_5_) );
  ADDFXL U79 ( .A(n261), .B(n262), .CI(n79), .CO(n78), .S(product_4_) );
  ADDFXL U80 ( .A(n263), .B(n389), .CI(n80), .CO(n79), .S(product_3_) );
  ADDFXL U81 ( .A(n406), .B(n390), .CI(n81), .CO(n80), .S(product_2_) );
  ADDHXL U82 ( .A(n271), .B(n407), .CO(n81), .S(product_1_) );
  CLKINVX1 U83 ( .A(n82), .Y(n83) );
  ADDFXL U84 ( .A(n273), .B(n88), .CI(n289), .CO(n84), .S(n85) );
  ADDFXL U85 ( .A(n89), .B(n274), .CI(n90), .CO(n86), .S(n87) );
  CLKINVX1 U86 ( .A(n88), .Y(n89) );
  CMPR42X1 U87 ( .A(n96), .B(n275), .C(n290), .D(n306), .ICI(n93), .S(n92), 
        .ICO(n90), .CO(n91) );
  CMPR42X1 U88 ( .A(n291), .B(n276), .C(n97), .D(n101), .ICI(n98), .S(n95), 
        .ICO(n93), .CO(n94) );
  CLKINVX1 U89 ( .A(n96), .Y(n97) );
  CMPR42X1 U90 ( .A(n307), .B(n292), .C(n106), .D(n102), .ICI(n103), .S(n100), 
        .ICO(n98), .CO(n99) );
  ADDFXL U91 ( .A(n108), .B(n277), .CI(n322), .CO(n101), .S(n102) );
  CMPR42X1 U92 ( .A(n308), .B(n113), .C(n107), .D(n114), .ICI(n110), .S(n105), 
        .ICO(n103), .CO(n104) );
  ADDFXL U93 ( .A(n293), .B(n278), .CI(n109), .CO(n106), .S(n107) );
  CLKINVX1 U94 ( .A(n108), .Y(n109) );
  CMPR42X1 U95 ( .A(n309), .B(n294), .C(n120), .D(n115), .ICI(n116), .S(n112), 
        .ICO(n110), .CO(n111) );
  CMPR42X1 U96 ( .A(n279), .B(n122), .C(n323), .D(n339), .ICI(n119), .S(n115), 
        .ICO(n113), .CO(n114) );
  CMPR42X1 U97 ( .A(n280), .B(n130), .C(n128), .D(n121), .ICI(n124), .S(n118), 
        .ICO(n116), .CO(n117) );
  CMPR42X1 U98 ( .A(n295), .B(n340), .C(n324), .D(n123), .ICI(n127), .S(n121), 
        .ICO(n119), .CO(n120) );
  CLKINVX1 U99 ( .A(n122), .Y(n123) );
  CMPR42X1 U100 ( .A(n138), .B(n131), .C(n136), .D(n129), .ICI(n132), .S(n126), 
        .ICO(n124), .CO(n125) );
  CMPR42X1 U101 ( .A(n296), .B(n325), .C(n310), .D(n140), .ICI(n135), .S(n129), 
        .ICO(n127), .CO(n128) );
  ADDFXL U102 ( .A(n341), .B(n281), .CI(n357), .CO(n130), .S(n131) );
  CMPR42X1 U103 ( .A(n139), .B(n149), .C(n146), .D(n137), .ICI(n142), .S(n134), 
        .ICO(n132), .CO(n133) );
  CMPR42X1 U104 ( .A(n342), .B(n311), .C(n326), .D(n145), .ICI(n148), .S(n137), 
        .ICO(n135), .CO(n136) );
  ADDFXL U105 ( .A(n282), .B(n297), .CI(n141), .CO(n138), .S(n139) );
  CLKINVX1 U106 ( .A(n140), .Y(n141) );
  CMPR42X1 U107 ( .A(n158), .B(n155), .C(n147), .D(n150), .ICI(n151), .S(n144), 
        .ICO(n142), .CO(n143) );
  CMPR42X1 U108 ( .A(n298), .B(n327), .C(n312), .D(n160), .ICI(n154), .S(n147), 
        .ICO(n145), .CO(n146) );
  CMPR42X1 U109 ( .A(n283), .B(n358), .C(n343), .D(n374), .ICI(n157), .S(n150), 
        .ICO(n148), .CO(n149) );
  CMPR42X1 U110 ( .A(n169), .B(n166), .C(n156), .D(n159), .ICI(n162), .S(n153), 
        .ICO(n151), .CO(n152) );
  CMPR42X1 U111 ( .A(n313), .B(n344), .C(n328), .D(n284), .ICI(n165), .S(n156), 
        .ICO(n154), .CO(n155) );
  CMPR42X1 U112 ( .A(n299), .B(n359), .C(n161), .D(n171), .ICI(n168), .S(n159), 
        .ICO(n157), .CO(n158) );
  CLKINVX1 U113 ( .A(n160), .Y(n161) );
  CMPR42X1 U114 ( .A(n180), .B(n177), .C(n167), .D(n170), .ICI(n173), .S(n164), 
        .ICO(n162), .CO(n163) );
  CMPR42X1 U115 ( .A(n285), .B(n360), .C(n329), .D(n182), .ICI(n176), .S(n167), 
        .ICO(n165), .CO(n166) );
  CMPR42X1 U116 ( .A(n314), .B(n375), .C(n391), .D(n172), .ICI(n179), .S(n170), 
        .ICO(n168), .CO(n169) );
  XNOR2X1 U117 ( .A(n345), .B(n300), .Y(n172) );
  OR2X1 U118 ( .A(n345), .B(n300), .Y(n171) );
  CMPR42X1 U119 ( .A(n191), .B(n188), .C(n181), .D(n178), .ICI(n184), .S(n175), 
        .ICO(n173), .CO(n174) );
  CMPR42X1 U120 ( .A(n301), .B(n315), .C(n346), .D(n183), .ICI(n190), .S(n178), 
        .ICO(n176), .CO(n177) );
  CMPR42X1 U121 ( .A(n330), .B(n376), .C(n361), .D(n193), .ICI(n187), .S(n181), 
        .ICO(n179), .CO(n180) );
  ADDHXL U122 ( .A(n392), .B(n286), .CO(n182), .S(n183) );
  CMPR42X1 U123 ( .A(n202), .B(n199), .C(n192), .D(n189), .ICI(n195), .S(n186), 
        .ICO(n184), .CO(n185) );
  CMPR42X1 U124 ( .A(n302), .B(n316), .C(n331), .D(n201), .ICI(n194), .S(n189), 
        .ICO(n187), .CO(n188) );
  CMPR42X1 U125 ( .A(n264), .B(n287), .C(n377), .D(n347), .ICI(n198), .S(n192), 
        .ICO(n190), .CO(n191) );
  ADDHXL U126 ( .A(n393), .B(n362), .CO(n193), .S(n194) );
  CMPR42X1 U127 ( .A(n210), .B(n203), .C(n208), .D(n200), .ICI(n204), .S(n197), 
        .ICO(n195), .CO(n196) );
  CMPR42X1 U128 ( .A(n378), .B(n332), .C(n348), .D(n363), .ICI(n212), .S(n200), 
        .ICO(n198), .CO(n199) );
  CMPR42X1 U129 ( .A(n288), .B(n394), .C(n303), .D(n317), .ICI(n207), .S(n203), 
        .ICO(n201), .CO(n202) );
  CMPR42X1 U130 ( .A(n220), .B(n211), .C(n218), .D(n209), .ICI(n214), .S(n206), 
        .ICO(n204), .CO(n205) );
  CMPR42X1 U131 ( .A(n318), .B(n349), .C(n333), .D(n304), .ICI(n217), .S(n209), 
        .ICO(n207), .CO(n208) );
  ADDFXL U132 ( .A(n379), .B(n265), .CI(n213), .CO(n210), .S(n211) );
  ADDHXL U133 ( .A(n395), .B(n364), .CO(n212), .S(n213) );
  CMPR42X1 U134 ( .A(n350), .B(n225), .C(n226), .D(n219), .ICI(n222), .S(n216), 
        .ICO(n214), .CO(n215) );
  CMPR42X1 U135 ( .A(n380), .B(n334), .C(n365), .D(n228), .ICI(n221), .S(n219), 
        .ICO(n217), .CO(n218) );
  ADDFXL U136 ( .A(n396), .B(n305), .CI(n319), .CO(n220), .S(n221) );
  CMPR42X1 U137 ( .A(n351), .B(n233), .C(n234), .D(n227), .ICI(n230), .S(n224), 
        .ICO(n222), .CO(n223) );
  CMPR42X1 U138 ( .A(n266), .B(n320), .C(n381), .D(n335), .ICI(n229), .S(n227), 
        .ICO(n225), .CO(n226) );
  ADDHXL U139 ( .A(n397), .B(n366), .CO(n228), .S(n229) );
  CMPR42X1 U140 ( .A(n382), .B(n367), .C(n239), .D(n236), .ICI(n235), .S(n232), 
        .ICO(n230), .CO(n231) );
  CMPR42X1 U141 ( .A(n321), .B(n398), .C(n336), .D(n352), .ICI(n241), .S(n235), 
        .ICO(n233), .CO(n234) );
  CMPR42X1 U142 ( .A(n383), .B(n353), .C(n243), .D(n246), .ICI(n240), .S(n238), 
        .ICO(n236), .CO(n237) );
  ADDFXL U143 ( .A(n337), .B(n267), .CI(n242), .CO(n239), .S(n240) );
  ADDHXL U144 ( .A(n399), .B(n368), .CO(n241), .S(n242) );
  CMPR42X1 U145 ( .A(n384), .B(n369), .C(n251), .D(n248), .ICI(n247), .S(n245), 
        .ICO(n243), .CO(n244) );
  ADDFXL U146 ( .A(n400), .B(n338), .CI(n354), .CO(n246), .S(n247) );
  CMPR42X1 U147 ( .A(n268), .B(n355), .C(n385), .D(n253), .ICI(n252), .S(n250), 
        .ICO(n248), .CO(n249) );
  ADDHXL U148 ( .A(n401), .B(n370), .CO(n251), .S(n252) );
  CMPR42X1 U149 ( .A(n356), .B(n402), .C(n371), .D(n386), .ICI(n258), .S(n255), 
        .ICO(n253), .CO(n254) );
  ADDFXL U150 ( .A(n387), .B(n269), .CI(n259), .CO(n256), .S(n257) );
  ADDHXL U151 ( .A(n403), .B(n372), .CO(n258), .S(n259) );
  ADDFXL U152 ( .A(n404), .B(n373), .CI(n388), .CO(n260), .S(n261) );
  ADDHXL U153 ( .A(n405), .B(n270), .CO(n262), .S(n263) );
  OAI22XL U154 ( .A0(n48), .A1(n593), .B0(n32), .B1(n425), .Y(n264) );
  AO21X1 U155 ( .A0(n48), .A1(n32), .B0(n408), .Y(n272) );
  OAI22XL U156 ( .A0(n48), .A1(n409), .B0(n32), .B1(n408), .Y(n82) );
  OAI22XL U157 ( .A0(n48), .A1(n410), .B0(n32), .B1(n409), .Y(n273) );
  OAI22XL U158 ( .A0(n48), .A1(n411), .B0(n32), .B1(n410), .Y(n274) );
  OAI22XL U159 ( .A0(n48), .A1(n412), .B0(n32), .B1(n411), .Y(n275) );
  OAI22XL U160 ( .A0(n48), .A1(n413), .B0(n32), .B1(n412), .Y(n276) );
  OAI22XL U161 ( .A0(n48), .A1(n414), .B0(n32), .B1(n413), .Y(n277) );
  OAI22XL U162 ( .A0(n48), .A1(n415), .B0(n32), .B1(n414), .Y(n278) );
  OAI22XL U163 ( .A0(n47), .A1(n416), .B0(n32), .B1(n415), .Y(n279) );
  OAI22XL U164 ( .A0(n47), .A1(n417), .B0(n31), .B1(n416), .Y(n280) );
  OAI22XL U165 ( .A0(n47), .A1(n418), .B0(n31), .B1(n417), .Y(n281) );
  OAI22XL U166 ( .A0(n47), .A1(n419), .B0(n31), .B1(n418), .Y(n282) );
  OAI22XL U167 ( .A0(n47), .A1(n420), .B0(n31), .B1(n419), .Y(n283) );
  OAI22XL U168 ( .A0(n47), .A1(n421), .B0(n31), .B1(n420), .Y(n284) );
  OAI22XL U169 ( .A0(n47), .A1(n422), .B0(n31), .B1(n421), .Y(n285) );
  OAI22XL U170 ( .A0(n47), .A1(n423), .B0(n31), .B1(n422), .Y(n286) );
  OAI22XL U171 ( .A0(n47), .A1(n424), .B0(n31), .B1(n423), .Y(n287) );
  NOR2BX1 U172 ( .AN(n49), .B(n31), .Y(n288) );
  XNOR2X1 U173 ( .A(n15), .B(n552), .Y(n408) );
  XNOR2X1 U174 ( .A(n15), .B(n553), .Y(n409) );
  XNOR2X1 U175 ( .A(n15), .B(n554), .Y(n410) );
  XNOR2X1 U176 ( .A(n15), .B(n555), .Y(n411) );
  XNOR2X1 U177 ( .A(n15), .B(n556), .Y(n412) );
  XNOR2X1 U178 ( .A(n15), .B(n557), .Y(n413) );
  XNOR2X1 U179 ( .A(n15), .B(n558), .Y(n414) );
  XNOR2X1 U180 ( .A(n15), .B(n559), .Y(n415) );
  XNOR2X1 U181 ( .A(n15), .B(n560), .Y(n416) );
  XNOR2X1 U182 ( .A(n15), .B(n561), .Y(n417) );
  XNOR2X1 U183 ( .A(n15), .B(n562), .Y(n418) );
  XNOR2X1 U184 ( .A(n15), .B(n563), .Y(n419) );
  XNOR2X1 U185 ( .A(n15), .B(n564), .Y(n420) );
  XNOR2X1 U186 ( .A(n15), .B(n565), .Y(n421) );
  XNOR2X1 U187 ( .A(n15), .B(n566), .Y(n422) );
  XNOR2X1 U188 ( .A(n15), .B(n567), .Y(n423) );
  XNOR2X1 U189 ( .A(n15), .B(n49), .Y(n424) );
  NAND2BX1 U190 ( .AN(n49), .B(n15), .Y(n425) );
  OAI22XL U191 ( .A0(n46), .A1(n594), .B0(n30), .B1(n443), .Y(n265) );
  AO21X1 U192 ( .A0(n46), .A1(n30), .B0(n426), .Y(n289) );
  OAI22XL U193 ( .A0(n46), .A1(n427), .B0(n30), .B1(n426), .Y(n88) );
  OAI22XL U194 ( .A0(n46), .A1(n428), .B0(n30), .B1(n427), .Y(n290) );
  OAI22XL U195 ( .A0(n46), .A1(n429), .B0(n30), .B1(n428), .Y(n291) );
  OAI22XL U196 ( .A0(n46), .A1(n430), .B0(n30), .B1(n429), .Y(n292) );
  OAI22XL U197 ( .A0(n46), .A1(n431), .B0(n30), .B1(n430), .Y(n293) );
  OAI22XL U198 ( .A0(n46), .A1(n432), .B0(n30), .B1(n431), .Y(n294) );
  OAI22XL U199 ( .A0(n46), .A1(n433), .B0(n30), .B1(n432), .Y(n295) );
  OAI22XL U200 ( .A0(n45), .A1(n434), .B0(n30), .B1(n433), .Y(n296) );
  OAI22XL U201 ( .A0(n45), .A1(n435), .B0(n29), .B1(n434), .Y(n297) );
  OAI22XL U202 ( .A0(n45), .A1(n436), .B0(n29), .B1(n435), .Y(n298) );
  OAI22XL U203 ( .A0(n45), .A1(n437), .B0(n29), .B1(n436), .Y(n299) );
  OAI22XL U204 ( .A0(n45), .A1(n438), .B0(n29), .B1(n437), .Y(n300) );
  OAI22XL U205 ( .A0(n45), .A1(n439), .B0(n29), .B1(n438), .Y(n301) );
  OAI22XL U206 ( .A0(n45), .A1(n440), .B0(n29), .B1(n439), .Y(n302) );
  OAI22XL U207 ( .A0(n45), .A1(n441), .B0(n29), .B1(n440), .Y(n303) );
  OAI22XL U208 ( .A0(n45), .A1(n442), .B0(n29), .B1(n441), .Y(n304) );
  NOR2BX1 U209 ( .AN(n49), .B(n29), .Y(n305) );
  XNOR2X1 U210 ( .A(n13), .B(n552), .Y(n426) );
  XNOR2X1 U211 ( .A(n13), .B(n553), .Y(n427) );
  XNOR2X1 U212 ( .A(n13), .B(n554), .Y(n428) );
  XNOR2X1 U213 ( .A(n13), .B(n555), .Y(n429) );
  XNOR2X1 U214 ( .A(n13), .B(n556), .Y(n430) );
  XNOR2X1 U215 ( .A(n13), .B(n557), .Y(n431) );
  XNOR2X1 U216 ( .A(n13), .B(n558), .Y(n432) );
  XNOR2X1 U217 ( .A(n13), .B(n559), .Y(n433) );
  XNOR2X1 U218 ( .A(n13), .B(n560), .Y(n434) );
  XNOR2X1 U219 ( .A(n13), .B(n561), .Y(n435) );
  XNOR2X1 U220 ( .A(n13), .B(n562), .Y(n436) );
  XNOR2X1 U221 ( .A(n13), .B(n563), .Y(n437) );
  XNOR2X1 U222 ( .A(n13), .B(n564), .Y(n438) );
  XNOR2X1 U223 ( .A(n13), .B(n565), .Y(n439) );
  XNOR2X1 U224 ( .A(n13), .B(n566), .Y(n440) );
  XNOR2X1 U225 ( .A(n13), .B(n567), .Y(n441) );
  XNOR2X1 U226 ( .A(n13), .B(n49), .Y(n442) );
  NAND2BX1 U227 ( .AN(n49), .B(n13), .Y(n443) );
  OAI22XL U228 ( .A0(n44), .A1(n595), .B0(n28), .B1(n461), .Y(n266) );
  AO21X1 U229 ( .A0(n44), .A1(n28), .B0(n444), .Y(n306) );
  OAI22XL U230 ( .A0(n44), .A1(n445), .B0(n28), .B1(n444), .Y(n96) );
  OAI22XL U231 ( .A0(n44), .A1(n446), .B0(n28), .B1(n445), .Y(n307) );
  OAI22XL U232 ( .A0(n44), .A1(n447), .B0(n28), .B1(n446), .Y(n308) );
  OAI22XL U233 ( .A0(n44), .A1(n448), .B0(n28), .B1(n447), .Y(n309) );
  OAI22XL U234 ( .A0(n44), .A1(n449), .B0(n28), .B1(n448), .Y(n122) );
  OAI22XL U235 ( .A0(n44), .A1(n450), .B0(n28), .B1(n449), .Y(n310) );
  OAI22XL U236 ( .A0(n44), .A1(n451), .B0(n28), .B1(n450), .Y(n311) );
  OAI22XL U237 ( .A0(n43), .A1(n452), .B0(n28), .B1(n451), .Y(n312) );
  OAI22XL U238 ( .A0(n43), .A1(n453), .B0(n27), .B1(n452), .Y(n313) );
  OAI22XL U239 ( .A0(n43), .A1(n454), .B0(n27), .B1(n453), .Y(n314) );
  OAI22XL U240 ( .A0(n43), .A1(n455), .B0(n27), .B1(n454), .Y(n315) );
  OAI22XL U241 ( .A0(n43), .A1(n456), .B0(n27), .B1(n455), .Y(n316) );
  OAI22XL U242 ( .A0(n43), .A1(n457), .B0(n27), .B1(n456), .Y(n317) );
  OAI22XL U243 ( .A0(n43), .A1(n458), .B0(n27), .B1(n457), .Y(n318) );
  OAI22XL U244 ( .A0(n43), .A1(n459), .B0(n27), .B1(n458), .Y(n319) );
  OAI22XL U245 ( .A0(n43), .A1(n460), .B0(n27), .B1(n459), .Y(n320) );
  NOR2BX1 U246 ( .AN(n49), .B(n27), .Y(n321) );
  XNOR2X1 U247 ( .A(n11), .B(n552), .Y(n444) );
  XNOR2X1 U248 ( .A(n11), .B(n553), .Y(n445) );
  XNOR2X1 U249 ( .A(n11), .B(n554), .Y(n446) );
  XNOR2X1 U250 ( .A(n11), .B(n555), .Y(n447) );
  XNOR2X1 U251 ( .A(n11), .B(n556), .Y(n448) );
  XNOR2X1 U252 ( .A(n11), .B(n557), .Y(n449) );
  XNOR2X1 U253 ( .A(n11), .B(n558), .Y(n450) );
  XNOR2X1 U254 ( .A(n11), .B(n559), .Y(n451) );
  XNOR2X1 U255 ( .A(n11), .B(n560), .Y(n452) );
  XNOR2X1 U256 ( .A(n11), .B(n561), .Y(n453) );
  XNOR2X1 U257 ( .A(n11), .B(n562), .Y(n454) );
  XNOR2X1 U258 ( .A(n11), .B(n563), .Y(n455) );
  XNOR2X1 U259 ( .A(n11), .B(n564), .Y(n456) );
  XNOR2X1 U260 ( .A(n11), .B(n565), .Y(n457) );
  XNOR2X1 U261 ( .A(n11), .B(n566), .Y(n458) );
  XNOR2X1 U262 ( .A(n11), .B(n567), .Y(n459) );
  XNOR2X1 U263 ( .A(n11), .B(n49), .Y(n460) );
  NAND2BX1 U264 ( .AN(n49), .B(n11), .Y(n461) );
  OAI22XL U265 ( .A0(n42), .A1(n596), .B0(n26), .B1(n479), .Y(n267) );
  AO21X1 U266 ( .A0(n42), .A1(n26), .B0(n462), .Y(n322) );
  OAI22XL U267 ( .A0(n42), .A1(n463), .B0(n26), .B1(n462), .Y(n108) );
  OAI22XL U268 ( .A0(n42), .A1(n464), .B0(n26), .B1(n463), .Y(n323) );
  OAI22XL U269 ( .A0(n42), .A1(n465), .B0(n26), .B1(n464), .Y(n324) );
  OAI22XL U270 ( .A0(n42), .A1(n466), .B0(n26), .B1(n465), .Y(n325) );
  OAI22XL U271 ( .A0(n42), .A1(n467), .B0(n26), .B1(n466), .Y(n326) );
  OAI22XL U272 ( .A0(n42), .A1(n468), .B0(n26), .B1(n467), .Y(n327) );
  OAI22XL U273 ( .A0(n42), .A1(n469), .B0(n26), .B1(n468), .Y(n328) );
  OAI22XL U274 ( .A0(n41), .A1(n470), .B0(n26), .B1(n469), .Y(n329) );
  OAI22XL U275 ( .A0(n41), .A1(n471), .B0(n25), .B1(n470), .Y(n330) );
  OAI22XL U276 ( .A0(n41), .A1(n472), .B0(n25), .B1(n471), .Y(n331) );
  OAI22XL U277 ( .A0(n41), .A1(n473), .B0(n25), .B1(n472), .Y(n332) );
  OAI22XL U278 ( .A0(n41), .A1(n474), .B0(n25), .B1(n473), .Y(n333) );
  OAI22XL U279 ( .A0(n41), .A1(n475), .B0(n25), .B1(n474), .Y(n334) );
  OAI22XL U280 ( .A0(n41), .A1(n476), .B0(n25), .B1(n475), .Y(n335) );
  OAI22XL U281 ( .A0(n41), .A1(n477), .B0(n25), .B1(n476), .Y(n336) );
  OAI22XL U282 ( .A0(n41), .A1(n478), .B0(n25), .B1(n477), .Y(n337) );
  NOR2BX1 U283 ( .AN(n49), .B(n25), .Y(n338) );
  XNOR2X1 U284 ( .A(n9), .B(n552), .Y(n462) );
  XNOR2X1 U285 ( .A(n9), .B(n553), .Y(n463) );
  XNOR2X1 U286 ( .A(n9), .B(n554), .Y(n464) );
  XNOR2X1 U287 ( .A(n9), .B(n555), .Y(n465) );
  XNOR2X1 U288 ( .A(n9), .B(n556), .Y(n466) );
  XNOR2X1 U289 ( .A(n9), .B(n557), .Y(n467) );
  XNOR2X1 U290 ( .A(n9), .B(n558), .Y(n468) );
  XNOR2X1 U291 ( .A(n9), .B(n559), .Y(n469) );
  XNOR2X1 U292 ( .A(n9), .B(n560), .Y(n470) );
  XNOR2X1 U293 ( .A(n9), .B(n561), .Y(n471) );
  XNOR2X1 U294 ( .A(n9), .B(n562), .Y(n472) );
  XNOR2X1 U295 ( .A(n9), .B(n563), .Y(n473) );
  XNOR2X1 U296 ( .A(n9), .B(n564), .Y(n474) );
  XNOR2X1 U297 ( .A(n9), .B(n565), .Y(n475) );
  XNOR2X1 U298 ( .A(n9), .B(n566), .Y(n476) );
  XNOR2X1 U299 ( .A(n9), .B(n567), .Y(n477) );
  XNOR2X1 U300 ( .A(n9), .B(n49), .Y(n478) );
  NAND2BX1 U301 ( .AN(n49), .B(n9), .Y(n479) );
  OAI22XL U302 ( .A0(n40), .A1(n597), .B0(n24), .B1(n497), .Y(n268) );
  AO21X1 U303 ( .A0(n40), .A1(n24), .B0(n480), .Y(n339) );
  OAI22XL U304 ( .A0(n40), .A1(n481), .B0(n24), .B1(n480), .Y(n340) );
  OAI22XL U305 ( .A0(n40), .A1(n482), .B0(n24), .B1(n481), .Y(n341) );
  OAI22XL U306 ( .A0(n40), .A1(n483), .B0(n24), .B1(n482), .Y(n342) );
  OAI22XL U307 ( .A0(n40), .A1(n484), .B0(n24), .B1(n483), .Y(n343) );
  OAI22XL U308 ( .A0(n40), .A1(n485), .B0(n24), .B1(n484), .Y(n344) );
  OAI22XL U309 ( .A0(n40), .A1(n486), .B0(n24), .B1(n485), .Y(n345) );
  OAI22XL U310 ( .A0(n40), .A1(n487), .B0(n24), .B1(n486), .Y(n346) );
  OAI22XL U311 ( .A0(n39), .A1(n488), .B0(n24), .B1(n487), .Y(n347) );
  OAI22XL U312 ( .A0(n39), .A1(n489), .B0(n23), .B1(n488), .Y(n348) );
  OAI22XL U313 ( .A0(n39), .A1(n490), .B0(n23), .B1(n489), .Y(n349) );
  OAI22XL U314 ( .A0(n39), .A1(n491), .B0(n23), .B1(n490), .Y(n350) );
  OAI22XL U315 ( .A0(n39), .A1(n492), .B0(n23), .B1(n491), .Y(n351) );
  OAI22XL U316 ( .A0(n39), .A1(n493), .B0(n23), .B1(n492), .Y(n352) );
  OAI22XL U317 ( .A0(n39), .A1(n494), .B0(n23), .B1(n493), .Y(n353) );
  OAI22XL U318 ( .A0(n39), .A1(n495), .B0(n23), .B1(n494), .Y(n354) );
  OAI22XL U319 ( .A0(n39), .A1(n496), .B0(n23), .B1(n495), .Y(n355) );
  NOR2BX1 U320 ( .AN(n49), .B(n23), .Y(n356) );
  XNOR2X1 U321 ( .A(n7), .B(n552), .Y(n480) );
  XNOR2X1 U322 ( .A(n7), .B(n553), .Y(n481) );
  XNOR2X1 U323 ( .A(n7), .B(n554), .Y(n482) );
  XNOR2X1 U324 ( .A(n7), .B(n555), .Y(n483) );
  XNOR2X1 U325 ( .A(n7), .B(n556), .Y(n484) );
  XNOR2X1 U326 ( .A(n7), .B(n557), .Y(n485) );
  XNOR2X1 U327 ( .A(n7), .B(n558), .Y(n486) );
  XNOR2X1 U328 ( .A(n7), .B(n559), .Y(n487) );
  XNOR2X1 U329 ( .A(n7), .B(n560), .Y(n488) );
  XNOR2X1 U330 ( .A(n7), .B(n561), .Y(n489) );
  XNOR2X1 U331 ( .A(n7), .B(n562), .Y(n490) );
  XNOR2X1 U332 ( .A(n7), .B(n563), .Y(n491) );
  XNOR2X1 U333 ( .A(n7), .B(n564), .Y(n492) );
  XNOR2X1 U334 ( .A(n7), .B(n565), .Y(n493) );
  XNOR2X1 U335 ( .A(n7), .B(n566), .Y(n494) );
  XNOR2X1 U336 ( .A(n7), .B(n567), .Y(n495) );
  XNOR2X1 U337 ( .A(n7), .B(n49), .Y(n496) );
  NAND2BX1 U338 ( .AN(n49), .B(n7), .Y(n497) );
  OAI22XL U339 ( .A0(n38), .A1(n598), .B0(n22), .B1(n515), .Y(n269) );
  AO21X1 U340 ( .A0(n38), .A1(n22), .B0(n498), .Y(n357) );
  OAI22XL U341 ( .A0(n38), .A1(n499), .B0(n22), .B1(n498), .Y(n140) );
  OAI22XL U342 ( .A0(n38), .A1(n500), .B0(n22), .B1(n499), .Y(n358) );
  OAI22XL U343 ( .A0(n38), .A1(n501), .B0(n22), .B1(n500), .Y(n359) );
  OAI22XL U344 ( .A0(n38), .A1(n502), .B0(n22), .B1(n501), .Y(n360) );
  OAI22XL U345 ( .A0(n38), .A1(n503), .B0(n22), .B1(n502), .Y(n361) );
  OAI22XL U346 ( .A0(n38), .A1(n504), .B0(n22), .B1(n503), .Y(n362) );
  OAI22XL U347 ( .A0(n38), .A1(n505), .B0(n22), .B1(n504), .Y(n363) );
  OAI22XL U348 ( .A0(n37), .A1(n506), .B0(n22), .B1(n505), .Y(n364) );
  OAI22XL U349 ( .A0(n37), .A1(n507), .B0(n21), .B1(n506), .Y(n365) );
  OAI22XL U350 ( .A0(n37), .A1(n508), .B0(n21), .B1(n507), .Y(n366) );
  OAI22XL U351 ( .A0(n37), .A1(n509), .B0(n21), .B1(n508), .Y(n367) );
  OAI22XL U352 ( .A0(n37), .A1(n510), .B0(n21), .B1(n509), .Y(n368) );
  OAI22XL U353 ( .A0(n37), .A1(n511), .B0(n21), .B1(n510), .Y(n369) );
  OAI22XL U354 ( .A0(n37), .A1(n512), .B0(n21), .B1(n511), .Y(n370) );
  OAI22XL U355 ( .A0(n37), .A1(n513), .B0(n21), .B1(n512), .Y(n371) );
  OAI22XL U356 ( .A0(n37), .A1(n514), .B0(n21), .B1(n513), .Y(n372) );
  NOR2BX1 U357 ( .AN(n49), .B(n21), .Y(n373) );
  XNOR2X1 U358 ( .A(n5), .B(n552), .Y(n498) );
  XNOR2X1 U359 ( .A(n5), .B(n553), .Y(n499) );
  XNOR2X1 U360 ( .A(n5), .B(n554), .Y(n500) );
  XNOR2X1 U361 ( .A(n5), .B(n555), .Y(n501) );
  XNOR2X1 U362 ( .A(n5), .B(n556), .Y(n502) );
  XNOR2X1 U363 ( .A(n5), .B(n557), .Y(n503) );
  XNOR2X1 U364 ( .A(n5), .B(n558), .Y(n504) );
  XNOR2X1 U365 ( .A(n5), .B(n559), .Y(n505) );
  XNOR2X1 U366 ( .A(n5), .B(n560), .Y(n506) );
  XNOR2X1 U367 ( .A(n5), .B(n561), .Y(n507) );
  XNOR2X1 U368 ( .A(n5), .B(n562), .Y(n508) );
  XNOR2X1 U369 ( .A(n5), .B(n563), .Y(n509) );
  XNOR2X1 U370 ( .A(n5), .B(n564), .Y(n510) );
  XNOR2X1 U371 ( .A(n5), .B(n565), .Y(n511) );
  XNOR2X1 U372 ( .A(n5), .B(n566), .Y(n512) );
  XNOR2X1 U373 ( .A(n5), .B(n567), .Y(n513) );
  XNOR2X1 U374 ( .A(n5), .B(n49), .Y(n514) );
  NAND2BX1 U375 ( .AN(n49), .B(n5), .Y(n515) );
  OAI22XL U376 ( .A0(n36), .A1(n599), .B0(n20), .B1(n533), .Y(n270) );
  AO21X1 U377 ( .A0(n36), .A1(n20), .B0(n516), .Y(n374) );
  OAI22XL U378 ( .A0(n36), .A1(n517), .B0(n20), .B1(n516), .Y(n160) );
  OAI22XL U379 ( .A0(n36), .A1(n518), .B0(n20), .B1(n517), .Y(n375) );
  OAI22XL U380 ( .A0(n36), .A1(n519), .B0(n20), .B1(n518), .Y(n376) );
  OAI22XL U381 ( .A0(n36), .A1(n520), .B0(n20), .B1(n519), .Y(n377) );
  OAI22XL U382 ( .A0(n36), .A1(n521), .B0(n20), .B1(n520), .Y(n378) );
  OAI22XL U383 ( .A0(n36), .A1(n522), .B0(n20), .B1(n521), .Y(n379) );
  OAI22XL U384 ( .A0(n36), .A1(n523), .B0(n20), .B1(n522), .Y(n380) );
  OAI22XL U385 ( .A0(n35), .A1(n524), .B0(n20), .B1(n523), .Y(n381) );
  OAI22XL U386 ( .A0(n35), .A1(n525), .B0(n19), .B1(n524), .Y(n382) );
  OAI22XL U387 ( .A0(n35), .A1(n526), .B0(n19), .B1(n525), .Y(n383) );
  OAI22XL U388 ( .A0(n35), .A1(n527), .B0(n19), .B1(n526), .Y(n384) );
  OAI22XL U389 ( .A0(n35), .A1(n528), .B0(n19), .B1(n527), .Y(n385) );
  OAI22XL U390 ( .A0(n35), .A1(n529), .B0(n19), .B1(n528), .Y(n386) );
  OAI22XL U391 ( .A0(n35), .A1(n530), .B0(n19), .B1(n529), .Y(n387) );
  OAI22XL U392 ( .A0(n35), .A1(n531), .B0(n19), .B1(n530), .Y(n388) );
  OAI22XL U393 ( .A0(n35), .A1(n532), .B0(n19), .B1(n531), .Y(n389) );
  NOR2BX1 U394 ( .AN(n49), .B(n19), .Y(n390) );
  XNOR2X1 U395 ( .A(n3), .B(n552), .Y(n516) );
  XNOR2X1 U396 ( .A(n3), .B(n553), .Y(n517) );
  XNOR2X1 U397 ( .A(n3), .B(n554), .Y(n518) );
  XNOR2X1 U398 ( .A(n3), .B(n555), .Y(n519) );
  XNOR2X1 U399 ( .A(n3), .B(n556), .Y(n520) );
  XNOR2X1 U400 ( .A(n3), .B(n557), .Y(n521) );
  XNOR2X1 U401 ( .A(n3), .B(n558), .Y(n522) );
  XNOR2X1 U402 ( .A(n3), .B(n559), .Y(n523) );
  XNOR2X1 U403 ( .A(n3), .B(n560), .Y(n524) );
  XNOR2X1 U404 ( .A(n3), .B(n561), .Y(n525) );
  XNOR2X1 U405 ( .A(n3), .B(n562), .Y(n526) );
  XNOR2X1 U406 ( .A(n3), .B(n563), .Y(n527) );
  XNOR2X1 U407 ( .A(n3), .B(n564), .Y(n528) );
  XNOR2X1 U408 ( .A(n3), .B(n565), .Y(n529) );
  XNOR2X1 U409 ( .A(n3), .B(n566), .Y(n530) );
  XNOR2X1 U410 ( .A(n3), .B(n567), .Y(n531) );
  XNOR2X1 U411 ( .A(n3), .B(n49), .Y(n532) );
  NAND2BX1 U412 ( .AN(n49), .B(n3), .Y(n533) );
  OAI22XL U413 ( .A0(n34), .A1(n600), .B0(n551), .B1(n18), .Y(n271) );
  AO21X1 U414 ( .A0(n34), .A1(n18), .B0(n534), .Y(n391) );
  OAI22XL U415 ( .A0(n34), .A1(n535), .B0(n534), .B1(n18), .Y(n392) );
  OAI22XL U416 ( .A0(n34), .A1(n536), .B0(n535), .B1(n18), .Y(n393) );
  OAI22XL U417 ( .A0(n34), .A1(n537), .B0(n536), .B1(n18), .Y(n394) );
  OAI22XL U418 ( .A0(n34), .A1(n538), .B0(n537), .B1(n18), .Y(n395) );
  OAI22XL U419 ( .A0(n34), .A1(n539), .B0(n538), .B1(n18), .Y(n396) );
  OAI22XL U420 ( .A0(n34), .A1(n540), .B0(n539), .B1(n18), .Y(n397) );
  OAI22XL U421 ( .A0(n34), .A1(n541), .B0(n540), .B1(n18), .Y(n398) );
  OAI22XL U422 ( .A0(n33), .A1(n542), .B0(n541), .B1(n18), .Y(n399) );
  OAI22XL U423 ( .A0(n33), .A1(n543), .B0(n542), .B1(n17), .Y(n400) );
  OAI22XL U424 ( .A0(n33), .A1(n544), .B0(n543), .B1(n17), .Y(n401) );
  OAI22XL U425 ( .A0(n33), .A1(n545), .B0(n544), .B1(n17), .Y(n402) );
  OAI22XL U426 ( .A0(n33), .A1(n546), .B0(n545), .B1(n17), .Y(n403) );
  OAI22XL U427 ( .A0(n33), .A1(n547), .B0(n546), .B1(n17), .Y(n404) );
  OAI22XL U428 ( .A0(n33), .A1(n548), .B0(n547), .B1(n17), .Y(n405) );
  OAI22XL U429 ( .A0(n33), .A1(n549), .B0(n548), .B1(n17), .Y(n406) );
  OAI22XL U430 ( .A0(n33), .A1(n550), .B0(n549), .B1(n17), .Y(n407) );
  NOR2BX1 U431 ( .AN(n49), .B(n17), .Y(product_0_) );
  XNOR2X1 U432 ( .A(n1), .B(n552), .Y(n534) );
  XNOR2X1 U433 ( .A(n1), .B(n553), .Y(n535) );
  XNOR2X1 U434 ( .A(n1), .B(n554), .Y(n536) );
  XNOR2X1 U435 ( .A(n1), .B(n555), .Y(n537) );
  XNOR2X1 U436 ( .A(n1), .B(n556), .Y(n538) );
  XNOR2X1 U437 ( .A(n1), .B(n557), .Y(n539) );
  XNOR2X1 U438 ( .A(n1), .B(n558), .Y(n540) );
  XNOR2X1 U439 ( .A(n1), .B(n559), .Y(n541) );
  XNOR2X1 U440 ( .A(n1), .B(n560), .Y(n542) );
  XNOR2X1 U441 ( .A(n1), .B(n561), .Y(n543) );
  XNOR2X1 U442 ( .A(n1), .B(n562), .Y(n544) );
  XNOR2X1 U443 ( .A(n1), .B(n563), .Y(n545) );
  XNOR2X1 U444 ( .A(n1), .B(n564), .Y(n546) );
  XNOR2X1 U445 ( .A(n1), .B(n565), .Y(n547) );
  XNOR2X1 U446 ( .A(n1), .B(n566), .Y(n548) );
  XNOR2X1 U447 ( .A(n1), .B(n567), .Y(n549) );
  XNOR2X1 U448 ( .A(n1), .B(n49), .Y(n550) );
  NAND2BX1 U449 ( .AN(n49), .B(n1), .Y(n551) );
  CLKINVX1 U466 ( .A(n15), .Y(n593) );
  CLKINVX1 U467 ( .A(n13), .Y(n594) );
  CLKINVX1 U468 ( .A(n11), .Y(n595) );
  CLKINVX1 U469 ( .A(n9), .Y(n596) );
  CLKINVX1 U470 ( .A(n7), .Y(n597) );
  CLKINVX1 U471 ( .A(n5), .Y(n598) );
  CLKINVX1 U472 ( .A(n3), .Y(n599) );
  CLKINVX1 U473 ( .A(n1), .Y(n600) );
  NAND2X1 U474 ( .A(n569), .B(n585), .Y(n577) );
  XOR2X1 U475 ( .A(a[14]), .B(a[15]), .Y(n569) );
  XNOR2X1 U476 ( .A(a[14]), .B(a[13]), .Y(n585) );
  NAND2X1 U477 ( .A(n570), .B(n586), .Y(n578) );
  XOR2X1 U478 ( .A(a[12]), .B(a[13]), .Y(n570) );
  XNOR2X1 U479 ( .A(a[12]), .B(a[11]), .Y(n586) );
  NAND2X1 U480 ( .A(n571), .B(n587), .Y(n579) );
  XOR2X1 U481 ( .A(a[10]), .B(a[11]), .Y(n571) );
  XNOR2X1 U482 ( .A(a[10]), .B(a[9]), .Y(n587) );
  NAND2X1 U483 ( .A(n572), .B(n588), .Y(n580) );
  XOR2X1 U484 ( .A(a[8]), .B(a[9]), .Y(n572) );
  XNOR2X1 U485 ( .A(a[8]), .B(a[7]), .Y(n588) );
  NAND2X1 U486 ( .A(n573), .B(n589), .Y(n581) );
  XOR2X1 U487 ( .A(a[6]), .B(a[7]), .Y(n573) );
  XNOR2X1 U488 ( .A(a[6]), .B(a[5]), .Y(n589) );
  NAND2X1 U489 ( .A(n574), .B(n590), .Y(n582) );
  XOR2X1 U490 ( .A(a[4]), .B(a[5]), .Y(n574) );
  XNOR2X1 U491 ( .A(a[4]), .B(a[3]), .Y(n590) );
  NAND2X1 U492 ( .A(n575), .B(n591), .Y(n583) );
  XOR2X1 U493 ( .A(a[2]), .B(a[3]), .Y(n575) );
  XNOR2X1 U494 ( .A(a[2]), .B(a[1]), .Y(n591) );
  NAND2X1 U495 ( .A(n576), .B(n592), .Y(n584) );
  XOR2X1 U496 ( .A(a[0]), .B(a[1]), .Y(n576) );
  CLKINVX1 U497 ( .A(a[0]), .Y(n592) );
  CLKBUFX3 U500 ( .A(b_2_), .Y(n566) );
  CLKBUFX3 U501 ( .A(b_4_), .Y(n564) );
  CLKBUFX3 U502 ( .A(b_5_), .Y(n563) );
  CLKBUFX3 U503 ( .A(b_6_), .Y(n562) );
  CLKBUFX3 U504 ( .A(b_0_), .Y(n49) );
  CLKBUFX3 U505 ( .A(b_3_), .Y(n565) );
  CLKBUFX3 U506 ( .A(b_9_), .Y(n559) );
  CLKBUFX3 U507 ( .A(b_12_), .Y(n556) );
  CLKBUFX3 U508 ( .A(b_7_), .Y(n561) );
  CLKBUFX3 U509 ( .A(b_14_), .Y(n554) );
  CLKBUFX3 U510 ( .A(n591), .Y(n20) );
  CLKBUFX3 U511 ( .A(n590), .Y(n22) );
  CLKBUFX3 U512 ( .A(n588), .Y(n26) );
  CLKBUFX3 U513 ( .A(n589), .Y(n24) );
  CLKBUFX3 U514 ( .A(n585), .Y(n32) );
  CLKBUFX3 U515 ( .A(n586), .Y(n30) );
  CLKBUFX3 U516 ( .A(n587), .Y(n28) );
  CLKBUFX3 U517 ( .A(b_10_), .Y(n558) );
  CLKBUFX3 U518 ( .A(b_15_), .Y(n553) );
  CLKBUFX3 U519 ( .A(n591), .Y(n19) );
  CLKBUFX3 U520 ( .A(n590), .Y(n21) );
  CLKBUFX3 U521 ( .A(n589), .Y(n23) );
  CLKBUFX3 U522 ( .A(n588), .Y(n25) );
  CLKBUFX3 U523 ( .A(n587), .Y(n27) );
  CLKBUFX3 U524 ( .A(n586), .Y(n29) );
  CLKBUFX3 U525 ( .A(n585), .Y(n31) );
  CLKBUFX3 U526 ( .A(b_8_), .Y(n560) );
  CLKBUFX3 U527 ( .A(b_11_), .Y(n557) );
  CLKBUFX3 U528 ( .A(b_16_), .Y(n552) );
  CLKBUFX3 U529 ( .A(n583), .Y(n35) );
  CLKBUFX3 U530 ( .A(n582), .Y(n37) );
  CLKBUFX3 U531 ( .A(n581), .Y(n39) );
  CLKBUFX3 U532 ( .A(n580), .Y(n41) );
  CLKBUFX3 U533 ( .A(n579), .Y(n43) );
  CLKBUFX3 U534 ( .A(n578), .Y(n45) );
  CLKBUFX3 U535 ( .A(n577), .Y(n47) );
  CLKBUFX3 U536 ( .A(n584), .Y(n33) );
  CLKBUFX3 U537 ( .A(n583), .Y(n36) );
  CLKBUFX3 U538 ( .A(n582), .Y(n38) );
  CLKBUFX3 U539 ( .A(n580), .Y(n42) );
  CLKBUFX3 U540 ( .A(n581), .Y(n40) );
  CLKBUFX3 U541 ( .A(n577), .Y(n48) );
  CLKBUFX3 U542 ( .A(n578), .Y(n46) );
  CLKBUFX3 U543 ( .A(n579), .Y(n44) );
  CLKBUFX3 U544 ( .A(n584), .Y(n34) );
  CLKBUFX3 U545 ( .A(n592), .Y(n18) );
  CLKBUFX3 U546 ( .A(n592), .Y(n17) );
  CLKBUFX3 U547 ( .A(b_1_), .Y(n567) );
  CLKBUFX3 U548 ( .A(b_13_), .Y(n555) );
  CLKBUFX3 U549 ( .A(a[1]), .Y(n1) );
  CLKBUFX3 U550 ( .A(a[3]), .Y(n3) );
  CLKBUFX3 U551 ( .A(a[5]), .Y(n5) );
  CLKBUFX3 U552 ( .A(a[7]), .Y(n7) );
  CLKBUFX3 U553 ( .A(a[9]), .Y(n9) );
  CLKBUFX3 U554 ( .A(a[11]), .Y(n11) );
  CLKBUFX3 U555 ( .A(a[13]), .Y(n13) );
  CLKBUFX3 U556 ( .A(a[15]), .Y(n15) );
endmodule


module FAS_DW_mult_uns_5 ( a, b, product_31_, product_30_, product_29_, 
        product_28_, product_27_, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_, product_14_, 
        product_13_, product_12_, product_11_, product_10_, product_9_, 
        product_8_, product_7_, product_6_, product_5_, product_4_, product_3_, 
        product_2_, product_1_, product_0_ );
  input [31:0] a;
  input b;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;

  NOR2X1 U3 ( .A(n2), .B(n3), .Y(product_31_) );
  NOR2X1 U4 ( .A(n2), .B(n4), .Y(product_30_) );
  NOR2X1 U5 ( .A(n2), .B(n5), .Y(product_29_) );
  NOR2X1 U6 ( .A(n2), .B(n6), .Y(product_28_) );
  NOR2X1 U7 ( .A(n2), .B(n7), .Y(product_27_) );
  NOR2X1 U8 ( .A(n2), .B(n8), .Y(product_26_) );
  NOR2X1 U9 ( .A(n2), .B(n9), .Y(product_25_) );
  NOR2X1 U10 ( .A(n2), .B(n10), .Y(product_24_) );
  NOR2X1 U11 ( .A(n2), .B(n11), .Y(product_23_) );
  NOR2X1 U12 ( .A(n2), .B(n12), .Y(product_22_) );
  NOR2X1 U13 ( .A(n2), .B(n13), .Y(product_21_) );
  NOR2X1 U14 ( .A(n2), .B(n14), .Y(product_20_) );
  NOR2X1 U15 ( .A(n2), .B(n15), .Y(product_19_) );
  NOR2X1 U16 ( .A(n2), .B(n16), .Y(product_18_) );
  NOR2X1 U17 ( .A(n2), .B(n17), .Y(product_17_) );
  NOR2X1 U18 ( .A(n2), .B(n18), .Y(product_16_) );
  NOR2X1 U19 ( .A(n1), .B(n19), .Y(product_15_) );
  NOR2X1 U20 ( .A(n1), .B(n20), .Y(product_14_) );
  NOR2X1 U21 ( .A(n1), .B(n21), .Y(product_13_) );
  NOR2X1 U22 ( .A(n1), .B(n22), .Y(product_12_) );
  NOR2X1 U23 ( .A(n1), .B(n23), .Y(product_11_) );
  NOR2X1 U24 ( .A(n1), .B(n24), .Y(product_10_) );
  NOR2X1 U25 ( .A(n1), .B(n25), .Y(product_9_) );
  NOR2X1 U26 ( .A(n1), .B(n26), .Y(product_8_) );
  NOR2X1 U27 ( .A(n1), .B(n27), .Y(product_7_) );
  NOR2X1 U28 ( .A(n1), .B(n28), .Y(product_6_) );
  NOR2X1 U29 ( .A(n1), .B(n29), .Y(product_5_) );
  NOR2X1 U30 ( .A(n1), .B(n30), .Y(product_4_) );
  NOR2X1 U31 ( .A(n1), .B(n31), .Y(product_3_) );
  NOR2X1 U32 ( .A(n1), .B(n32), .Y(product_2_) );
  NOR2X1 U33 ( .A(n1), .B(n33), .Y(product_1_) );
  NOR2X1 U34 ( .A(n1), .B(n34), .Y(product_0_) );
  CLKINVX1 U70 ( .A(a[1]), .Y(n33) );
  CLKINVX1 U71 ( .A(a[0]), .Y(n34) );
  CLKBUFX3 U72 ( .A(n35), .Y(n1) );
  CLKBUFX3 U73 ( .A(n35), .Y(n2) );
  CLKINVX1 U74 ( .A(b), .Y(n35) );
  CLKINVX1 U75 ( .A(a[2]), .Y(n32) );
  CLKINVX1 U76 ( .A(a[3]), .Y(n31) );
  CLKINVX1 U77 ( .A(a[4]), .Y(n30) );
  CLKINVX1 U78 ( .A(a[5]), .Y(n29) );
  CLKINVX1 U79 ( .A(a[6]), .Y(n28) );
  CLKINVX1 U80 ( .A(a[7]), .Y(n27) );
  CLKINVX1 U81 ( .A(a[8]), .Y(n26) );
  CLKINVX1 U82 ( .A(a[9]), .Y(n25) );
  CLKINVX1 U83 ( .A(a[10]), .Y(n24) );
  CLKINVX1 U84 ( .A(a[11]), .Y(n23) );
  CLKINVX1 U85 ( .A(a[12]), .Y(n22) );
  CLKINVX1 U86 ( .A(a[13]), .Y(n21) );
  CLKINVX1 U87 ( .A(a[14]), .Y(n20) );
  CLKINVX1 U88 ( .A(a[15]), .Y(n19) );
  CLKINVX1 U89 ( .A(a[16]), .Y(n18) );
  CLKINVX1 U90 ( .A(a[17]), .Y(n17) );
  CLKINVX1 U91 ( .A(a[18]), .Y(n16) );
  CLKINVX1 U92 ( .A(a[19]), .Y(n15) );
  CLKINVX1 U93 ( .A(a[20]), .Y(n14) );
  CLKINVX1 U94 ( .A(a[21]), .Y(n13) );
  CLKINVX1 U95 ( .A(a[22]), .Y(n12) );
  CLKINVX1 U96 ( .A(a[23]), .Y(n11) );
  CLKINVX1 U97 ( .A(a[24]), .Y(n10) );
  CLKINVX1 U98 ( .A(a[25]), .Y(n9) );
  CLKINVX1 U99 ( .A(a[26]), .Y(n8) );
  CLKINVX1 U100 ( .A(a[27]), .Y(n7) );
  CLKINVX1 U101 ( .A(a[28]), .Y(n6) );
  CLKINVX1 U102 ( .A(a[29]), .Y(n5) );
  CLKINVX1 U103 ( .A(a[30]), .Y(n4) );
  CLKINVX1 U104 ( .A(a[31]), .Y(n3) );
endmodule


module FAS_DW_mult_tc_27 ( a, b_17_, b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, 
        b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input [15:0] a;
  input b_17_, b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_, b_8_,
         b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n3, n5, n7, n9, n11, n13, n15, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n697;

  XOR2X1 U51 ( .A(n52), .B(n51), .Y(product_31_) );
  XOR2X1 U52 ( .A(n83), .B(n697), .Y(n51) );
  ADDFXL U53 ( .A(n84), .B(n85), .CI(n53), .CO(n52), .S(product_30_) );
  ADDFXL U54 ( .A(n90), .B(n86), .CI(n54), .CO(n53), .S(product_29_) );
  ADDFXL U55 ( .A(n93), .B(n91), .CI(n55), .CO(n54), .S(product_28_) );
  ADDFXL U56 ( .A(n94), .B(n98), .CI(n56), .CO(n55), .S(product_27_) );
  ADDFXL U57 ( .A(n99), .B(n103), .CI(n57), .CO(n56), .S(product_26_) );
  ADDFXL U58 ( .A(n104), .B(n110), .CI(n58), .CO(n57), .S(product_25_) );
  ADDFXL U59 ( .A(n111), .B(n116), .CI(n59), .CO(n58), .S(product_24_) );
  ADDFXL U60 ( .A(n117), .B(n124), .CI(n60), .CO(n59), .S(product_23_) );
  ADDFXL U61 ( .A(n132), .B(n125), .CI(n61), .CO(n60), .S(product_22_) );
  ADDFXL U62 ( .A(n142), .B(n133), .CI(n62), .CO(n61), .S(product_21_) );
  ADDFXL U63 ( .A(n143), .B(n151), .CI(n63), .CO(n62), .S(product_20_) );
  ADDFXL U64 ( .A(n152), .B(n162), .CI(n64), .CO(n63), .S(product_19_) );
  ADDFXL U65 ( .A(n163), .B(n173), .CI(n65), .CO(n64), .S(product_18_) );
  ADDFXL U66 ( .A(n174), .B(n184), .CI(n66), .CO(n65), .S(product_17_) );
  ADDFXL U67 ( .A(n185), .B(n195), .CI(n67), .CO(n66), .S(product_16_) );
  ADDFXL U68 ( .A(n196), .B(n206), .CI(n68), .CO(n67), .S(product_15_) );
  ADDFXL U69 ( .A(n207), .B(n215), .CI(n69), .CO(n68), .S(product_14_) );
  ADDFXL U70 ( .A(n216), .B(n225), .CI(n70), .CO(n69), .S(product_13_) );
  ADDFXL U71 ( .A(n226), .B(n233), .CI(n71), .CO(n70), .S(product_12_) );
  ADDFXL U72 ( .A(n234), .B(n241), .CI(n72), .CO(n71), .S(product_11_) );
  ADDFXL U73 ( .A(n242), .B(n247), .CI(n73), .CO(n72), .S(product_10_) );
  ADDFXL U74 ( .A(n248), .B(n254), .CI(n74), .CO(n73), .S(product_9_) );
  ADDFXL U75 ( .A(n255), .B(n259), .CI(n75), .CO(n74), .S(product_8_) );
  ADDFXL U76 ( .A(n260), .B(n264), .CI(n76), .CO(n75), .S(product_7_) );
  ADDFXL U77 ( .A(n265), .B(n266), .CI(n77), .CO(n76), .S(product_6_) );
  ADDFXL U78 ( .A(n267), .B(n270), .CI(n78), .CO(n77), .S(product_5_) );
  ADDFXL U79 ( .A(n271), .B(n272), .CI(n79), .CO(n78), .S(product_4_) );
  ADDFXL U80 ( .A(n273), .B(n406), .CI(n80), .CO(n79), .S(product_3_) );
  ADDFXL U81 ( .A(n424), .B(n407), .CI(n81), .CO(n80), .S(product_2_) );
  ADDHXL U82 ( .A(n281), .B(n425), .CO(n81), .S(product_1_) );
  ADDFXL U84 ( .A(n283), .B(n87), .CI(n300), .CO(n83), .S(n84) );
  ADDFXL U85 ( .A(n88), .B(n284), .CI(n89), .CO(n85), .S(n86) );
  CLKINVX1 U86 ( .A(n87), .Y(n88) );
  CMPR42X1 U87 ( .A(n95), .B(n285), .C(n301), .D(n318), .ICI(n92), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U88 ( .A(n302), .B(n286), .C(n96), .D(n100), .ICI(n97), .S(n94), 
        .ICO(n92), .CO(n93) );
  CLKINVX1 U89 ( .A(n95), .Y(n96) );
  CMPR42X1 U90 ( .A(n319), .B(n303), .C(n105), .D(n101), .ICI(n102), .S(n99), 
        .ICO(n97), .CO(n98) );
  ADDFXL U91 ( .A(n107), .B(n287), .CI(n335), .CO(n100), .S(n101) );
  CMPR42X1 U92 ( .A(n320), .B(n112), .C(n106), .D(n113), .ICI(n109), .S(n104), 
        .ICO(n102), .CO(n103) );
  ADDFXL U93 ( .A(n304), .B(n288), .CI(n108), .CO(n105), .S(n106) );
  CLKINVX1 U94 ( .A(n107), .Y(n108) );
  CMPR42X1 U95 ( .A(n321), .B(n305), .C(n119), .D(n114), .ICI(n115), .S(n111), 
        .ICO(n109), .CO(n110) );
  CMPR42X1 U96 ( .A(n289), .B(n121), .C(n336), .D(n353), .ICI(n118), .S(n114), 
        .ICO(n112), .CO(n113) );
  CMPR42X1 U97 ( .A(n290), .B(n129), .C(n127), .D(n120), .ICI(n123), .S(n117), 
        .ICO(n115), .CO(n116) );
  CMPR42X1 U98 ( .A(n306), .B(n354), .C(n337), .D(n122), .ICI(n126), .S(n120), 
        .ICO(n118), .CO(n119) );
  CLKINVX1 U99 ( .A(n121), .Y(n122) );
  CMPR42X1 U100 ( .A(n137), .B(n130), .C(n135), .D(n128), .ICI(n131), .S(n125), 
        .ICO(n123), .CO(n124) );
  CMPR42X1 U101 ( .A(n307), .B(n338), .C(n322), .D(n139), .ICI(n134), .S(n128), 
        .ICO(n126), .CO(n127) );
  ADDFXL U102 ( .A(n355), .B(n291), .CI(n372), .CO(n129), .S(n130) );
  CMPR42X1 U103 ( .A(n138), .B(n148), .C(n145), .D(n136), .ICI(n141), .S(n133), 
        .ICO(n131), .CO(n132) );
  CMPR42X1 U104 ( .A(n356), .B(n323), .C(n339), .D(n144), .ICI(n147), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFXL U105 ( .A(n292), .B(n308), .CI(n140), .CO(n137), .S(n138) );
  CLKINVX1 U106 ( .A(n139), .Y(n140) );
  CMPR42X1 U107 ( .A(n157), .B(n154), .C(n146), .D(n149), .ICI(n150), .S(n143), 
        .ICO(n141), .CO(n142) );
  CMPR42X1 U108 ( .A(n309), .B(n340), .C(n324), .D(n159), .ICI(n153), .S(n146), 
        .ICO(n144), .CO(n145) );
  CMPR42X1 U109 ( .A(n293), .B(n373), .C(n357), .D(n390), .ICI(n156), .S(n149), 
        .ICO(n147), .CO(n148) );
  CMPR42X1 U110 ( .A(n168), .B(n165), .C(n155), .D(n158), .ICI(n161), .S(n152), 
        .ICO(n150), .CO(n151) );
  CMPR42X1 U111 ( .A(n325), .B(n358), .C(n341), .D(n294), .ICI(n164), .S(n155), 
        .ICO(n153), .CO(n154) );
  CMPR42X1 U112 ( .A(n310), .B(n374), .C(n160), .D(n170), .ICI(n167), .S(n158), 
        .ICO(n156), .CO(n157) );
  CLKINVX1 U113 ( .A(n159), .Y(n160) );
  CMPR42X1 U114 ( .A(n179), .B(n176), .C(n166), .D(n169), .ICI(n172), .S(n163), 
        .ICO(n161), .CO(n162) );
  CMPR42X1 U115 ( .A(n295), .B(n375), .C(n342), .D(n181), .ICI(n175), .S(n166), 
        .ICO(n164), .CO(n165) );
  CMPR42X1 U116 ( .A(n326), .B(n391), .C(n408), .D(n171), .ICI(n178), .S(n169), 
        .ICO(n167), .CO(n168) );
  XNOR2X1 U117 ( .A(n359), .B(n311), .Y(n171) );
  OR2X1 U118 ( .A(n359), .B(n311), .Y(n170) );
  CMPR42X1 U119 ( .A(n190), .B(n187), .C(n180), .D(n177), .ICI(n183), .S(n174), 
        .ICO(n172), .CO(n173) );
  CMPR42X1 U120 ( .A(n312), .B(n360), .C(n343), .D(n182), .ICI(n186), .S(n177), 
        .ICO(n175), .CO(n176) );
  CMPR42X1 U121 ( .A(n327), .B(n392), .C(n376), .D(n192), .ICI(n189), .S(n180), 
        .ICO(n178), .CO(n179) );
  ADDHXL U122 ( .A(n409), .B(n296), .CO(n181), .S(n182) );
  CMPR42X1 U123 ( .A(n201), .B(n198), .C(n191), .D(n188), .ICI(n194), .S(n185), 
        .ICO(n183), .CO(n184) );
  CMPR42X1 U124 ( .A(n313), .B(n328), .C(n361), .D(n193), .ICI(n200), .S(n188), 
        .ICO(n186), .CO(n187) );
  CMPR42X1 U125 ( .A(n344), .B(n393), .C(n377), .D(n203), .ICI(n197), .S(n191), 
        .ICO(n189), .CO(n190) );
  ADDHXL U126 ( .A(n410), .B(n297), .CO(n192), .S(n193) );
  CMPR42X1 U127 ( .A(n212), .B(n209), .C(n202), .D(n199), .ICI(n205), .S(n196), 
        .ICO(n194), .CO(n195) );
  CMPR42X1 U128 ( .A(n314), .B(n329), .C(n345), .D(n211), .ICI(n204), .S(n199), 
        .ICO(n197), .CO(n198) );
  CMPR42X1 U129 ( .A(n274), .B(n298), .C(n394), .D(n362), .ICI(n208), .S(n202), 
        .ICO(n200), .CO(n201) );
  ADDHXL U130 ( .A(n411), .B(n378), .CO(n203), .S(n204) );
  CMPR42X1 U131 ( .A(n220), .B(n213), .C(n218), .D(n210), .ICI(n214), .S(n207), 
        .ICO(n205), .CO(n206) );
  CMPR42X1 U132 ( .A(n395), .B(n346), .C(n363), .D(n379), .ICI(n222), .S(n210), 
        .ICO(n208), .CO(n209) );
  CMPR42X1 U133 ( .A(n299), .B(n412), .C(n315), .D(n330), .ICI(n217), .S(n213), 
        .ICO(n211), .CO(n212) );
  CMPR42X1 U134 ( .A(n230), .B(n221), .C(n228), .D(n219), .ICI(n224), .S(n216), 
        .ICO(n214), .CO(n215) );
  CMPR42X1 U135 ( .A(n331), .B(n364), .C(n347), .D(n316), .ICI(n227), .S(n219), 
        .ICO(n217), .CO(n218) );
  ADDFXL U136 ( .A(n396), .B(n275), .CI(n223), .CO(n220), .S(n221) );
  ADDHXL U137 ( .A(n413), .B(n380), .CO(n222), .S(n223) );
  CMPR42X1 U138 ( .A(n365), .B(n235), .C(n236), .D(n229), .ICI(n232), .S(n226), 
        .ICO(n224), .CO(n225) );
  CMPR42X1 U139 ( .A(n397), .B(n348), .C(n381), .D(n238), .ICI(n231), .S(n229), 
        .ICO(n227), .CO(n228) );
  ADDFXL U140 ( .A(n414), .B(n317), .CI(n332), .CO(n230), .S(n231) );
  CMPR42X1 U141 ( .A(n366), .B(n243), .C(n244), .D(n237), .ICI(n240), .S(n234), 
        .ICO(n232), .CO(n233) );
  CMPR42X1 U142 ( .A(n276), .B(n333), .C(n398), .D(n349), .ICI(n239), .S(n237), 
        .ICO(n235), .CO(n236) );
  ADDHXL U143 ( .A(n415), .B(n382), .CO(n238), .S(n239) );
  CMPR42X1 U144 ( .A(n399), .B(n383), .C(n249), .D(n246), .ICI(n245), .S(n242), 
        .ICO(n240), .CO(n241) );
  CMPR42X1 U145 ( .A(n334), .B(n416), .C(n350), .D(n367), .ICI(n251), .S(n245), 
        .ICO(n243), .CO(n244) );
  CMPR42X1 U146 ( .A(n400), .B(n368), .C(n253), .D(n256), .ICI(n250), .S(n248), 
        .ICO(n246), .CO(n247) );
  ADDFXL U147 ( .A(n351), .B(n277), .CI(n252), .CO(n249), .S(n250) );
  ADDHXL U148 ( .A(n417), .B(n384), .CO(n251), .S(n252) );
  CMPR42X1 U149 ( .A(n401), .B(n385), .C(n261), .D(n258), .ICI(n257), .S(n255), 
        .ICO(n253), .CO(n254) );
  ADDFXL U150 ( .A(n418), .B(n352), .CI(n369), .CO(n256), .S(n257) );
  CMPR42X1 U151 ( .A(n278), .B(n370), .C(n402), .D(n263), .ICI(n262), .S(n260), 
        .ICO(n258), .CO(n259) );
  ADDHXL U152 ( .A(n419), .B(n386), .CO(n261), .S(n262) );
  CMPR42X1 U153 ( .A(n371), .B(n420), .C(n387), .D(n403), .ICI(n268), .S(n265), 
        .ICO(n263), .CO(n264) );
  ADDFXL U154 ( .A(n404), .B(n279), .CI(n269), .CO(n266), .S(n267) );
  ADDHXL U155 ( .A(n421), .B(n388), .CO(n268), .S(n269) );
  ADDFXL U156 ( .A(n422), .B(n389), .CI(n405), .CO(n270), .S(n271) );
  ADDHXL U157 ( .A(n423), .B(n280), .CO(n272), .S(n273) );
  OAI22XL U158 ( .A0(n48), .A1(n620), .B0(n32), .B1(n444), .Y(n274) );
  OAI22XL U160 ( .A0(n48), .A1(n428), .B0(n32), .B1(n427), .Y(n283) );
  OAI22XL U161 ( .A0(n48), .A1(n429), .B0(n32), .B1(n428), .Y(n284) );
  OAI22XL U162 ( .A0(n48), .A1(n430), .B0(n32), .B1(n429), .Y(n285) );
  OAI22XL U163 ( .A0(n48), .A1(n431), .B0(n32), .B1(n430), .Y(n286) );
  OAI22XL U164 ( .A0(n48), .A1(n432), .B0(n32), .B1(n431), .Y(n287) );
  OAI22XL U165 ( .A0(n48), .A1(n433), .B0(n32), .B1(n432), .Y(n288) );
  OAI22XL U166 ( .A0(n48), .A1(n434), .B0(n32), .B1(n433), .Y(n289) );
  OAI22XL U167 ( .A0(n47), .A1(n435), .B0(n31), .B1(n434), .Y(n290) );
  OAI22XL U168 ( .A0(n47), .A1(n436), .B0(n31), .B1(n435), .Y(n291) );
  OAI22XL U169 ( .A0(n47), .A1(n437), .B0(n31), .B1(n436), .Y(n292) );
  OAI22XL U170 ( .A0(n47), .A1(n438), .B0(n31), .B1(n437), .Y(n293) );
  OAI22XL U171 ( .A0(n47), .A1(n439), .B0(n31), .B1(n438), .Y(n294) );
  OAI22XL U172 ( .A0(n47), .A1(n440), .B0(n31), .B1(n439), .Y(n295) );
  OAI22XL U173 ( .A0(n47), .A1(n441), .B0(n31), .B1(n440), .Y(n296) );
  OAI22XL U174 ( .A0(n47), .A1(n442), .B0(n31), .B1(n441), .Y(n297) );
  OAI22XL U175 ( .A0(n47), .A1(n443), .B0(n31), .B1(n442), .Y(n298) );
  NOR2BX1 U176 ( .AN(n49), .B(n31), .Y(n299) );
  XNOR2X1 U177 ( .A(n15), .B(n578), .Y(n426) );
  XNOR2X1 U178 ( .A(n15), .B(n579), .Y(n427) );
  XNOR2X1 U179 ( .A(n15), .B(n580), .Y(n428) );
  XNOR2X1 U180 ( .A(n15), .B(n581), .Y(n429) );
  XNOR2X1 U181 ( .A(n15), .B(n582), .Y(n430) );
  XNOR2X1 U182 ( .A(n15), .B(n583), .Y(n431) );
  XNOR2X1 U183 ( .A(n15), .B(n584), .Y(n432) );
  XNOR2X1 U184 ( .A(n15), .B(n585), .Y(n433) );
  XNOR2X1 U185 ( .A(n15), .B(n586), .Y(n434) );
  XNOR2X1 U186 ( .A(n15), .B(n587), .Y(n435) );
  XNOR2X1 U187 ( .A(n15), .B(n588), .Y(n436) );
  XNOR2X1 U188 ( .A(n15), .B(n589), .Y(n437) );
  XNOR2X1 U189 ( .A(n15), .B(n590), .Y(n438) );
  XNOR2X1 U190 ( .A(n15), .B(n591), .Y(n439) );
  XNOR2X1 U191 ( .A(n15), .B(n592), .Y(n440) );
  XNOR2X1 U192 ( .A(n15), .B(n593), .Y(n441) );
  XNOR2X1 U193 ( .A(n15), .B(n594), .Y(n442) );
  XNOR2X1 U194 ( .A(n15), .B(n49), .Y(n443) );
  NAND2BX1 U195 ( .AN(n49), .B(n15), .Y(n444) );
  OAI22XL U196 ( .A0(n46), .A1(n621), .B0(n30), .B1(n463), .Y(n275) );
  AO21X1 U197 ( .A0(n46), .A1(n30), .B0(n445), .Y(n300) );
  OAI22XL U198 ( .A0(n46), .A1(n446), .B0(n30), .B1(n445), .Y(n87) );
  OAI22XL U199 ( .A0(n46), .A1(n447), .B0(n30), .B1(n446), .Y(n301) );
  OAI22XL U200 ( .A0(n46), .A1(n448), .B0(n30), .B1(n447), .Y(n302) );
  OAI22XL U201 ( .A0(n46), .A1(n449), .B0(n30), .B1(n448), .Y(n303) );
  OAI22XL U202 ( .A0(n46), .A1(n450), .B0(n30), .B1(n449), .Y(n304) );
  OAI22XL U203 ( .A0(n46), .A1(n451), .B0(n30), .B1(n450), .Y(n305) );
  OAI22XL U204 ( .A0(n46), .A1(n452), .B0(n30), .B1(n451), .Y(n306) );
  OAI22XL U205 ( .A0(n46), .A1(n453), .B0(n30), .B1(n452), .Y(n307) );
  OAI22XL U206 ( .A0(n45), .A1(n454), .B0(n29), .B1(n453), .Y(n308) );
  OAI22XL U207 ( .A0(n45), .A1(n455), .B0(n29), .B1(n454), .Y(n309) );
  OAI22XL U208 ( .A0(n45), .A1(n456), .B0(n29), .B1(n455), .Y(n310) );
  OAI22XL U209 ( .A0(n45), .A1(n457), .B0(n29), .B1(n456), .Y(n311) );
  OAI22XL U210 ( .A0(n45), .A1(n458), .B0(n29), .B1(n457), .Y(n312) );
  OAI22XL U211 ( .A0(n45), .A1(n459), .B0(n29), .B1(n458), .Y(n313) );
  OAI22XL U212 ( .A0(n45), .A1(n460), .B0(n29), .B1(n459), .Y(n314) );
  OAI22XL U213 ( .A0(n45), .A1(n461), .B0(n29), .B1(n460), .Y(n315) );
  OAI22XL U214 ( .A0(n45), .A1(n462), .B0(n29), .B1(n461), .Y(n316) );
  NOR2BX1 U215 ( .AN(n49), .B(n29), .Y(n317) );
  XNOR2X1 U216 ( .A(n13), .B(n578), .Y(n445) );
  XNOR2X1 U217 ( .A(n13), .B(n579), .Y(n446) );
  XNOR2X1 U218 ( .A(n13), .B(n580), .Y(n447) );
  XNOR2X1 U219 ( .A(n13), .B(n581), .Y(n448) );
  XNOR2X1 U220 ( .A(n13), .B(n582), .Y(n449) );
  XNOR2X1 U221 ( .A(n13), .B(n583), .Y(n450) );
  XNOR2X1 U222 ( .A(n13), .B(n584), .Y(n451) );
  XNOR2X1 U223 ( .A(n13), .B(n585), .Y(n452) );
  XNOR2X1 U224 ( .A(n13), .B(n586), .Y(n453) );
  XNOR2X1 U225 ( .A(n13), .B(n587), .Y(n454) );
  XNOR2X1 U226 ( .A(n13), .B(n588), .Y(n455) );
  XNOR2X1 U227 ( .A(n13), .B(n589), .Y(n456) );
  XNOR2X1 U228 ( .A(n13), .B(n590), .Y(n457) );
  XNOR2X1 U229 ( .A(n13), .B(n591), .Y(n458) );
  XNOR2X1 U230 ( .A(n13), .B(n592), .Y(n459) );
  XNOR2X1 U231 ( .A(n13), .B(n593), .Y(n460) );
  XNOR2X1 U232 ( .A(n13), .B(n594), .Y(n461) );
  XNOR2X1 U233 ( .A(n13), .B(n49), .Y(n462) );
  NAND2BX1 U234 ( .AN(n49), .B(n13), .Y(n463) );
  OAI22XL U235 ( .A0(n44), .A1(n622), .B0(n28), .B1(n482), .Y(n276) );
  AO21X1 U236 ( .A0(n44), .A1(n28), .B0(n464), .Y(n318) );
  OAI22XL U237 ( .A0(n44), .A1(n465), .B0(n28), .B1(n464), .Y(n95) );
  OAI22XL U238 ( .A0(n44), .A1(n466), .B0(n28), .B1(n465), .Y(n319) );
  OAI22XL U239 ( .A0(n44), .A1(n467), .B0(n28), .B1(n466), .Y(n320) );
  OAI22XL U240 ( .A0(n44), .A1(n468), .B0(n28), .B1(n467), .Y(n321) );
  OAI22XL U241 ( .A0(n44), .A1(n469), .B0(n28), .B1(n468), .Y(n121) );
  OAI22XL U242 ( .A0(n44), .A1(n470), .B0(n28), .B1(n469), .Y(n322) );
  OAI22XL U243 ( .A0(n44), .A1(n471), .B0(n28), .B1(n470), .Y(n323) );
  OAI22XL U244 ( .A0(n44), .A1(n472), .B0(n28), .B1(n471), .Y(n324) );
  OAI22XL U245 ( .A0(n43), .A1(n473), .B0(n27), .B1(n472), .Y(n325) );
  OAI22XL U246 ( .A0(n43), .A1(n474), .B0(n27), .B1(n473), .Y(n326) );
  OAI22XL U247 ( .A0(n43), .A1(n475), .B0(n27), .B1(n474), .Y(n327) );
  OAI22XL U248 ( .A0(n43), .A1(n476), .B0(n27), .B1(n475), .Y(n328) );
  OAI22XL U249 ( .A0(n43), .A1(n477), .B0(n27), .B1(n476), .Y(n329) );
  OAI22XL U250 ( .A0(n43), .A1(n478), .B0(n27), .B1(n477), .Y(n330) );
  OAI22XL U251 ( .A0(n43), .A1(n479), .B0(n27), .B1(n478), .Y(n331) );
  OAI22XL U252 ( .A0(n43), .A1(n480), .B0(n27), .B1(n479), .Y(n332) );
  OAI22XL U253 ( .A0(n43), .A1(n481), .B0(n27), .B1(n480), .Y(n333) );
  NOR2BX1 U254 ( .AN(n49), .B(n27), .Y(n334) );
  XNOR2X1 U255 ( .A(n11), .B(n578), .Y(n464) );
  XNOR2X1 U256 ( .A(n11), .B(n579), .Y(n465) );
  XNOR2X1 U257 ( .A(n11), .B(n580), .Y(n466) );
  XNOR2X1 U258 ( .A(n11), .B(n581), .Y(n467) );
  XNOR2X1 U259 ( .A(n11), .B(n582), .Y(n468) );
  XNOR2X1 U260 ( .A(n11), .B(n583), .Y(n469) );
  XNOR2X1 U261 ( .A(n11), .B(n584), .Y(n470) );
  XNOR2X1 U262 ( .A(n11), .B(n585), .Y(n471) );
  XNOR2X1 U263 ( .A(n11), .B(n586), .Y(n472) );
  XNOR2X1 U264 ( .A(n11), .B(n587), .Y(n473) );
  XNOR2X1 U265 ( .A(n11), .B(n588), .Y(n474) );
  XNOR2X1 U266 ( .A(n11), .B(n589), .Y(n475) );
  XNOR2X1 U267 ( .A(n11), .B(n590), .Y(n476) );
  XNOR2X1 U268 ( .A(n11), .B(n591), .Y(n477) );
  XNOR2X1 U269 ( .A(n11), .B(n592), .Y(n478) );
  XNOR2X1 U270 ( .A(n11), .B(n593), .Y(n479) );
  XNOR2X1 U271 ( .A(n11), .B(n594), .Y(n480) );
  XNOR2X1 U272 ( .A(n11), .B(n49), .Y(n481) );
  NAND2BX1 U273 ( .AN(n49), .B(n11), .Y(n482) );
  OAI22XL U274 ( .A0(n42), .A1(n623), .B0(n26), .B1(n501), .Y(n277) );
  AO21X1 U275 ( .A0(n42), .A1(n26), .B0(n483), .Y(n335) );
  OAI22XL U276 ( .A0(n42), .A1(n484), .B0(n26), .B1(n483), .Y(n107) );
  OAI22XL U277 ( .A0(n42), .A1(n485), .B0(n26), .B1(n484), .Y(n336) );
  OAI22XL U278 ( .A0(n42), .A1(n486), .B0(n26), .B1(n485), .Y(n337) );
  OAI22XL U279 ( .A0(n42), .A1(n487), .B0(n26), .B1(n486), .Y(n338) );
  OAI22XL U280 ( .A0(n42), .A1(n488), .B0(n26), .B1(n487), .Y(n339) );
  OAI22XL U281 ( .A0(n42), .A1(n489), .B0(n26), .B1(n488), .Y(n340) );
  OAI22XL U282 ( .A0(n42), .A1(n490), .B0(n26), .B1(n489), .Y(n341) );
  OAI22XL U283 ( .A0(n42), .A1(n491), .B0(n26), .B1(n490), .Y(n342) );
  OAI22XL U284 ( .A0(n41), .A1(n492), .B0(n25), .B1(n491), .Y(n343) );
  OAI22XL U285 ( .A0(n41), .A1(n493), .B0(n25), .B1(n492), .Y(n344) );
  OAI22XL U286 ( .A0(n41), .A1(n494), .B0(n25), .B1(n493), .Y(n345) );
  OAI22XL U287 ( .A0(n41), .A1(n495), .B0(n25), .B1(n494), .Y(n346) );
  OAI22XL U288 ( .A0(n41), .A1(n496), .B0(n25), .B1(n495), .Y(n347) );
  OAI22XL U289 ( .A0(n41), .A1(n497), .B0(n25), .B1(n496), .Y(n348) );
  OAI22XL U290 ( .A0(n41), .A1(n498), .B0(n25), .B1(n497), .Y(n349) );
  OAI22XL U291 ( .A0(n41), .A1(n499), .B0(n25), .B1(n498), .Y(n350) );
  OAI22XL U292 ( .A0(n41), .A1(n500), .B0(n25), .B1(n499), .Y(n351) );
  NOR2BX1 U293 ( .AN(n49), .B(n25), .Y(n352) );
  XNOR2X1 U294 ( .A(n9), .B(n578), .Y(n483) );
  XNOR2X1 U295 ( .A(n9), .B(n579), .Y(n484) );
  XNOR2X1 U296 ( .A(n9), .B(n580), .Y(n485) );
  XNOR2X1 U297 ( .A(n9), .B(n581), .Y(n486) );
  XNOR2X1 U298 ( .A(n9), .B(n582), .Y(n487) );
  XNOR2X1 U299 ( .A(n9), .B(n583), .Y(n488) );
  XNOR2X1 U300 ( .A(n9), .B(n584), .Y(n489) );
  XNOR2X1 U301 ( .A(n9), .B(n585), .Y(n490) );
  XNOR2X1 U302 ( .A(n9), .B(n586), .Y(n491) );
  XNOR2X1 U303 ( .A(n9), .B(n587), .Y(n492) );
  XNOR2X1 U304 ( .A(n9), .B(n588), .Y(n493) );
  XNOR2X1 U305 ( .A(n9), .B(n589), .Y(n494) );
  XNOR2X1 U306 ( .A(n9), .B(n590), .Y(n495) );
  XNOR2X1 U307 ( .A(n9), .B(n591), .Y(n496) );
  XNOR2X1 U308 ( .A(n9), .B(n592), .Y(n497) );
  XNOR2X1 U309 ( .A(n9), .B(n593), .Y(n498) );
  XNOR2X1 U310 ( .A(n9), .B(n594), .Y(n499) );
  XNOR2X1 U311 ( .A(n9), .B(n49), .Y(n500) );
  NAND2BX1 U312 ( .AN(n49), .B(n9), .Y(n501) );
  OAI22XL U313 ( .A0(n40), .A1(n624), .B0(n24), .B1(n520), .Y(n278) );
  AO21X1 U314 ( .A0(n40), .A1(n24), .B0(n502), .Y(n353) );
  OAI22XL U315 ( .A0(n40), .A1(n503), .B0(n24), .B1(n502), .Y(n354) );
  OAI22XL U316 ( .A0(n40), .A1(n504), .B0(n24), .B1(n503), .Y(n355) );
  OAI22XL U317 ( .A0(n40), .A1(n505), .B0(n24), .B1(n504), .Y(n356) );
  OAI22XL U318 ( .A0(n40), .A1(n506), .B0(n24), .B1(n505), .Y(n357) );
  OAI22XL U319 ( .A0(n40), .A1(n507), .B0(n24), .B1(n506), .Y(n358) );
  OAI22XL U320 ( .A0(n40), .A1(n508), .B0(n24), .B1(n507), .Y(n359) );
  OAI22XL U321 ( .A0(n40), .A1(n509), .B0(n24), .B1(n508), .Y(n360) );
  OAI22XL U322 ( .A0(n40), .A1(n510), .B0(n24), .B1(n509), .Y(n361) );
  OAI22XL U323 ( .A0(n39), .A1(n511), .B0(n23), .B1(n510), .Y(n362) );
  OAI22XL U324 ( .A0(n39), .A1(n512), .B0(n23), .B1(n511), .Y(n363) );
  OAI22XL U325 ( .A0(n39), .A1(n513), .B0(n23), .B1(n512), .Y(n364) );
  OAI22XL U326 ( .A0(n39), .A1(n514), .B0(n23), .B1(n513), .Y(n365) );
  OAI22XL U327 ( .A0(n39), .A1(n515), .B0(n23), .B1(n514), .Y(n366) );
  OAI22XL U328 ( .A0(n39), .A1(n516), .B0(n23), .B1(n515), .Y(n367) );
  OAI22XL U329 ( .A0(n39), .A1(n517), .B0(n23), .B1(n516), .Y(n368) );
  OAI22XL U330 ( .A0(n39), .A1(n518), .B0(n23), .B1(n517), .Y(n369) );
  OAI22XL U331 ( .A0(n39), .A1(n519), .B0(n23), .B1(n518), .Y(n370) );
  NOR2BX1 U332 ( .AN(n49), .B(n23), .Y(n371) );
  XNOR2X1 U333 ( .A(n7), .B(n578), .Y(n502) );
  XNOR2X1 U334 ( .A(n7), .B(n579), .Y(n503) );
  XNOR2X1 U335 ( .A(n7), .B(n580), .Y(n504) );
  XNOR2X1 U336 ( .A(n7), .B(n581), .Y(n505) );
  XNOR2X1 U337 ( .A(n7), .B(n582), .Y(n506) );
  XNOR2X1 U338 ( .A(n7), .B(n583), .Y(n507) );
  XNOR2X1 U339 ( .A(n7), .B(n584), .Y(n508) );
  XNOR2X1 U340 ( .A(n7), .B(n585), .Y(n509) );
  XNOR2X1 U341 ( .A(n7), .B(n586), .Y(n510) );
  XNOR2X1 U342 ( .A(n7), .B(n587), .Y(n511) );
  XNOR2X1 U343 ( .A(n7), .B(n588), .Y(n512) );
  XNOR2X1 U344 ( .A(n7), .B(n589), .Y(n513) );
  XNOR2X1 U345 ( .A(n7), .B(n590), .Y(n514) );
  XNOR2X1 U346 ( .A(n7), .B(n591), .Y(n515) );
  XNOR2X1 U347 ( .A(n7), .B(n592), .Y(n516) );
  XNOR2X1 U348 ( .A(n7), .B(n593), .Y(n517) );
  XNOR2X1 U349 ( .A(n7), .B(n594), .Y(n518) );
  XNOR2X1 U350 ( .A(n7), .B(n49), .Y(n519) );
  NAND2BX1 U351 ( .AN(n49), .B(n7), .Y(n520) );
  OAI22XL U352 ( .A0(n38), .A1(n625), .B0(n22), .B1(n539), .Y(n279) );
  AO21X1 U353 ( .A0(n38), .A1(n22), .B0(n521), .Y(n372) );
  OAI22XL U354 ( .A0(n38), .A1(n522), .B0(n22), .B1(n521), .Y(n139) );
  OAI22XL U355 ( .A0(n38), .A1(n523), .B0(n22), .B1(n522), .Y(n373) );
  OAI22XL U356 ( .A0(n38), .A1(n524), .B0(n22), .B1(n523), .Y(n374) );
  OAI22XL U357 ( .A0(n38), .A1(n525), .B0(n22), .B1(n524), .Y(n375) );
  OAI22XL U358 ( .A0(n38), .A1(n526), .B0(n22), .B1(n525), .Y(n376) );
  OAI22XL U359 ( .A0(n38), .A1(n527), .B0(n22), .B1(n526), .Y(n377) );
  OAI22XL U360 ( .A0(n38), .A1(n528), .B0(n22), .B1(n527), .Y(n378) );
  OAI22XL U361 ( .A0(n38), .A1(n529), .B0(n22), .B1(n528), .Y(n379) );
  OAI22XL U362 ( .A0(n37), .A1(n530), .B0(n21), .B1(n529), .Y(n380) );
  OAI22XL U363 ( .A0(n37), .A1(n531), .B0(n21), .B1(n530), .Y(n381) );
  OAI22XL U364 ( .A0(n37), .A1(n532), .B0(n21), .B1(n531), .Y(n382) );
  OAI22XL U365 ( .A0(n37), .A1(n533), .B0(n21), .B1(n532), .Y(n383) );
  OAI22XL U366 ( .A0(n37), .A1(n534), .B0(n21), .B1(n533), .Y(n384) );
  OAI22XL U367 ( .A0(n37), .A1(n535), .B0(n21), .B1(n534), .Y(n385) );
  OAI22XL U368 ( .A0(n37), .A1(n536), .B0(n21), .B1(n535), .Y(n386) );
  OAI22XL U369 ( .A0(n37), .A1(n537), .B0(n21), .B1(n536), .Y(n387) );
  OAI22XL U370 ( .A0(n37), .A1(n538), .B0(n21), .B1(n537), .Y(n388) );
  NOR2BX1 U371 ( .AN(n49), .B(n21), .Y(n389) );
  XNOR2X1 U372 ( .A(n5), .B(n578), .Y(n521) );
  XNOR2X1 U373 ( .A(n5), .B(n579), .Y(n522) );
  XNOR2X1 U374 ( .A(n5), .B(n580), .Y(n523) );
  XNOR2X1 U375 ( .A(n5), .B(n581), .Y(n524) );
  XNOR2X1 U376 ( .A(n5), .B(n582), .Y(n525) );
  XNOR2X1 U377 ( .A(n5), .B(n583), .Y(n526) );
  XNOR2X1 U378 ( .A(n5), .B(n584), .Y(n527) );
  XNOR2X1 U379 ( .A(n5), .B(n585), .Y(n528) );
  XNOR2X1 U380 ( .A(n5), .B(n586), .Y(n529) );
  XNOR2X1 U381 ( .A(n5), .B(n587), .Y(n530) );
  XNOR2X1 U382 ( .A(n5), .B(n588), .Y(n531) );
  XNOR2X1 U383 ( .A(n5), .B(n589), .Y(n532) );
  XNOR2X1 U384 ( .A(n5), .B(n590), .Y(n533) );
  XNOR2X1 U385 ( .A(n5), .B(n591), .Y(n534) );
  XNOR2X1 U386 ( .A(n5), .B(n592), .Y(n535) );
  XNOR2X1 U387 ( .A(n5), .B(n593), .Y(n536) );
  XNOR2X1 U388 ( .A(n5), .B(n594), .Y(n537) );
  XNOR2X1 U389 ( .A(n5), .B(n49), .Y(n538) );
  NAND2BX1 U390 ( .AN(n49), .B(n5), .Y(n539) );
  OAI22XL U391 ( .A0(n36), .A1(n626), .B0(n20), .B1(n558), .Y(n280) );
  AO21X1 U392 ( .A0(n36), .A1(n20), .B0(n540), .Y(n390) );
  OAI22XL U393 ( .A0(n36), .A1(n541), .B0(n20), .B1(n540), .Y(n159) );
  OAI22XL U394 ( .A0(n36), .A1(n542), .B0(n20), .B1(n541), .Y(n391) );
  OAI22XL U395 ( .A0(n36), .A1(n543), .B0(n20), .B1(n542), .Y(n392) );
  OAI22XL U396 ( .A0(n36), .A1(n544), .B0(n20), .B1(n543), .Y(n393) );
  OAI22XL U397 ( .A0(n36), .A1(n545), .B0(n20), .B1(n544), .Y(n394) );
  OAI22XL U398 ( .A0(n36), .A1(n546), .B0(n20), .B1(n545), .Y(n395) );
  OAI22XL U399 ( .A0(n36), .A1(n547), .B0(n20), .B1(n546), .Y(n396) );
  OAI22XL U400 ( .A0(n36), .A1(n548), .B0(n20), .B1(n547), .Y(n397) );
  OAI22XL U401 ( .A0(n35), .A1(n549), .B0(n19), .B1(n548), .Y(n398) );
  OAI22XL U402 ( .A0(n35), .A1(n550), .B0(n19), .B1(n549), .Y(n399) );
  OAI22XL U403 ( .A0(n35), .A1(n551), .B0(n19), .B1(n550), .Y(n400) );
  OAI22XL U404 ( .A0(n35), .A1(n552), .B0(n19), .B1(n551), .Y(n401) );
  OAI22XL U405 ( .A0(n35), .A1(n553), .B0(n19), .B1(n552), .Y(n402) );
  OAI22XL U406 ( .A0(n35), .A1(n554), .B0(n19), .B1(n553), .Y(n403) );
  OAI22XL U407 ( .A0(n35), .A1(n555), .B0(n19), .B1(n554), .Y(n404) );
  OAI22XL U408 ( .A0(n35), .A1(n556), .B0(n19), .B1(n555), .Y(n405) );
  OAI22XL U409 ( .A0(n35), .A1(n557), .B0(n19), .B1(n556), .Y(n406) );
  NOR2BX1 U410 ( .AN(n49), .B(n19), .Y(n407) );
  XNOR2X1 U411 ( .A(n3), .B(n578), .Y(n540) );
  XNOR2X1 U412 ( .A(n3), .B(n579), .Y(n541) );
  XNOR2X1 U413 ( .A(n3), .B(n580), .Y(n542) );
  XNOR2X1 U414 ( .A(n3), .B(n581), .Y(n543) );
  XNOR2X1 U415 ( .A(n3), .B(n582), .Y(n544) );
  XNOR2X1 U416 ( .A(n3), .B(n583), .Y(n545) );
  XNOR2X1 U417 ( .A(n3), .B(n584), .Y(n546) );
  XNOR2X1 U418 ( .A(n3), .B(n585), .Y(n547) );
  XNOR2X1 U419 ( .A(n3), .B(n586), .Y(n548) );
  XNOR2X1 U420 ( .A(n3), .B(n587), .Y(n549) );
  XNOR2X1 U421 ( .A(n3), .B(n588), .Y(n550) );
  XNOR2X1 U422 ( .A(n3), .B(n589), .Y(n551) );
  XNOR2X1 U423 ( .A(n3), .B(n590), .Y(n552) );
  XNOR2X1 U424 ( .A(n3), .B(n591), .Y(n553) );
  XNOR2X1 U425 ( .A(n3), .B(n592), .Y(n554) );
  XNOR2X1 U426 ( .A(n3), .B(n593), .Y(n555) );
  XNOR2X1 U427 ( .A(n3), .B(n594), .Y(n556) );
  XNOR2X1 U428 ( .A(n3), .B(n49), .Y(n557) );
  NAND2BX1 U429 ( .AN(n49), .B(n3), .Y(n558) );
  OAI22XL U430 ( .A0(n34), .A1(n627), .B0(n577), .B1(n18), .Y(n281) );
  AO21X1 U431 ( .A0(n34), .A1(n18), .B0(n559), .Y(n408) );
  OAI22XL U432 ( .A0(n34), .A1(n560), .B0(n559), .B1(n18), .Y(n409) );
  OAI22XL U433 ( .A0(n34), .A1(n561), .B0(n560), .B1(n18), .Y(n410) );
  OAI22XL U434 ( .A0(n34), .A1(n562), .B0(n561), .B1(n18), .Y(n411) );
  OAI22XL U435 ( .A0(n34), .A1(n563), .B0(n562), .B1(n18), .Y(n412) );
  OAI22XL U436 ( .A0(n34), .A1(n564), .B0(n563), .B1(n18), .Y(n413) );
  OAI22XL U437 ( .A0(n34), .A1(n565), .B0(n564), .B1(n18), .Y(n414) );
  OAI22XL U438 ( .A0(n34), .A1(n566), .B0(n565), .B1(n18), .Y(n415) );
  OAI22XL U439 ( .A0(n34), .A1(n567), .B0(n566), .B1(n18), .Y(n416) );
  OAI22XL U440 ( .A0(n33), .A1(n568), .B0(n567), .B1(n17), .Y(n417) );
  OAI22XL U441 ( .A0(n33), .A1(n569), .B0(n568), .B1(n17), .Y(n418) );
  OAI22XL U442 ( .A0(n33), .A1(n570), .B0(n569), .B1(n17), .Y(n419) );
  OAI22XL U443 ( .A0(n33), .A1(n571), .B0(n570), .B1(n17), .Y(n420) );
  OAI22XL U444 ( .A0(n33), .A1(n572), .B0(n571), .B1(n17), .Y(n421) );
  OAI22XL U445 ( .A0(n33), .A1(n573), .B0(n572), .B1(n17), .Y(n422) );
  OAI22XL U446 ( .A0(n33), .A1(n574), .B0(n573), .B1(n17), .Y(n423) );
  OAI22XL U447 ( .A0(n33), .A1(n575), .B0(n574), .B1(n17), .Y(n424) );
  OAI22XL U448 ( .A0(n33), .A1(n576), .B0(n575), .B1(n17), .Y(n425) );
  NOR2BX1 U449 ( .AN(n49), .B(n17), .Y(product_0_) );
  XNOR2X1 U450 ( .A(n1), .B(n578), .Y(n559) );
  XNOR2X1 U451 ( .A(n1), .B(n579), .Y(n560) );
  XNOR2X1 U452 ( .A(n1), .B(n580), .Y(n561) );
  XNOR2X1 U453 ( .A(n1), .B(n581), .Y(n562) );
  XNOR2X1 U454 ( .A(n1), .B(n582), .Y(n563) );
  XNOR2X1 U455 ( .A(n1), .B(n583), .Y(n564) );
  XNOR2X1 U456 ( .A(n1), .B(n584), .Y(n565) );
  XNOR2X1 U457 ( .A(n1), .B(n585), .Y(n566) );
  XNOR2X1 U458 ( .A(n1), .B(n586), .Y(n567) );
  XNOR2X1 U459 ( .A(n1), .B(n587), .Y(n568) );
  XNOR2X1 U460 ( .A(n1), .B(n588), .Y(n569) );
  XNOR2X1 U461 ( .A(n1), .B(n589), .Y(n570) );
  XNOR2X1 U462 ( .A(n1), .B(n590), .Y(n571) );
  XNOR2X1 U463 ( .A(n1), .B(n591), .Y(n572) );
  XNOR2X1 U464 ( .A(n1), .B(n592), .Y(n573) );
  XNOR2X1 U465 ( .A(n1), .B(n593), .Y(n574) );
  XNOR2X1 U466 ( .A(n1), .B(n594), .Y(n575) );
  XNOR2X1 U467 ( .A(n1), .B(n49), .Y(n576) );
  NAND2BX1 U468 ( .AN(n49), .B(n1), .Y(n577) );
  CLKINVX1 U486 ( .A(n15), .Y(n620) );
  CLKINVX1 U487 ( .A(n13), .Y(n621) );
  CLKINVX1 U488 ( .A(n11), .Y(n622) );
  CLKINVX1 U489 ( .A(n9), .Y(n623) );
  CLKINVX1 U490 ( .A(n7), .Y(n624) );
  CLKINVX1 U491 ( .A(n5), .Y(n625) );
  CLKINVX1 U492 ( .A(n3), .Y(n626) );
  CLKINVX1 U493 ( .A(n1), .Y(n627) );
  NAND2X1 U494 ( .A(n596), .B(n612), .Y(n604) );
  XOR2X1 U495 ( .A(a[14]), .B(a[15]), .Y(n596) );
  XNOR2X1 U496 ( .A(a[14]), .B(a[13]), .Y(n612) );
  NAND2X1 U497 ( .A(n597), .B(n613), .Y(n605) );
  XOR2X1 U498 ( .A(a[12]), .B(a[13]), .Y(n597) );
  XNOR2X1 U499 ( .A(a[12]), .B(a[11]), .Y(n613) );
  NAND2X1 U500 ( .A(n598), .B(n614), .Y(n606) );
  XOR2X1 U501 ( .A(a[10]), .B(a[11]), .Y(n598) );
  XNOR2X1 U502 ( .A(a[10]), .B(a[9]), .Y(n614) );
  NAND2X1 U503 ( .A(n599), .B(n615), .Y(n607) );
  XOR2X1 U504 ( .A(a[8]), .B(a[9]), .Y(n599) );
  XNOR2X1 U505 ( .A(a[8]), .B(a[7]), .Y(n615) );
  NAND2X1 U506 ( .A(n600), .B(n616), .Y(n608) );
  XOR2X1 U507 ( .A(a[6]), .B(a[7]), .Y(n600) );
  XNOR2X1 U508 ( .A(a[6]), .B(a[5]), .Y(n616) );
  NAND2X1 U509 ( .A(n601), .B(n617), .Y(n609) );
  XOR2X1 U510 ( .A(a[4]), .B(a[5]), .Y(n601) );
  XNOR2X1 U511 ( .A(a[4]), .B(a[3]), .Y(n617) );
  NAND2X1 U512 ( .A(n602), .B(n618), .Y(n610) );
  XOR2X1 U513 ( .A(a[2]), .B(a[3]), .Y(n602) );
  XNOR2X1 U514 ( .A(a[2]), .B(a[1]), .Y(n618) );
  NAND2X1 U515 ( .A(n603), .B(n619), .Y(n611) );
  XOR2X1 U516 ( .A(a[0]), .B(a[1]), .Y(n603) );
  CLKINVX1 U517 ( .A(a[0]), .Y(n619) );
  OA22X1 U520 ( .A0(n48), .A1(n427), .B0(n32), .B1(n426), .Y(n697) );
  CLKBUFX3 U521 ( .A(b_2_), .Y(n593) );
  CLKBUFX3 U522 ( .A(b_0_), .Y(n49) );
  CLKBUFX3 U523 ( .A(b_3_), .Y(n592) );
  CLKBUFX3 U524 ( .A(b_9_), .Y(n586) );
  CLKBUFX3 U525 ( .A(b_17_), .Y(n578) );
  CLKBUFX3 U526 ( .A(b_4_), .Y(n591) );
  CLKBUFX3 U527 ( .A(b_5_), .Y(n590) );
  CLKBUFX3 U528 ( .A(b_6_), .Y(n589) );
  CLKBUFX3 U529 ( .A(b_10_), .Y(n585) );
  CLKBUFX3 U530 ( .A(b_15_), .Y(n580) );
  CLKBUFX3 U531 ( .A(b_7_), .Y(n588) );
  CLKBUFX3 U532 ( .A(b_14_), .Y(n581) );
  CLKBUFX3 U533 ( .A(b_1_), .Y(n594) );
  CLKBUFX3 U534 ( .A(b_16_), .Y(n579) );
  CLKBUFX3 U535 ( .A(n618), .Y(n19) );
  CLKBUFX3 U536 ( .A(n617), .Y(n21) );
  CLKBUFX3 U537 ( .A(n616), .Y(n23) );
  CLKBUFX3 U538 ( .A(n615), .Y(n25) );
  CLKBUFX3 U539 ( .A(n614), .Y(n27) );
  CLKBUFX3 U540 ( .A(n613), .Y(n29) );
  CLKBUFX3 U541 ( .A(n612), .Y(n31) );
  CLKBUFX3 U542 ( .A(n618), .Y(n20) );
  CLKBUFX3 U543 ( .A(n617), .Y(n22) );
  CLKBUFX3 U544 ( .A(n615), .Y(n26) );
  CLKBUFX3 U545 ( .A(n616), .Y(n24) );
  CLKBUFX3 U546 ( .A(n613), .Y(n30) );
  CLKBUFX3 U547 ( .A(n614), .Y(n28) );
  CLKBUFX3 U548 ( .A(b_13_), .Y(n582) );
  CLKBUFX3 U549 ( .A(b_8_), .Y(n587) );
  CLKBUFX3 U550 ( .A(n612), .Y(n32) );
  CLKBUFX3 U551 ( .A(b_11_), .Y(n584) );
  CLKBUFX3 U552 ( .A(b_12_), .Y(n583) );
  CLKBUFX3 U553 ( .A(n610), .Y(n36) );
  CLKBUFX3 U554 ( .A(n609), .Y(n38) );
  CLKBUFX3 U555 ( .A(n607), .Y(n42) );
  CLKBUFX3 U556 ( .A(n608), .Y(n40) );
  CLKBUFX3 U557 ( .A(n605), .Y(n46) );
  CLKBUFX3 U558 ( .A(n606), .Y(n44) );
  CLKBUFX3 U559 ( .A(n611), .Y(n34) );
  CLKBUFX3 U560 ( .A(n610), .Y(n35) );
  CLKBUFX3 U561 ( .A(n609), .Y(n37) );
  CLKBUFX3 U562 ( .A(n608), .Y(n39) );
  CLKBUFX3 U563 ( .A(n607), .Y(n41) );
  CLKBUFX3 U564 ( .A(n606), .Y(n43) );
  CLKBUFX3 U565 ( .A(n605), .Y(n45) );
  CLKBUFX3 U566 ( .A(n604), .Y(n47) );
  CLKBUFX3 U567 ( .A(n604), .Y(n48) );
  CLKBUFX3 U568 ( .A(n611), .Y(n33) );
  CLKBUFX3 U569 ( .A(n619), .Y(n17) );
  CLKBUFX3 U570 ( .A(n619), .Y(n18) );
  CLKBUFX3 U571 ( .A(a[1]), .Y(n1) );
  CLKBUFX3 U572 ( .A(a[3]), .Y(n3) );
  CLKBUFX3 U573 ( .A(a[5]), .Y(n5) );
  CLKBUFX3 U574 ( .A(a[7]), .Y(n7) );
  CLKBUFX3 U575 ( .A(a[9]), .Y(n9) );
  CLKBUFX3 U576 ( .A(a[11]), .Y(n11) );
  CLKBUFX3 U577 ( .A(a[13]), .Y(n13) );
  CLKBUFX3 U578 ( .A(a[15]), .Y(n15) );
endmodule


module FAS_DW_mult_tc_28 ( a, b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, 
        b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input [15:0] a;
  input b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_, b_8_, b_7_,
         b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n3, n5, n7, n9, n11, n13, n15, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600;

  XOR2X1 U51 ( .A(n52), .B(n51), .Y(product_31_) );
  XOR2X1 U52 ( .A(n272), .B(n82), .Y(n51) );
  ADDFXL U53 ( .A(n84), .B(n83), .CI(n53), .CO(n52), .S(product_30_) );
  ADDFXL U54 ( .A(n85), .B(n86), .CI(n54), .CO(n53), .S(product_29_) );
  ADDFXL U55 ( .A(n91), .B(n87), .CI(n55), .CO(n54), .S(product_28_) );
  ADDFXL U56 ( .A(n94), .B(n92), .CI(n56), .CO(n55), .S(product_27_) );
  ADDFXL U57 ( .A(n95), .B(n99), .CI(n57), .CO(n56), .S(product_26_) );
  ADDFXL U58 ( .A(n100), .B(n104), .CI(n58), .CO(n57), .S(product_25_) );
  ADDFXL U59 ( .A(n105), .B(n111), .CI(n59), .CO(n58), .S(product_24_) );
  ADDFXL U60 ( .A(n112), .B(n117), .CI(n60), .CO(n59), .S(product_23_) );
  ADDFXL U61 ( .A(n118), .B(n125), .CI(n61), .CO(n60), .S(product_22_) );
  ADDFXL U62 ( .A(n133), .B(n126), .CI(n62), .CO(n61), .S(product_21_) );
  ADDFXL U63 ( .A(n143), .B(n134), .CI(n63), .CO(n62), .S(product_20_) );
  ADDFXL U64 ( .A(n144), .B(n152), .CI(n64), .CO(n63), .S(product_19_) );
  ADDFXL U65 ( .A(n153), .B(n163), .CI(n65), .CO(n64), .S(product_18_) );
  ADDFXL U66 ( .A(n164), .B(n174), .CI(n66), .CO(n65), .S(product_17_) );
  ADDFXL U67 ( .A(n175), .B(n185), .CI(n67), .CO(n66), .S(product_16_) );
  ADDFXL U68 ( .A(n186), .B(n196), .CI(n68), .CO(n67), .S(product_15_) );
  ADDFXL U69 ( .A(n197), .B(n205), .CI(n69), .CO(n68), .S(product_14_) );
  ADDFXL U70 ( .A(n206), .B(n215), .CI(n70), .CO(n69), .S(product_13_) );
  ADDFXL U71 ( .A(n216), .B(n223), .CI(n71), .CO(n70), .S(product_12_) );
  ADDFXL U72 ( .A(n224), .B(n231), .CI(n72), .CO(n71), .S(product_11_) );
  ADDFXL U73 ( .A(n232), .B(n237), .CI(n73), .CO(n72), .S(product_10_) );
  ADDFXL U74 ( .A(n238), .B(n244), .CI(n74), .CO(n73), .S(product_9_) );
  ADDFXL U75 ( .A(n245), .B(n249), .CI(n75), .CO(n74), .S(product_8_) );
  ADDFXL U76 ( .A(n250), .B(n254), .CI(n76), .CO(n75), .S(product_7_) );
  ADDFXL U77 ( .A(n255), .B(n256), .CI(n77), .CO(n76), .S(product_6_) );
  ADDFXL U78 ( .A(n257), .B(n260), .CI(n78), .CO(n77), .S(product_5_) );
  ADDFXL U79 ( .A(n261), .B(n262), .CI(n79), .CO(n78), .S(product_4_) );
  ADDFXL U80 ( .A(n263), .B(n389), .CI(n80), .CO(n79), .S(product_3_) );
  ADDFXL U81 ( .A(n406), .B(n390), .CI(n81), .CO(n80), .S(product_2_) );
  ADDHXL U82 ( .A(n271), .B(n407), .CO(n81), .S(product_1_) );
  CLKINVX1 U83 ( .A(n82), .Y(n83) );
  ADDFXL U84 ( .A(n273), .B(n88), .CI(n289), .CO(n84), .S(n85) );
  ADDFXL U85 ( .A(n89), .B(n274), .CI(n90), .CO(n86), .S(n87) );
  CLKINVX1 U86 ( .A(n88), .Y(n89) );
  CMPR42X1 U87 ( .A(n96), .B(n275), .C(n290), .D(n306), .ICI(n93), .S(n92), 
        .ICO(n90), .CO(n91) );
  CMPR42X1 U88 ( .A(n291), .B(n276), .C(n97), .D(n101), .ICI(n98), .S(n95), 
        .ICO(n93), .CO(n94) );
  CLKINVX1 U89 ( .A(n96), .Y(n97) );
  CMPR42X1 U90 ( .A(n307), .B(n292), .C(n106), .D(n102), .ICI(n103), .S(n100), 
        .ICO(n98), .CO(n99) );
  ADDFXL U91 ( .A(n108), .B(n277), .CI(n322), .CO(n101), .S(n102) );
  CMPR42X1 U92 ( .A(n308), .B(n113), .C(n107), .D(n114), .ICI(n110), .S(n105), 
        .ICO(n103), .CO(n104) );
  ADDFXL U93 ( .A(n293), .B(n278), .CI(n109), .CO(n106), .S(n107) );
  CLKINVX1 U94 ( .A(n108), .Y(n109) );
  CMPR42X1 U95 ( .A(n309), .B(n294), .C(n120), .D(n115), .ICI(n116), .S(n112), 
        .ICO(n110), .CO(n111) );
  CMPR42X1 U96 ( .A(n279), .B(n122), .C(n323), .D(n339), .ICI(n119), .S(n115), 
        .ICO(n113), .CO(n114) );
  CMPR42X1 U97 ( .A(n280), .B(n130), .C(n128), .D(n121), .ICI(n124), .S(n118), 
        .ICO(n116), .CO(n117) );
  CMPR42X1 U98 ( .A(n295), .B(n340), .C(n324), .D(n123), .ICI(n127), .S(n121), 
        .ICO(n119), .CO(n120) );
  CLKINVX1 U99 ( .A(n122), .Y(n123) );
  CMPR42X1 U100 ( .A(n138), .B(n131), .C(n136), .D(n129), .ICI(n132), .S(n126), 
        .ICO(n124), .CO(n125) );
  CMPR42X1 U101 ( .A(n296), .B(n325), .C(n310), .D(n140), .ICI(n135), .S(n129), 
        .ICO(n127), .CO(n128) );
  ADDFXL U102 ( .A(n341), .B(n281), .CI(n357), .CO(n130), .S(n131) );
  CMPR42X1 U103 ( .A(n139), .B(n149), .C(n146), .D(n137), .ICI(n142), .S(n134), 
        .ICO(n132), .CO(n133) );
  CMPR42X1 U104 ( .A(n342), .B(n311), .C(n326), .D(n145), .ICI(n148), .S(n137), 
        .ICO(n135), .CO(n136) );
  ADDFXL U105 ( .A(n282), .B(n297), .CI(n141), .CO(n138), .S(n139) );
  CLKINVX1 U106 ( .A(n140), .Y(n141) );
  CMPR42X1 U107 ( .A(n158), .B(n155), .C(n147), .D(n150), .ICI(n151), .S(n144), 
        .ICO(n142), .CO(n143) );
  CMPR42X1 U108 ( .A(n298), .B(n327), .C(n312), .D(n160), .ICI(n154), .S(n147), 
        .ICO(n145), .CO(n146) );
  CMPR42X1 U109 ( .A(n283), .B(n358), .C(n343), .D(n374), .ICI(n157), .S(n150), 
        .ICO(n148), .CO(n149) );
  CMPR42X1 U110 ( .A(n169), .B(n166), .C(n156), .D(n159), .ICI(n162), .S(n153), 
        .ICO(n151), .CO(n152) );
  CMPR42X1 U111 ( .A(n313), .B(n344), .C(n328), .D(n284), .ICI(n165), .S(n156), 
        .ICO(n154), .CO(n155) );
  CMPR42X1 U112 ( .A(n299), .B(n359), .C(n161), .D(n171), .ICI(n168), .S(n159), 
        .ICO(n157), .CO(n158) );
  CLKINVX1 U113 ( .A(n160), .Y(n161) );
  CMPR42X1 U114 ( .A(n180), .B(n177), .C(n167), .D(n170), .ICI(n173), .S(n164), 
        .ICO(n162), .CO(n163) );
  CMPR42X1 U115 ( .A(n285), .B(n360), .C(n329), .D(n182), .ICI(n176), .S(n167), 
        .ICO(n165), .CO(n166) );
  CMPR42X1 U116 ( .A(n314), .B(n375), .C(n391), .D(n172), .ICI(n179), .S(n170), 
        .ICO(n168), .CO(n169) );
  XNOR2X1 U117 ( .A(n345), .B(n300), .Y(n172) );
  OR2X1 U118 ( .A(n345), .B(n300), .Y(n171) );
  CMPR42X1 U119 ( .A(n191), .B(n188), .C(n181), .D(n178), .ICI(n184), .S(n175), 
        .ICO(n173), .CO(n174) );
  CMPR42X1 U120 ( .A(n301), .B(n315), .C(n346), .D(n183), .ICI(n190), .S(n178), 
        .ICO(n176), .CO(n177) );
  CMPR42X1 U121 ( .A(n330), .B(n376), .C(n361), .D(n193), .ICI(n187), .S(n181), 
        .ICO(n179), .CO(n180) );
  ADDHXL U122 ( .A(n392), .B(n286), .CO(n182), .S(n183) );
  CMPR42X1 U123 ( .A(n202), .B(n199), .C(n192), .D(n189), .ICI(n195), .S(n186), 
        .ICO(n184), .CO(n185) );
  CMPR42X1 U124 ( .A(n302), .B(n316), .C(n331), .D(n201), .ICI(n194), .S(n189), 
        .ICO(n187), .CO(n188) );
  CMPR42X1 U125 ( .A(n264), .B(n287), .C(n377), .D(n347), .ICI(n198), .S(n192), 
        .ICO(n190), .CO(n191) );
  ADDHXL U126 ( .A(n393), .B(n362), .CO(n193), .S(n194) );
  CMPR42X1 U127 ( .A(n210), .B(n203), .C(n208), .D(n200), .ICI(n204), .S(n197), 
        .ICO(n195), .CO(n196) );
  CMPR42X1 U128 ( .A(n378), .B(n332), .C(n348), .D(n363), .ICI(n212), .S(n200), 
        .ICO(n198), .CO(n199) );
  CMPR42X1 U129 ( .A(n288), .B(n394), .C(n303), .D(n317), .ICI(n207), .S(n203), 
        .ICO(n201), .CO(n202) );
  CMPR42X1 U130 ( .A(n220), .B(n211), .C(n218), .D(n209), .ICI(n214), .S(n206), 
        .ICO(n204), .CO(n205) );
  CMPR42X1 U131 ( .A(n318), .B(n349), .C(n333), .D(n304), .ICI(n217), .S(n209), 
        .ICO(n207), .CO(n208) );
  ADDFXL U132 ( .A(n379), .B(n265), .CI(n213), .CO(n210), .S(n211) );
  ADDHXL U133 ( .A(n395), .B(n364), .CO(n212), .S(n213) );
  CMPR42X1 U134 ( .A(n350), .B(n225), .C(n226), .D(n219), .ICI(n222), .S(n216), 
        .ICO(n214), .CO(n215) );
  CMPR42X1 U135 ( .A(n380), .B(n334), .C(n365), .D(n228), .ICI(n221), .S(n219), 
        .ICO(n217), .CO(n218) );
  ADDFXL U136 ( .A(n396), .B(n305), .CI(n319), .CO(n220), .S(n221) );
  CMPR42X1 U137 ( .A(n351), .B(n233), .C(n234), .D(n227), .ICI(n230), .S(n224), 
        .ICO(n222), .CO(n223) );
  CMPR42X1 U138 ( .A(n266), .B(n320), .C(n381), .D(n335), .ICI(n229), .S(n227), 
        .ICO(n225), .CO(n226) );
  ADDHXL U139 ( .A(n397), .B(n366), .CO(n228), .S(n229) );
  CMPR42X1 U140 ( .A(n382), .B(n367), .C(n239), .D(n236), .ICI(n235), .S(n232), 
        .ICO(n230), .CO(n231) );
  CMPR42X1 U141 ( .A(n321), .B(n398), .C(n336), .D(n352), .ICI(n241), .S(n235), 
        .ICO(n233), .CO(n234) );
  CMPR42X1 U142 ( .A(n383), .B(n353), .C(n243), .D(n246), .ICI(n240), .S(n238), 
        .ICO(n236), .CO(n237) );
  ADDFXL U143 ( .A(n337), .B(n267), .CI(n242), .CO(n239), .S(n240) );
  ADDHXL U144 ( .A(n399), .B(n368), .CO(n241), .S(n242) );
  CMPR42X1 U145 ( .A(n384), .B(n369), .C(n251), .D(n248), .ICI(n247), .S(n245), 
        .ICO(n243), .CO(n244) );
  ADDFXL U146 ( .A(n400), .B(n338), .CI(n354), .CO(n246), .S(n247) );
  CMPR42X1 U147 ( .A(n268), .B(n355), .C(n385), .D(n253), .ICI(n252), .S(n250), 
        .ICO(n248), .CO(n249) );
  ADDHXL U148 ( .A(n401), .B(n370), .CO(n251), .S(n252) );
  CMPR42X1 U149 ( .A(n356), .B(n402), .C(n371), .D(n386), .ICI(n258), .S(n255), 
        .ICO(n253), .CO(n254) );
  ADDFXL U150 ( .A(n387), .B(n269), .CI(n259), .CO(n256), .S(n257) );
  ADDHXL U151 ( .A(n403), .B(n372), .CO(n258), .S(n259) );
  ADDFXL U152 ( .A(n404), .B(n373), .CI(n388), .CO(n260), .S(n261) );
  ADDHXL U153 ( .A(n405), .B(n270), .CO(n262), .S(n263) );
  OAI22XL U154 ( .A0(n48), .A1(n593), .B0(n32), .B1(n425), .Y(n264) );
  AO21X1 U155 ( .A0(n48), .A1(n32), .B0(n408), .Y(n272) );
  OAI22XL U156 ( .A0(n48), .A1(n409), .B0(n32), .B1(n408), .Y(n82) );
  OAI22XL U157 ( .A0(n48), .A1(n410), .B0(n32), .B1(n409), .Y(n273) );
  OAI22XL U158 ( .A0(n48), .A1(n411), .B0(n32), .B1(n410), .Y(n274) );
  OAI22XL U159 ( .A0(n48), .A1(n412), .B0(n32), .B1(n411), .Y(n275) );
  OAI22XL U160 ( .A0(n48), .A1(n413), .B0(n32), .B1(n412), .Y(n276) );
  OAI22XL U161 ( .A0(n48), .A1(n414), .B0(n32), .B1(n413), .Y(n277) );
  OAI22XL U162 ( .A0(n48), .A1(n415), .B0(n32), .B1(n414), .Y(n278) );
  OAI22XL U163 ( .A0(n47), .A1(n416), .B0(n32), .B1(n415), .Y(n279) );
  OAI22XL U164 ( .A0(n47), .A1(n417), .B0(n31), .B1(n416), .Y(n280) );
  OAI22XL U165 ( .A0(n47), .A1(n418), .B0(n31), .B1(n417), .Y(n281) );
  OAI22XL U166 ( .A0(n47), .A1(n419), .B0(n31), .B1(n418), .Y(n282) );
  OAI22XL U167 ( .A0(n47), .A1(n420), .B0(n31), .B1(n419), .Y(n283) );
  OAI22XL U168 ( .A0(n47), .A1(n421), .B0(n31), .B1(n420), .Y(n284) );
  OAI22XL U169 ( .A0(n47), .A1(n422), .B0(n31), .B1(n421), .Y(n285) );
  OAI22XL U170 ( .A0(n47), .A1(n423), .B0(n31), .B1(n422), .Y(n286) );
  OAI22XL U171 ( .A0(n47), .A1(n424), .B0(n31), .B1(n423), .Y(n287) );
  NOR2BX1 U172 ( .AN(n49), .B(n31), .Y(n288) );
  XNOR2X1 U173 ( .A(n15), .B(n552), .Y(n408) );
  XNOR2X1 U174 ( .A(n15), .B(n553), .Y(n409) );
  XNOR2X1 U175 ( .A(n15), .B(n554), .Y(n410) );
  XNOR2X1 U176 ( .A(n15), .B(n555), .Y(n411) );
  XNOR2X1 U177 ( .A(n15), .B(n556), .Y(n412) );
  XNOR2X1 U178 ( .A(n15), .B(n557), .Y(n413) );
  XNOR2X1 U179 ( .A(n15), .B(n558), .Y(n414) );
  XNOR2X1 U180 ( .A(n15), .B(n559), .Y(n415) );
  XNOR2X1 U181 ( .A(n15), .B(n560), .Y(n416) );
  XNOR2X1 U182 ( .A(n15), .B(n561), .Y(n417) );
  XNOR2X1 U183 ( .A(n15), .B(n562), .Y(n418) );
  XNOR2X1 U184 ( .A(n15), .B(n563), .Y(n419) );
  XNOR2X1 U185 ( .A(n15), .B(n564), .Y(n420) );
  XNOR2X1 U186 ( .A(n15), .B(n565), .Y(n421) );
  XNOR2X1 U187 ( .A(n15), .B(n566), .Y(n422) );
  XNOR2X1 U188 ( .A(n15), .B(n567), .Y(n423) );
  XNOR2X1 U189 ( .A(n15), .B(n49), .Y(n424) );
  NAND2BX1 U190 ( .AN(n49), .B(n15), .Y(n425) );
  OAI22XL U191 ( .A0(n46), .A1(n594), .B0(n30), .B1(n443), .Y(n265) );
  AO21X1 U192 ( .A0(n46), .A1(n30), .B0(n426), .Y(n289) );
  OAI22XL U193 ( .A0(n46), .A1(n427), .B0(n30), .B1(n426), .Y(n88) );
  OAI22XL U194 ( .A0(n46), .A1(n428), .B0(n30), .B1(n427), .Y(n290) );
  OAI22XL U195 ( .A0(n46), .A1(n429), .B0(n30), .B1(n428), .Y(n291) );
  OAI22XL U196 ( .A0(n46), .A1(n430), .B0(n30), .B1(n429), .Y(n292) );
  OAI22XL U197 ( .A0(n46), .A1(n431), .B0(n30), .B1(n430), .Y(n293) );
  OAI22XL U198 ( .A0(n46), .A1(n432), .B0(n30), .B1(n431), .Y(n294) );
  OAI22XL U199 ( .A0(n46), .A1(n433), .B0(n30), .B1(n432), .Y(n295) );
  OAI22XL U200 ( .A0(n45), .A1(n434), .B0(n30), .B1(n433), .Y(n296) );
  OAI22XL U201 ( .A0(n45), .A1(n435), .B0(n29), .B1(n434), .Y(n297) );
  OAI22XL U202 ( .A0(n45), .A1(n436), .B0(n29), .B1(n435), .Y(n298) );
  OAI22XL U203 ( .A0(n45), .A1(n437), .B0(n29), .B1(n436), .Y(n299) );
  OAI22XL U204 ( .A0(n45), .A1(n438), .B0(n29), .B1(n437), .Y(n300) );
  OAI22XL U205 ( .A0(n45), .A1(n439), .B0(n29), .B1(n438), .Y(n301) );
  OAI22XL U206 ( .A0(n45), .A1(n440), .B0(n29), .B1(n439), .Y(n302) );
  OAI22XL U207 ( .A0(n45), .A1(n441), .B0(n29), .B1(n440), .Y(n303) );
  OAI22XL U208 ( .A0(n45), .A1(n442), .B0(n29), .B1(n441), .Y(n304) );
  NOR2BX1 U209 ( .AN(n49), .B(n29), .Y(n305) );
  XNOR2X1 U210 ( .A(n13), .B(n552), .Y(n426) );
  XNOR2X1 U211 ( .A(n13), .B(n553), .Y(n427) );
  XNOR2X1 U212 ( .A(n13), .B(n554), .Y(n428) );
  XNOR2X1 U213 ( .A(n13), .B(n555), .Y(n429) );
  XNOR2X1 U214 ( .A(n13), .B(n556), .Y(n430) );
  XNOR2X1 U215 ( .A(n13), .B(n557), .Y(n431) );
  XNOR2X1 U216 ( .A(n13), .B(n558), .Y(n432) );
  XNOR2X1 U217 ( .A(n13), .B(n559), .Y(n433) );
  XNOR2X1 U218 ( .A(n13), .B(n560), .Y(n434) );
  XNOR2X1 U219 ( .A(n13), .B(n561), .Y(n435) );
  XNOR2X1 U220 ( .A(n13), .B(n562), .Y(n436) );
  XNOR2X1 U221 ( .A(n13), .B(n563), .Y(n437) );
  XNOR2X1 U222 ( .A(n13), .B(n564), .Y(n438) );
  XNOR2X1 U223 ( .A(n13), .B(n565), .Y(n439) );
  XNOR2X1 U224 ( .A(n13), .B(n566), .Y(n440) );
  XNOR2X1 U225 ( .A(n13), .B(n567), .Y(n441) );
  XNOR2X1 U226 ( .A(n13), .B(n49), .Y(n442) );
  NAND2BX1 U227 ( .AN(n49), .B(n13), .Y(n443) );
  OAI22XL U228 ( .A0(n44), .A1(n595), .B0(n28), .B1(n461), .Y(n266) );
  AO21X1 U229 ( .A0(n44), .A1(n28), .B0(n444), .Y(n306) );
  OAI22XL U230 ( .A0(n44), .A1(n445), .B0(n28), .B1(n444), .Y(n96) );
  OAI22XL U231 ( .A0(n44), .A1(n446), .B0(n28), .B1(n445), .Y(n307) );
  OAI22XL U232 ( .A0(n44), .A1(n447), .B0(n28), .B1(n446), .Y(n308) );
  OAI22XL U233 ( .A0(n44), .A1(n448), .B0(n28), .B1(n447), .Y(n309) );
  OAI22XL U234 ( .A0(n44), .A1(n449), .B0(n28), .B1(n448), .Y(n122) );
  OAI22XL U235 ( .A0(n44), .A1(n450), .B0(n28), .B1(n449), .Y(n310) );
  OAI22XL U236 ( .A0(n44), .A1(n451), .B0(n28), .B1(n450), .Y(n311) );
  OAI22XL U237 ( .A0(n43), .A1(n452), .B0(n28), .B1(n451), .Y(n312) );
  OAI22XL U238 ( .A0(n43), .A1(n453), .B0(n27), .B1(n452), .Y(n313) );
  OAI22XL U239 ( .A0(n43), .A1(n454), .B0(n27), .B1(n453), .Y(n314) );
  OAI22XL U240 ( .A0(n43), .A1(n455), .B0(n27), .B1(n454), .Y(n315) );
  OAI22XL U241 ( .A0(n43), .A1(n456), .B0(n27), .B1(n455), .Y(n316) );
  OAI22XL U242 ( .A0(n43), .A1(n457), .B0(n27), .B1(n456), .Y(n317) );
  OAI22XL U243 ( .A0(n43), .A1(n458), .B0(n27), .B1(n457), .Y(n318) );
  OAI22XL U244 ( .A0(n43), .A1(n459), .B0(n27), .B1(n458), .Y(n319) );
  OAI22XL U245 ( .A0(n43), .A1(n460), .B0(n27), .B1(n459), .Y(n320) );
  NOR2BX1 U246 ( .AN(n49), .B(n27), .Y(n321) );
  XNOR2X1 U247 ( .A(n11), .B(n552), .Y(n444) );
  XNOR2X1 U248 ( .A(n11), .B(n553), .Y(n445) );
  XNOR2X1 U249 ( .A(n11), .B(n554), .Y(n446) );
  XNOR2X1 U250 ( .A(n11), .B(n555), .Y(n447) );
  XNOR2X1 U251 ( .A(n11), .B(n556), .Y(n448) );
  XNOR2X1 U252 ( .A(n11), .B(n557), .Y(n449) );
  XNOR2X1 U253 ( .A(n11), .B(n558), .Y(n450) );
  XNOR2X1 U254 ( .A(n11), .B(n559), .Y(n451) );
  XNOR2X1 U255 ( .A(n11), .B(n560), .Y(n452) );
  XNOR2X1 U256 ( .A(n11), .B(n561), .Y(n453) );
  XNOR2X1 U257 ( .A(n11), .B(n562), .Y(n454) );
  XNOR2X1 U258 ( .A(n11), .B(n563), .Y(n455) );
  XNOR2X1 U259 ( .A(n11), .B(n564), .Y(n456) );
  XNOR2X1 U260 ( .A(n11), .B(n565), .Y(n457) );
  XNOR2X1 U261 ( .A(n11), .B(n566), .Y(n458) );
  XNOR2X1 U262 ( .A(n11), .B(n567), .Y(n459) );
  XNOR2X1 U263 ( .A(n11), .B(n49), .Y(n460) );
  NAND2BX1 U264 ( .AN(n49), .B(n11), .Y(n461) );
  OAI22XL U265 ( .A0(n42), .A1(n596), .B0(n26), .B1(n479), .Y(n267) );
  AO21X1 U266 ( .A0(n42), .A1(n26), .B0(n462), .Y(n322) );
  OAI22XL U267 ( .A0(n42), .A1(n463), .B0(n26), .B1(n462), .Y(n108) );
  OAI22XL U268 ( .A0(n42), .A1(n464), .B0(n26), .B1(n463), .Y(n323) );
  OAI22XL U269 ( .A0(n42), .A1(n465), .B0(n26), .B1(n464), .Y(n324) );
  OAI22XL U270 ( .A0(n42), .A1(n466), .B0(n26), .B1(n465), .Y(n325) );
  OAI22XL U271 ( .A0(n42), .A1(n467), .B0(n26), .B1(n466), .Y(n326) );
  OAI22XL U272 ( .A0(n42), .A1(n468), .B0(n26), .B1(n467), .Y(n327) );
  OAI22XL U273 ( .A0(n42), .A1(n469), .B0(n26), .B1(n468), .Y(n328) );
  OAI22XL U274 ( .A0(n41), .A1(n470), .B0(n26), .B1(n469), .Y(n329) );
  OAI22XL U275 ( .A0(n41), .A1(n471), .B0(n25), .B1(n470), .Y(n330) );
  OAI22XL U276 ( .A0(n41), .A1(n472), .B0(n25), .B1(n471), .Y(n331) );
  OAI22XL U277 ( .A0(n41), .A1(n473), .B0(n25), .B1(n472), .Y(n332) );
  OAI22XL U278 ( .A0(n41), .A1(n474), .B0(n25), .B1(n473), .Y(n333) );
  OAI22XL U279 ( .A0(n41), .A1(n475), .B0(n25), .B1(n474), .Y(n334) );
  OAI22XL U280 ( .A0(n41), .A1(n476), .B0(n25), .B1(n475), .Y(n335) );
  OAI22XL U281 ( .A0(n41), .A1(n477), .B0(n25), .B1(n476), .Y(n336) );
  OAI22XL U282 ( .A0(n41), .A1(n478), .B0(n25), .B1(n477), .Y(n337) );
  NOR2BX1 U283 ( .AN(n49), .B(n25), .Y(n338) );
  XNOR2X1 U284 ( .A(n9), .B(n552), .Y(n462) );
  XNOR2X1 U285 ( .A(n9), .B(n553), .Y(n463) );
  XNOR2X1 U286 ( .A(n9), .B(n554), .Y(n464) );
  XNOR2X1 U287 ( .A(n9), .B(n555), .Y(n465) );
  XNOR2X1 U288 ( .A(n9), .B(n556), .Y(n466) );
  XNOR2X1 U289 ( .A(n9), .B(n557), .Y(n467) );
  XNOR2X1 U290 ( .A(n9), .B(n558), .Y(n468) );
  XNOR2X1 U291 ( .A(n9), .B(n559), .Y(n469) );
  XNOR2X1 U292 ( .A(n9), .B(n560), .Y(n470) );
  XNOR2X1 U293 ( .A(n9), .B(n561), .Y(n471) );
  XNOR2X1 U294 ( .A(n9), .B(n562), .Y(n472) );
  XNOR2X1 U295 ( .A(n9), .B(n563), .Y(n473) );
  XNOR2X1 U296 ( .A(n9), .B(n564), .Y(n474) );
  XNOR2X1 U297 ( .A(n9), .B(n565), .Y(n475) );
  XNOR2X1 U298 ( .A(n9), .B(n566), .Y(n476) );
  XNOR2X1 U299 ( .A(n9), .B(n567), .Y(n477) );
  XNOR2X1 U300 ( .A(n9), .B(n49), .Y(n478) );
  NAND2BX1 U301 ( .AN(n49), .B(n9), .Y(n479) );
  OAI22XL U302 ( .A0(n40), .A1(n597), .B0(n24), .B1(n497), .Y(n268) );
  AO21X1 U303 ( .A0(n40), .A1(n24), .B0(n480), .Y(n339) );
  OAI22XL U304 ( .A0(n40), .A1(n481), .B0(n24), .B1(n480), .Y(n340) );
  OAI22XL U305 ( .A0(n40), .A1(n482), .B0(n24), .B1(n481), .Y(n341) );
  OAI22XL U306 ( .A0(n40), .A1(n483), .B0(n24), .B1(n482), .Y(n342) );
  OAI22XL U307 ( .A0(n40), .A1(n484), .B0(n24), .B1(n483), .Y(n343) );
  OAI22XL U308 ( .A0(n40), .A1(n485), .B0(n24), .B1(n484), .Y(n344) );
  OAI22XL U309 ( .A0(n40), .A1(n486), .B0(n24), .B1(n485), .Y(n345) );
  OAI22XL U310 ( .A0(n40), .A1(n487), .B0(n24), .B1(n486), .Y(n346) );
  OAI22XL U311 ( .A0(n39), .A1(n488), .B0(n24), .B1(n487), .Y(n347) );
  OAI22XL U312 ( .A0(n39), .A1(n489), .B0(n23), .B1(n488), .Y(n348) );
  OAI22XL U313 ( .A0(n39), .A1(n490), .B0(n23), .B1(n489), .Y(n349) );
  OAI22XL U314 ( .A0(n39), .A1(n491), .B0(n23), .B1(n490), .Y(n350) );
  OAI22XL U315 ( .A0(n39), .A1(n492), .B0(n23), .B1(n491), .Y(n351) );
  OAI22XL U316 ( .A0(n39), .A1(n493), .B0(n23), .B1(n492), .Y(n352) );
  OAI22XL U317 ( .A0(n39), .A1(n494), .B0(n23), .B1(n493), .Y(n353) );
  OAI22XL U318 ( .A0(n39), .A1(n495), .B0(n23), .B1(n494), .Y(n354) );
  OAI22XL U319 ( .A0(n39), .A1(n496), .B0(n23), .B1(n495), .Y(n355) );
  NOR2BX1 U320 ( .AN(n49), .B(n23), .Y(n356) );
  XNOR2X1 U321 ( .A(n7), .B(n552), .Y(n480) );
  XNOR2X1 U322 ( .A(n7), .B(n553), .Y(n481) );
  XNOR2X1 U323 ( .A(n7), .B(n554), .Y(n482) );
  XNOR2X1 U324 ( .A(n7), .B(n555), .Y(n483) );
  XNOR2X1 U325 ( .A(n7), .B(n556), .Y(n484) );
  XNOR2X1 U326 ( .A(n7), .B(n557), .Y(n485) );
  XNOR2X1 U327 ( .A(n7), .B(n558), .Y(n486) );
  XNOR2X1 U328 ( .A(n7), .B(n559), .Y(n487) );
  XNOR2X1 U329 ( .A(n7), .B(n560), .Y(n488) );
  XNOR2X1 U330 ( .A(n7), .B(n561), .Y(n489) );
  XNOR2X1 U331 ( .A(n7), .B(n562), .Y(n490) );
  XNOR2X1 U332 ( .A(n7), .B(n563), .Y(n491) );
  XNOR2X1 U333 ( .A(n7), .B(n564), .Y(n492) );
  XNOR2X1 U334 ( .A(n7), .B(n565), .Y(n493) );
  XNOR2X1 U335 ( .A(n7), .B(n566), .Y(n494) );
  XNOR2X1 U336 ( .A(n7), .B(n567), .Y(n495) );
  XNOR2X1 U337 ( .A(n7), .B(n49), .Y(n496) );
  NAND2BX1 U338 ( .AN(n49), .B(n7), .Y(n497) );
  OAI22XL U339 ( .A0(n38), .A1(n598), .B0(n22), .B1(n515), .Y(n269) );
  AO21X1 U340 ( .A0(n38), .A1(n22), .B0(n498), .Y(n357) );
  OAI22XL U341 ( .A0(n38), .A1(n499), .B0(n22), .B1(n498), .Y(n140) );
  OAI22XL U342 ( .A0(n38), .A1(n500), .B0(n22), .B1(n499), .Y(n358) );
  OAI22XL U343 ( .A0(n38), .A1(n501), .B0(n22), .B1(n500), .Y(n359) );
  OAI22XL U344 ( .A0(n38), .A1(n502), .B0(n22), .B1(n501), .Y(n360) );
  OAI22XL U345 ( .A0(n38), .A1(n503), .B0(n22), .B1(n502), .Y(n361) );
  OAI22XL U346 ( .A0(n38), .A1(n504), .B0(n22), .B1(n503), .Y(n362) );
  OAI22XL U347 ( .A0(n38), .A1(n505), .B0(n22), .B1(n504), .Y(n363) );
  OAI22XL U348 ( .A0(n37), .A1(n506), .B0(n22), .B1(n505), .Y(n364) );
  OAI22XL U349 ( .A0(n37), .A1(n507), .B0(n21), .B1(n506), .Y(n365) );
  OAI22XL U350 ( .A0(n37), .A1(n508), .B0(n21), .B1(n507), .Y(n366) );
  OAI22XL U351 ( .A0(n37), .A1(n509), .B0(n21), .B1(n508), .Y(n367) );
  OAI22XL U352 ( .A0(n37), .A1(n510), .B0(n21), .B1(n509), .Y(n368) );
  OAI22XL U353 ( .A0(n37), .A1(n511), .B0(n21), .B1(n510), .Y(n369) );
  OAI22XL U354 ( .A0(n37), .A1(n512), .B0(n21), .B1(n511), .Y(n370) );
  OAI22XL U355 ( .A0(n37), .A1(n513), .B0(n21), .B1(n512), .Y(n371) );
  OAI22XL U356 ( .A0(n37), .A1(n514), .B0(n21), .B1(n513), .Y(n372) );
  NOR2BX1 U357 ( .AN(n49), .B(n21), .Y(n373) );
  XNOR2X1 U358 ( .A(n5), .B(n552), .Y(n498) );
  XNOR2X1 U359 ( .A(n5), .B(n553), .Y(n499) );
  XNOR2X1 U360 ( .A(n5), .B(n554), .Y(n500) );
  XNOR2X1 U361 ( .A(n5), .B(n555), .Y(n501) );
  XNOR2X1 U362 ( .A(n5), .B(n556), .Y(n502) );
  XNOR2X1 U363 ( .A(n5), .B(n557), .Y(n503) );
  XNOR2X1 U364 ( .A(n5), .B(n558), .Y(n504) );
  XNOR2X1 U365 ( .A(n5), .B(n559), .Y(n505) );
  XNOR2X1 U366 ( .A(n5), .B(n560), .Y(n506) );
  XNOR2X1 U367 ( .A(n5), .B(n561), .Y(n507) );
  XNOR2X1 U368 ( .A(n5), .B(n562), .Y(n508) );
  XNOR2X1 U369 ( .A(n5), .B(n563), .Y(n509) );
  XNOR2X1 U370 ( .A(n5), .B(n564), .Y(n510) );
  XNOR2X1 U371 ( .A(n5), .B(n565), .Y(n511) );
  XNOR2X1 U372 ( .A(n5), .B(n566), .Y(n512) );
  XNOR2X1 U373 ( .A(n5), .B(n567), .Y(n513) );
  XNOR2X1 U374 ( .A(n5), .B(n49), .Y(n514) );
  NAND2BX1 U375 ( .AN(n49), .B(n5), .Y(n515) );
  OAI22XL U376 ( .A0(n36), .A1(n599), .B0(n20), .B1(n533), .Y(n270) );
  AO21X1 U377 ( .A0(n36), .A1(n20), .B0(n516), .Y(n374) );
  OAI22XL U378 ( .A0(n36), .A1(n517), .B0(n20), .B1(n516), .Y(n160) );
  OAI22XL U379 ( .A0(n36), .A1(n518), .B0(n20), .B1(n517), .Y(n375) );
  OAI22XL U380 ( .A0(n36), .A1(n519), .B0(n20), .B1(n518), .Y(n376) );
  OAI22XL U381 ( .A0(n36), .A1(n520), .B0(n20), .B1(n519), .Y(n377) );
  OAI22XL U382 ( .A0(n36), .A1(n521), .B0(n20), .B1(n520), .Y(n378) );
  OAI22XL U383 ( .A0(n36), .A1(n522), .B0(n20), .B1(n521), .Y(n379) );
  OAI22XL U384 ( .A0(n36), .A1(n523), .B0(n20), .B1(n522), .Y(n380) );
  OAI22XL U385 ( .A0(n35), .A1(n524), .B0(n20), .B1(n523), .Y(n381) );
  OAI22XL U386 ( .A0(n35), .A1(n525), .B0(n19), .B1(n524), .Y(n382) );
  OAI22XL U387 ( .A0(n35), .A1(n526), .B0(n19), .B1(n525), .Y(n383) );
  OAI22XL U388 ( .A0(n35), .A1(n527), .B0(n19), .B1(n526), .Y(n384) );
  OAI22XL U389 ( .A0(n35), .A1(n528), .B0(n19), .B1(n527), .Y(n385) );
  OAI22XL U390 ( .A0(n35), .A1(n529), .B0(n19), .B1(n528), .Y(n386) );
  OAI22XL U391 ( .A0(n35), .A1(n530), .B0(n19), .B1(n529), .Y(n387) );
  OAI22XL U392 ( .A0(n35), .A1(n531), .B0(n19), .B1(n530), .Y(n388) );
  OAI22XL U393 ( .A0(n35), .A1(n532), .B0(n19), .B1(n531), .Y(n389) );
  NOR2BX1 U394 ( .AN(n49), .B(n19), .Y(n390) );
  XNOR2X1 U395 ( .A(n3), .B(n552), .Y(n516) );
  XNOR2X1 U396 ( .A(n3), .B(n553), .Y(n517) );
  XNOR2X1 U397 ( .A(n3), .B(n554), .Y(n518) );
  XNOR2X1 U398 ( .A(n3), .B(n555), .Y(n519) );
  XNOR2X1 U399 ( .A(n3), .B(n556), .Y(n520) );
  XNOR2X1 U400 ( .A(n3), .B(n557), .Y(n521) );
  XNOR2X1 U401 ( .A(n3), .B(n558), .Y(n522) );
  XNOR2X1 U402 ( .A(n3), .B(n559), .Y(n523) );
  XNOR2X1 U403 ( .A(n3), .B(n560), .Y(n524) );
  XNOR2X1 U404 ( .A(n3), .B(n561), .Y(n525) );
  XNOR2X1 U405 ( .A(n3), .B(n562), .Y(n526) );
  XNOR2X1 U406 ( .A(n3), .B(n563), .Y(n527) );
  XNOR2X1 U407 ( .A(n3), .B(n564), .Y(n528) );
  XNOR2X1 U408 ( .A(n3), .B(n565), .Y(n529) );
  XNOR2X1 U409 ( .A(n3), .B(n566), .Y(n530) );
  XNOR2X1 U410 ( .A(n3), .B(n567), .Y(n531) );
  XNOR2X1 U411 ( .A(n3), .B(n49), .Y(n532) );
  NAND2BX1 U412 ( .AN(n49), .B(n3), .Y(n533) );
  OAI22XL U413 ( .A0(n34), .A1(n600), .B0(n551), .B1(n18), .Y(n271) );
  AO21X1 U414 ( .A0(n34), .A1(n18), .B0(n534), .Y(n391) );
  OAI22XL U415 ( .A0(n34), .A1(n535), .B0(n534), .B1(n18), .Y(n392) );
  OAI22XL U416 ( .A0(n34), .A1(n536), .B0(n535), .B1(n18), .Y(n393) );
  OAI22XL U417 ( .A0(n34), .A1(n537), .B0(n536), .B1(n18), .Y(n394) );
  OAI22XL U418 ( .A0(n34), .A1(n538), .B0(n537), .B1(n18), .Y(n395) );
  OAI22XL U419 ( .A0(n34), .A1(n539), .B0(n538), .B1(n18), .Y(n396) );
  OAI22XL U420 ( .A0(n34), .A1(n540), .B0(n539), .B1(n18), .Y(n397) );
  OAI22XL U421 ( .A0(n34), .A1(n541), .B0(n540), .B1(n18), .Y(n398) );
  OAI22XL U422 ( .A0(n33), .A1(n542), .B0(n541), .B1(n18), .Y(n399) );
  OAI22XL U423 ( .A0(n33), .A1(n543), .B0(n542), .B1(n17), .Y(n400) );
  OAI22XL U424 ( .A0(n33), .A1(n544), .B0(n543), .B1(n17), .Y(n401) );
  OAI22XL U425 ( .A0(n33), .A1(n545), .B0(n544), .B1(n17), .Y(n402) );
  OAI22XL U426 ( .A0(n33), .A1(n546), .B0(n545), .B1(n17), .Y(n403) );
  OAI22XL U427 ( .A0(n33), .A1(n547), .B0(n546), .B1(n17), .Y(n404) );
  OAI22XL U428 ( .A0(n33), .A1(n548), .B0(n547), .B1(n17), .Y(n405) );
  OAI22XL U429 ( .A0(n33), .A1(n549), .B0(n548), .B1(n17), .Y(n406) );
  OAI22XL U430 ( .A0(n33), .A1(n550), .B0(n549), .B1(n17), .Y(n407) );
  NOR2BX1 U431 ( .AN(n49), .B(n17), .Y(product_0_) );
  XNOR2X1 U432 ( .A(n1), .B(n552), .Y(n534) );
  XNOR2X1 U433 ( .A(n1), .B(n553), .Y(n535) );
  XNOR2X1 U434 ( .A(n1), .B(n554), .Y(n536) );
  XNOR2X1 U435 ( .A(n1), .B(n555), .Y(n537) );
  XNOR2X1 U436 ( .A(n1), .B(n556), .Y(n538) );
  XNOR2X1 U437 ( .A(n1), .B(n557), .Y(n539) );
  XNOR2X1 U438 ( .A(n1), .B(n558), .Y(n540) );
  XNOR2X1 U439 ( .A(n1), .B(n559), .Y(n541) );
  XNOR2X1 U440 ( .A(n1), .B(n560), .Y(n542) );
  XNOR2X1 U441 ( .A(n1), .B(n561), .Y(n543) );
  XNOR2X1 U442 ( .A(n1), .B(n562), .Y(n544) );
  XNOR2X1 U443 ( .A(n1), .B(n563), .Y(n545) );
  XNOR2X1 U444 ( .A(n1), .B(n564), .Y(n546) );
  XNOR2X1 U445 ( .A(n1), .B(n565), .Y(n547) );
  XNOR2X1 U446 ( .A(n1), .B(n566), .Y(n548) );
  XNOR2X1 U447 ( .A(n1), .B(n567), .Y(n549) );
  XNOR2X1 U448 ( .A(n1), .B(n49), .Y(n550) );
  NAND2BX1 U449 ( .AN(n49), .B(n1), .Y(n551) );
  CLKINVX1 U466 ( .A(n15), .Y(n593) );
  CLKINVX1 U467 ( .A(n13), .Y(n594) );
  CLKINVX1 U468 ( .A(n11), .Y(n595) );
  CLKINVX1 U469 ( .A(n9), .Y(n596) );
  CLKINVX1 U470 ( .A(n7), .Y(n597) );
  CLKINVX1 U471 ( .A(n5), .Y(n598) );
  CLKINVX1 U472 ( .A(n3), .Y(n599) );
  CLKINVX1 U473 ( .A(n1), .Y(n600) );
  NAND2X1 U474 ( .A(n569), .B(n585), .Y(n577) );
  XOR2X1 U475 ( .A(a[14]), .B(a[15]), .Y(n569) );
  XNOR2X1 U476 ( .A(a[14]), .B(a[13]), .Y(n585) );
  NAND2X1 U477 ( .A(n570), .B(n586), .Y(n578) );
  XOR2X1 U478 ( .A(a[12]), .B(a[13]), .Y(n570) );
  XNOR2X1 U479 ( .A(a[12]), .B(a[11]), .Y(n586) );
  NAND2X1 U480 ( .A(n571), .B(n587), .Y(n579) );
  XOR2X1 U481 ( .A(a[10]), .B(a[11]), .Y(n571) );
  XNOR2X1 U482 ( .A(a[10]), .B(a[9]), .Y(n587) );
  NAND2X1 U483 ( .A(n572), .B(n588), .Y(n580) );
  XOR2X1 U484 ( .A(a[8]), .B(a[9]), .Y(n572) );
  XNOR2X1 U485 ( .A(a[8]), .B(a[7]), .Y(n588) );
  NAND2X1 U486 ( .A(n573), .B(n589), .Y(n581) );
  XOR2X1 U487 ( .A(a[6]), .B(a[7]), .Y(n573) );
  XNOR2X1 U488 ( .A(a[6]), .B(a[5]), .Y(n589) );
  NAND2X1 U489 ( .A(n574), .B(n590), .Y(n582) );
  XOR2X1 U490 ( .A(a[4]), .B(a[5]), .Y(n574) );
  XNOR2X1 U491 ( .A(a[4]), .B(a[3]), .Y(n590) );
  NAND2X1 U492 ( .A(n575), .B(n591), .Y(n583) );
  XOR2X1 U493 ( .A(a[2]), .B(a[3]), .Y(n575) );
  XNOR2X1 U494 ( .A(a[2]), .B(a[1]), .Y(n591) );
  NAND2X1 U495 ( .A(n576), .B(n592), .Y(n584) );
  XOR2X1 U496 ( .A(a[0]), .B(a[1]), .Y(n576) );
  CLKINVX1 U497 ( .A(a[0]), .Y(n592) );
  CLKBUFX3 U500 ( .A(b_2_), .Y(n566) );
  CLKBUFX3 U501 ( .A(b_4_), .Y(n564) );
  CLKBUFX3 U502 ( .A(b_5_), .Y(n563) );
  CLKBUFX3 U503 ( .A(b_6_), .Y(n562) );
  CLKBUFX3 U504 ( .A(b_0_), .Y(n49) );
  CLKBUFX3 U505 ( .A(b_3_), .Y(n565) );
  CLKBUFX3 U506 ( .A(b_9_), .Y(n559) );
  CLKBUFX3 U507 ( .A(b_12_), .Y(n556) );
  CLKBUFX3 U508 ( .A(b_7_), .Y(n561) );
  CLKBUFX3 U509 ( .A(b_14_), .Y(n554) );
  CLKBUFX3 U510 ( .A(n591), .Y(n20) );
  CLKBUFX3 U511 ( .A(n590), .Y(n22) );
  CLKBUFX3 U512 ( .A(n588), .Y(n26) );
  CLKBUFX3 U513 ( .A(n589), .Y(n24) );
  CLKBUFX3 U514 ( .A(n585), .Y(n32) );
  CLKBUFX3 U515 ( .A(n586), .Y(n30) );
  CLKBUFX3 U516 ( .A(n587), .Y(n28) );
  CLKBUFX3 U517 ( .A(b_10_), .Y(n558) );
  CLKBUFX3 U518 ( .A(b_15_), .Y(n553) );
  CLKBUFX3 U519 ( .A(n591), .Y(n19) );
  CLKBUFX3 U520 ( .A(n590), .Y(n21) );
  CLKBUFX3 U521 ( .A(n589), .Y(n23) );
  CLKBUFX3 U522 ( .A(n588), .Y(n25) );
  CLKBUFX3 U523 ( .A(n587), .Y(n27) );
  CLKBUFX3 U524 ( .A(n586), .Y(n29) );
  CLKBUFX3 U525 ( .A(n585), .Y(n31) );
  CLKBUFX3 U526 ( .A(b_8_), .Y(n560) );
  CLKBUFX3 U527 ( .A(b_11_), .Y(n557) );
  CLKBUFX3 U528 ( .A(b_16_), .Y(n552) );
  CLKBUFX3 U529 ( .A(n583), .Y(n35) );
  CLKBUFX3 U530 ( .A(n582), .Y(n37) );
  CLKBUFX3 U531 ( .A(n581), .Y(n39) );
  CLKBUFX3 U532 ( .A(n580), .Y(n41) );
  CLKBUFX3 U533 ( .A(n579), .Y(n43) );
  CLKBUFX3 U534 ( .A(n578), .Y(n45) );
  CLKBUFX3 U535 ( .A(n577), .Y(n47) );
  CLKBUFX3 U536 ( .A(n584), .Y(n33) );
  CLKBUFX3 U537 ( .A(n583), .Y(n36) );
  CLKBUFX3 U538 ( .A(n582), .Y(n38) );
  CLKBUFX3 U539 ( .A(n580), .Y(n42) );
  CLKBUFX3 U540 ( .A(n581), .Y(n40) );
  CLKBUFX3 U541 ( .A(n577), .Y(n48) );
  CLKBUFX3 U542 ( .A(n578), .Y(n46) );
  CLKBUFX3 U543 ( .A(n579), .Y(n44) );
  CLKBUFX3 U544 ( .A(n584), .Y(n34) );
  CLKBUFX3 U545 ( .A(n592), .Y(n18) );
  CLKBUFX3 U546 ( .A(n592), .Y(n17) );
  CLKBUFX3 U547 ( .A(b_1_), .Y(n567) );
  CLKBUFX3 U548 ( .A(b_13_), .Y(n555) );
  CLKBUFX3 U549 ( .A(a[1]), .Y(n1) );
  CLKBUFX3 U550 ( .A(a[3]), .Y(n3) );
  CLKBUFX3 U551 ( .A(a[5]), .Y(n5) );
  CLKBUFX3 U552 ( .A(a[7]), .Y(n7) );
  CLKBUFX3 U553 ( .A(a[9]), .Y(n9) );
  CLKBUFX3 U554 ( .A(a[11]), .Y(n11) );
  CLKBUFX3 U555 ( .A(a[13]), .Y(n13) );
  CLKBUFX3 U556 ( .A(a[15]), .Y(n15) );
endmodule


module FAS_DW_mult_uns_6 ( a, b, product_31_, product_30_, product_29_, 
        product_28_, product_27_, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_, product_14_, 
        product_13_, product_12_, product_11_, product_10_, product_9_, 
        product_8_, product_7_, product_6_, product_5_, product_4_, product_3_, 
        product_2_, product_1_, product_0_ );
  input [31:0] a;
  input b;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;

  NOR2X1 U3 ( .A(n2), .B(n3), .Y(product_31_) );
  NOR2X1 U4 ( .A(n2), .B(n4), .Y(product_30_) );
  NOR2X1 U5 ( .A(n2), .B(n5), .Y(product_29_) );
  NOR2X1 U6 ( .A(n2), .B(n6), .Y(product_28_) );
  NOR2X1 U7 ( .A(n2), .B(n7), .Y(product_27_) );
  NOR2X1 U8 ( .A(n2), .B(n8), .Y(product_26_) );
  NOR2X1 U9 ( .A(n2), .B(n9), .Y(product_25_) );
  NOR2X1 U10 ( .A(n2), .B(n10), .Y(product_24_) );
  NOR2X1 U11 ( .A(n2), .B(n11), .Y(product_23_) );
  NOR2X1 U12 ( .A(n2), .B(n12), .Y(product_22_) );
  NOR2X1 U13 ( .A(n2), .B(n13), .Y(product_21_) );
  NOR2X1 U14 ( .A(n2), .B(n14), .Y(product_20_) );
  NOR2X1 U15 ( .A(n2), .B(n15), .Y(product_19_) );
  NOR2X1 U16 ( .A(n2), .B(n16), .Y(product_18_) );
  NOR2X1 U17 ( .A(n2), .B(n17), .Y(product_17_) );
  NOR2X1 U18 ( .A(n2), .B(n18), .Y(product_16_) );
  NOR2X1 U19 ( .A(n1), .B(n19), .Y(product_15_) );
  NOR2X1 U20 ( .A(n1), .B(n20), .Y(product_14_) );
  NOR2X1 U21 ( .A(n1), .B(n21), .Y(product_13_) );
  NOR2X1 U22 ( .A(n1), .B(n22), .Y(product_12_) );
  NOR2X1 U23 ( .A(n1), .B(n23), .Y(product_11_) );
  NOR2X1 U24 ( .A(n1), .B(n24), .Y(product_10_) );
  NOR2X1 U25 ( .A(n1), .B(n25), .Y(product_9_) );
  NOR2X1 U26 ( .A(n1), .B(n26), .Y(product_8_) );
  NOR2X1 U27 ( .A(n1), .B(n27), .Y(product_7_) );
  NOR2X1 U28 ( .A(n1), .B(n28), .Y(product_6_) );
  NOR2X1 U29 ( .A(n1), .B(n29), .Y(product_5_) );
  NOR2X1 U30 ( .A(n1), .B(n30), .Y(product_4_) );
  NOR2X1 U31 ( .A(n1), .B(n31), .Y(product_3_) );
  NOR2X1 U32 ( .A(n1), .B(n32), .Y(product_2_) );
  NOR2X1 U33 ( .A(n1), .B(n33), .Y(product_1_) );
  NOR2X1 U34 ( .A(n1), .B(n34), .Y(product_0_) );
  CLKINVX1 U70 ( .A(a[1]), .Y(n33) );
  CLKINVX1 U71 ( .A(a[0]), .Y(n34) );
  CLKBUFX3 U72 ( .A(n35), .Y(n1) );
  CLKBUFX3 U73 ( .A(n35), .Y(n2) );
  CLKINVX1 U74 ( .A(b), .Y(n35) );
  CLKINVX1 U75 ( .A(a[2]), .Y(n32) );
  CLKINVX1 U76 ( .A(a[3]), .Y(n31) );
  CLKINVX1 U77 ( .A(a[4]), .Y(n30) );
  CLKINVX1 U78 ( .A(a[5]), .Y(n29) );
  CLKINVX1 U79 ( .A(a[6]), .Y(n28) );
  CLKINVX1 U80 ( .A(a[7]), .Y(n27) );
  CLKINVX1 U81 ( .A(a[8]), .Y(n26) );
  CLKINVX1 U82 ( .A(a[9]), .Y(n25) );
  CLKINVX1 U83 ( .A(a[10]), .Y(n24) );
  CLKINVX1 U84 ( .A(a[11]), .Y(n23) );
  CLKINVX1 U85 ( .A(a[12]), .Y(n22) );
  CLKINVX1 U86 ( .A(a[13]), .Y(n21) );
  CLKINVX1 U87 ( .A(a[14]), .Y(n20) );
  CLKINVX1 U88 ( .A(a[16]), .Y(n18) );
  CLKINVX1 U89 ( .A(a[15]), .Y(n19) );
  CLKINVX1 U90 ( .A(a[17]), .Y(n17) );
  CLKINVX1 U91 ( .A(a[18]), .Y(n16) );
  CLKINVX1 U92 ( .A(a[19]), .Y(n15) );
  CLKINVX1 U93 ( .A(a[20]), .Y(n14) );
  CLKINVX1 U94 ( .A(a[21]), .Y(n13) );
  CLKINVX1 U95 ( .A(a[22]), .Y(n12) );
  CLKINVX1 U96 ( .A(a[23]), .Y(n11) );
  CLKINVX1 U97 ( .A(a[24]), .Y(n10) );
  CLKINVX1 U98 ( .A(a[25]), .Y(n9) );
  CLKINVX1 U99 ( .A(a[26]), .Y(n8) );
  CLKINVX1 U100 ( .A(a[27]), .Y(n7) );
  CLKINVX1 U101 ( .A(a[28]), .Y(n6) );
  CLKINVX1 U102 ( .A(a[29]), .Y(n5) );
  CLKINVX1 U103 ( .A(a[30]), .Y(n4) );
  CLKINVX1 U104 ( .A(a[31]), .Y(n3) );
endmodule


module FAS_DW_mult_tc_29 ( a, product_23_, product_22_, product_21_, 
        product_20_, product_19_, product_18_, product_17_, product_16_, 
        product_15_, product_14_, product_13_, product_12_, product_11_, 
        product_10_, product_9_, product_8_, product_7_, product_6_, 
        product_5_, product_4_, product_3_, product_2_, product_1_ );
  input [15:0] a;
  output product_23_, product_22_, product_21_, product_20_, product_19_,
         product_18_, product_17_, product_16_, product_15_, product_14_,
         product_13_, product_12_, product_11_, product_10_, product_9_,
         product_8_, product_7_, product_6_, product_5_, product_4_,
         product_3_, product_2_, product_1_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  CLKINVX1 U1 ( .A(n1), .Y(product_23_) );
  ADDFXL U2 ( .A(a[15]), .B(n43), .CI(n2), .CO(n1), .S(product_22_) );
  ADDFXL U3 ( .A(n44), .B(a[14]), .CI(n3), .CO(n2), .S(product_21_) );
  ADDFXL U4 ( .A(n45), .B(a[13]), .CI(n4), .CO(n3), .S(product_20_) );
  ADDFXL U5 ( .A(n46), .B(a[12]), .CI(n5), .CO(n4), .S(product_19_) );
  ADDFXL U6 ( .A(n42), .B(a[11]), .CI(n6), .CO(n5), .S(product_18_) );
  ADDFXL U7 ( .A(n22), .B(n47), .CI(n7), .CO(n6), .S(product_17_) );
  ADDFXL U8 ( .A(n24), .B(n23), .CI(n8), .CO(n7), .S(product_16_) );
  ADDFXL U9 ( .A(n25), .B(n26), .CI(n9), .CO(n8), .S(product_15_) );
  ADDFXL U10 ( .A(n27), .B(n28), .CI(n10), .CO(n9), .S(product_14_) );
  ADDFXL U11 ( .A(n29), .B(n30), .CI(n11), .CO(n10), .S(product_13_) );
  ADDFXL U12 ( .A(n31), .B(n32), .CI(n12), .CO(n11), .S(product_12_) );
  ADDFXL U13 ( .A(n33), .B(n34), .CI(n13), .CO(n12), .S(product_11_) );
  ADDFXL U14 ( .A(n35), .B(n36), .CI(n14), .CO(n13), .S(product_10_) );
  ADDFXL U15 ( .A(n37), .B(n38), .CI(n15), .CO(n14), .S(product_9_) );
  ADDFXL U16 ( .A(n39), .B(n40), .CI(n16), .CO(n15), .S(product_8_) );
  ADDFXL U17 ( .A(n41), .B(a[5]), .CI(n17), .CO(n16), .S(product_7_) );
  ADDFXL U18 ( .A(a[5]), .B(a[4]), .CI(n18), .CO(n17), .S(product_6_) );
  ADDFXL U19 ( .A(a[4]), .B(a[3]), .CI(n19), .CO(n18), .S(product_5_) );
  ADDFXL U20 ( .A(a[3]), .B(a[2]), .CI(n20), .CO(n19), .S(product_4_) );
  ADDFXL U21 ( .A(a[2]), .B(a[1]), .CI(n21), .CO(n20), .S(product_3_) );
  ADDHXL U22 ( .A(a[0]), .B(a[1]), .CO(n21), .S(product_2_) );
  ADDFXL U23 ( .A(n48), .B(a[15]), .CI(a[14]), .CO(n22), .S(n23) );
  ADDFXL U24 ( .A(a[13]), .B(n49), .CI(a[14]), .CO(n24), .S(n25) );
  ADDFXL U25 ( .A(a[12]), .B(n50), .CI(a[13]), .CO(n26), .S(n27) );
  ADDFXL U26 ( .A(a[11]), .B(n51), .CI(a[12]), .CO(n28), .S(n29) );
  ADDFXL U27 ( .A(a[10]), .B(n52), .CI(a[11]), .CO(n30), .S(n31) );
  ADDFXL U28 ( .A(a[9]), .B(n53), .CI(a[10]), .CO(n32), .S(n33) );
  ADDFXL U29 ( .A(a[8]), .B(n54), .CI(a[9]), .CO(n34), .S(n35) );
  ADDFXL U30 ( .A(a[7]), .B(n55), .CI(a[8]), .CO(n36), .S(n37) );
  ADDFXL U31 ( .A(a[6]), .B(n56), .CI(a[7]), .CO(n38), .S(n39) );
  XNOR2X1 U32 ( .A(a[6]), .B(n57), .Y(n41) );
  OR2X1 U33 ( .A(a[6]), .B(n57), .Y(n40) );
  CLKINVX1 U54 ( .A(a[10]), .Y(n47) );
  CLKINVX1 U55 ( .A(a[15]), .Y(n42) );
  CLKINVX1 U56 ( .A(a[11]), .Y(n46) );
  CLKINVX1 U57 ( .A(a[12]), .Y(n45) );
  CLKINVX1 U58 ( .A(a[13]), .Y(n44) );
  CLKINVX1 U59 ( .A(a[14]), .Y(n43) );
  CLKINVX1 U60 ( .A(a[1]), .Y(n56) );
  CLKINVX1 U61 ( .A(a[2]), .Y(n55) );
  CLKINVX1 U62 ( .A(a[3]), .Y(n54) );
  CLKINVX1 U63 ( .A(a[4]), .Y(n53) );
  CLKINVX1 U64 ( .A(a[5]), .Y(n52) );
  CLKINVX1 U65 ( .A(a[6]), .Y(n51) );
  CLKINVX1 U66 ( .A(a[7]), .Y(n50) );
  CLKINVX1 U67 ( .A(a[9]), .Y(n48) );
  CLKINVX1 U68 ( .A(a[8]), .Y(n49) );
  CLKINVX1 U69 ( .A(a[0]), .Y(n57) );
  BUFX2 U70 ( .A(a[0]), .Y(product_1_) );
endmodule


module FAS_DW_mult_tc_30 ( a, product );
  input [15:0] a;
  output [27:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84, n85, n86;

  CLKINVX1 U3 ( .A(n2), .Y(product[26]) );
  ADDFXL U4 ( .A(a[15]), .B(n68), .CI(n3), .CO(n2), .S(product[25]) );
  ADDFXL U5 ( .A(n69), .B(a[14]), .CI(n4), .CO(n3), .S(product[24]) );
  ADDFXL U6 ( .A(n70), .B(a[13]), .CI(n5), .CO(n4), .S(product[23]) );
  ADDFXL U7 ( .A(n26), .B(a[12]), .CI(n6), .CO(n5), .S(product[22]) );
  ADDFXL U8 ( .A(n27), .B(n28), .CI(n7), .CO(n6), .S(product[21]) );
  ADDFXL U9 ( .A(n29), .B(n30), .CI(n8), .CO(n7), .S(product[20]) );
  ADDFXL U10 ( .A(n32), .B(n31), .CI(n9), .CO(n8), .S(product[19]) );
  ADDFXL U11 ( .A(n35), .B(n33), .CI(n10), .CO(n9), .S(product[18]) );
  ADDFXL U12 ( .A(n36), .B(n38), .CI(n11), .CO(n10), .S(product[17]) );
  ADDFXL U13 ( .A(n39), .B(n41), .CI(n12), .CO(n11), .S(product[16]) );
  ADDFXL U14 ( .A(n42), .B(n44), .CI(n13), .CO(n12), .S(product[15]) );
  ADDFXL U15 ( .A(n45), .B(n47), .CI(n14), .CO(n13), .S(product[14]) );
  ADDFXL U16 ( .A(n48), .B(n50), .CI(n15), .CO(n14), .S(product[13]) );
  ADDFXL U17 ( .A(n51), .B(n53), .CI(n16), .CO(n15), .S(product[12]) );
  ADDFXL U18 ( .A(n54), .B(n55), .CI(n17), .CO(n16), .S(product[11]) );
  ADDFXL U19 ( .A(n56), .B(n59), .CI(n18), .CO(n17), .S(product[10]) );
  ADDFXL U20 ( .A(n60), .B(n61), .CI(n19), .CO(n18), .S(product[9]) );
  ADDFXL U21 ( .A(n62), .B(n63), .CI(n20), .CO(n19), .S(product[8]) );
  ADDFXL U22 ( .A(n64), .B(n65), .CI(n21), .CO(n20), .S(product[7]) );
  ADDFXL U23 ( .A(n66), .B(a[4]), .CI(n22), .CO(n21), .S(product[6]) );
  ADDFXL U24 ( .A(a[5]), .B(a[3]), .CI(n23), .CO(n22), .S(product[5]) );
  ADDFXL U25 ( .A(a[4]), .B(a[2]), .CI(n24), .CO(n23), .S(product[4]) );
  ADDFXL U26 ( .A(a[3]), .B(a[1]), .CI(n25), .CO(n24), .S(product[3]) );
  ADDHXL U27 ( .A(a[0]), .B(a[2]), .CO(n25), .S(product[2]) );
  ADDFXL U28 ( .A(n71), .B(n68), .CI(a[15]), .CO(n26), .S(n27) );
  ADDFXL U29 ( .A(n69), .B(a[14]), .CI(n72), .CO(n28), .S(n29) );
  ADDFXL U30 ( .A(n70), .B(a[13]), .CI(n73), .CO(n30), .S(n31) );
  ADDFXL U31 ( .A(n74), .B(a[12]), .CI(n34), .CO(n32), .S(n33) );
  CMPR42X1 U32 ( .A(n75), .B(n72), .C(n71), .D(n67), .ICI(n37), .S(n36), .ICO(
        n34), .CO(n35) );
  CMPR42X1 U33 ( .A(a[10]), .B(n76), .C(n67), .D(n84), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U34 ( .A(a[15]), .B(n73), .C(n77), .D(n85), .ICI(n43), .S(n42), 
        .ICO(n40), .CO(n41) );
  CMPR42X1 U35 ( .A(n78), .B(n74), .C(n86), .D(n84), .ICI(n46), .S(n45), .ICO(
        n43), .CO(n44) );
  CMPR42X1 U36 ( .A(n79), .B(n75), .C(a[11]), .D(n85), .ICI(n49), .S(n48), 
        .ICO(n46), .CO(n47) );
  CMPR42X1 U37 ( .A(n80), .B(n76), .C(a[10]), .D(n86), .ICI(n52), .S(n51), 
        .ICO(n49), .CO(n50) );
  CMPR42X1 U38 ( .A(n81), .B(n77), .C(a[9]), .D(a[11]), .ICI(n57), .S(n54), 
        .ICO(n52), .CO(n53) );
  ADDFXL U39 ( .A(a[8]), .B(a[10]), .CI(n58), .CO(n55), .S(n56) );
  XNOR2X1 U40 ( .A(n78), .B(n82), .Y(n58) );
  OR2X1 U41 ( .A(n78), .B(n82), .Y(n57) );
  ADDFXL U42 ( .A(a[7]), .B(n79), .CI(a[9]), .CO(n59), .S(n60) );
  ADDFXL U43 ( .A(a[6]), .B(n80), .CI(a[8]), .CO(n61), .S(n62) );
  ADDFXL U44 ( .A(a[5]), .B(n81), .CI(a[7]), .CO(n63), .S(n64) );
  XNOR2X1 U45 ( .A(a[6]), .B(n82), .Y(n66) );
  OR2X1 U46 ( .A(a[6]), .B(n82), .Y(n65) );
  CLKBUFX3 U70 ( .A(product[26]), .Y(product[27]) );
  CLKBUFX3 U71 ( .A(a[12]), .Y(n86) );
  CLKBUFX3 U72 ( .A(a[13]), .Y(n85) );
  CLKBUFX3 U73 ( .A(a[14]), .Y(n84) );
  CLKINVX1 U74 ( .A(a[6]), .Y(n76) );
  CLKINVX1 U75 ( .A(a[7]), .Y(n75) );
  CLKINVX1 U76 ( .A(a[5]), .Y(n77) );
  CLKINVX1 U77 ( .A(a[4]), .Y(n78) );
  CLKINVX1 U78 ( .A(a[9]), .Y(n73) );
  CLKINVX1 U79 ( .A(a[10]), .Y(n72) );
  CLKINVX1 U80 ( .A(a[15]), .Y(n67) );
  CLKINVX1 U81 ( .A(a[8]), .Y(n74) );
  CLKINVX1 U82 ( .A(a[0]), .Y(n82) );
  CLKINVX1 U83 ( .A(a[1]), .Y(n81) );
  CLKINVX1 U84 ( .A(a[2]), .Y(n80) );
  CLKINVX1 U85 ( .A(a[3]), .Y(n79) );
  CLKINVX1 U86 ( .A(a[11]), .Y(n71) );
  CLKINVX1 U87 ( .A(a[14]), .Y(n68) );
  CLKINVX1 U88 ( .A(a[12]), .Y(n70) );
  CLKINVX1 U89 ( .A(a[13]), .Y(n69) );
  BUFX2 U90 ( .A(a[0]), .Y(product[0]) );
  BUFX2 U91 ( .A(a[1]), .Y(product[1]) );
endmodule


module FAS_DW_mult_tc_31 ( a, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_, product_14_, 
        product_13_, product_12_, product_11_, product_10_, product_9_, 
        product_8_, product_7_, product_6_, product_5_, product_4_, product_3_, 
        product_2_, product_1_ );
  input [15:0] a;
  output product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;

  CLKINVX1 U1 ( .A(n43), .Y(product_26_) );
  ADDFXL U3 ( .A(a[14]), .B(a[15]), .CI(n3), .CO(product_24_), .S(product_23_)
         );
  ADDFXL U4 ( .A(a[13]), .B(a[15]), .CI(n4), .CO(n3), .S(product_22_) );
  ADDFXL U5 ( .A(a[12]), .B(a[15]), .CI(n5), .CO(n4), .S(product_21_) );
  ADDFXL U6 ( .A(n21), .B(a[11]), .CI(n6), .CO(n5), .S(product_20_) );
  ADDFXL U7 ( .A(n23), .B(n22), .CI(n7), .CO(n6), .S(product_19_) );
  ADDFXL U8 ( .A(n25), .B(n24), .CI(n8), .CO(n7), .S(product_18_) );
  ADDFXL U9 ( .A(n27), .B(n26), .CI(n9), .CO(n8), .S(product_17_) );
  ADDFXL U10 ( .A(n29), .B(n28), .CI(n10), .CO(n9), .S(product_16_) );
  ADDFXL U11 ( .A(n30), .B(n31), .CI(n11), .CO(n10), .S(product_15_) );
  ADDFXL U12 ( .A(n32), .B(n33), .CI(n12), .CO(n11), .S(product_14_) );
  ADDFXL U13 ( .A(n34), .B(n35), .CI(n13), .CO(n12), .S(product_13_) );
  ADDFXL U14 ( .A(n36), .B(n37), .CI(n14), .CO(n13), .S(product_12_) );
  ADDFXL U15 ( .A(n38), .B(n39), .CI(n15), .CO(n14), .S(product_11_) );
  ADDFXL U16 ( .A(n40), .B(n41), .CI(n16), .CO(n15), .S(product_10_) );
  ADDFXL U17 ( .A(n42), .B(a[0]), .CI(n17), .CO(n16), .S(product_9_) );
  ADDFXL U18 ( .A(a[7]), .B(a[3]), .CI(n18), .CO(n17), .S(product_8_) );
  ADDFXL U19 ( .A(a[6]), .B(a[2]), .CI(n19), .CO(n18), .S(product_7_) );
  ADDFXL U20 ( .A(a[5]), .B(a[1]), .CI(n20), .CO(n19), .S(product_6_) );
  ADDHXL U21 ( .A(a[0]), .B(a[4]), .CO(n20), .S(product_5_) );
  ADDFXL U22 ( .A(a[10]), .B(a[15]), .CI(a[14]), .CO(n21), .S(n22) );
  ADDFXL U23 ( .A(a[9]), .B(a[15]), .CI(a[13]), .CO(n23), .S(n24) );
  ADDFXL U24 ( .A(a[8]), .B(a[15]), .CI(a[12]), .CO(n25), .S(n26) );
  ADDFXL U25 ( .A(a[7]), .B(a[15]), .CI(a[11]), .CO(n27), .S(n28) );
  ADDFXL U26 ( .A(a[6]), .B(a[14]), .CI(a[10]), .CO(n29), .S(n30) );
  ADDFXL U27 ( .A(a[5]), .B(a[13]), .CI(a[9]), .CO(n31), .S(n32) );
  ADDFXL U28 ( .A(a[4]), .B(a[12]), .CI(a[8]), .CO(n33), .S(n34) );
  ADDFXL U29 ( .A(a[3]), .B(a[11]), .CI(a[7]), .CO(n35), .S(n36) );
  ADDFXL U30 ( .A(a[2]), .B(a[10]), .CI(a[6]), .CO(n37), .S(n38) );
  ADDFXL U31 ( .A(a[1]), .B(a[9]), .CI(a[5]), .CO(n39), .S(n40) );
  ADDHXL U32 ( .A(a[8]), .B(a[4]), .CO(n41), .S(n42) );
  CLKINVX1 U38 ( .A(a[15]), .Y(n43) );
  BUFX2 U39 ( .A(a[0]), .Y(product_1_) );
  BUFX2 U40 ( .A(a[1]), .Y(product_2_) );
  BUFX2 U41 ( .A(a[2]), .Y(product_3_) );
  BUFX2 U42 ( .A(a[3]), .Y(product_4_) );
  BUFX2 U43 ( .A(product_26_), .Y(product_25_) );
endmodule


module FAS_DW_mult_tc_32 ( a, product_23_, product_22_, product_21_, 
        product_20_, product_19_, product_18_, product_17_, product_16_, 
        product_15_, product_14_, product_13_, product_12_, product_11_, 
        product_10_, product_9_, product_8_, product_7_, product_6_, 
        product_5_, product_4_, product_3_, product_2_, product_1_ );
  input [15:0] a;
  output product_23_, product_22_, product_21_, product_20_, product_19_,
         product_18_, product_17_, product_16_, product_15_, product_14_,
         product_13_, product_12_, product_11_, product_10_, product_9_,
         product_8_, product_7_, product_6_, product_5_, product_4_,
         product_3_, product_2_, product_1_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65;

  CLKINVX1 U1 ( .A(n1), .Y(product_23_) );
  ADDFXL U2 ( .A(a[15]), .B(n52), .CI(n2), .CO(n1), .S(product_22_) );
  ADDFXL U3 ( .A(n23), .B(a[14]), .CI(n3), .CO(n2), .S(product_21_) );
  ADDFXL U4 ( .A(n24), .B(n25), .CI(n4), .CO(n3), .S(product_20_) );
  ADDFXL U5 ( .A(n26), .B(n27), .CI(n5), .CO(n4), .S(product_19_) );
  ADDFXL U6 ( .A(n28), .B(n29), .CI(n6), .CO(n5), .S(product_18_) );
  ADDFXL U7 ( .A(n30), .B(n31), .CI(n7), .CO(n6), .S(product_17_) );
  ADDFXL U8 ( .A(n33), .B(n32), .CI(n8), .CO(n7), .S(product_16_) );
  ADDFXL U9 ( .A(n34), .B(n35), .CI(n9), .CO(n8), .S(product_15_) );
  ADDFXL U10 ( .A(n36), .B(n37), .CI(n10), .CO(n9), .S(product_14_) );
  ADDFXL U11 ( .A(n38), .B(n39), .CI(n11), .CO(n10), .S(product_13_) );
  ADDFXL U12 ( .A(n40), .B(n41), .CI(n12), .CO(n11), .S(product_12_) );
  ADDFXL U13 ( .A(n42), .B(n43), .CI(n13), .CO(n12), .S(product_11_) );
  ADDFXL U14 ( .A(n44), .B(n45), .CI(n14), .CO(n13), .S(product_10_) );
  ADDFXL U15 ( .A(n46), .B(n47), .CI(n15), .CO(n14), .S(product_9_) );
  ADDFXL U16 ( .A(n48), .B(n49), .CI(n16), .CO(n15), .S(product_8_) );
  ADDFXL U17 ( .A(n50), .B(a[2]), .CI(n17), .CO(n16), .S(product_7_) );
  ADDFXL U18 ( .A(a[1]), .B(n61), .CI(n18), .CO(n17), .S(product_6_) );
  ADDFXL U19 ( .A(a[0]), .B(n62), .CI(n19), .CO(n18), .S(product_5_) );
  ADDHXL U20 ( .A(n63), .B(n20), .CO(n19), .S(product_4_) );
  ADDHXL U21 ( .A(n64), .B(n21), .CO(n20), .S(product_3_) );
  ADDHXL U22 ( .A(n65), .B(n22), .CO(n21), .S(product_2_) );
  CLKINVX1 U23 ( .A(n22), .Y(product_1_) );
  ADDFXL U24 ( .A(n54), .B(n51), .CI(n53), .CO(n23), .S(n24) );
  ADDFXL U25 ( .A(n55), .B(a[12]), .CI(a[14]), .CO(n25), .S(n26) );
  ADDFXL U26 ( .A(n56), .B(a[11]), .CI(a[13]), .CO(n27), .S(n28) );
  ADDFXL U27 ( .A(n57), .B(a[10]), .CI(a[12]), .CO(n29), .S(n30) );
  ADDFXL U28 ( .A(a[11]), .B(a[9]), .CI(a[15]), .CO(n31), .S(n32) );
  ADDFXL U29 ( .A(n58), .B(n52), .CI(a[10]), .CO(n33), .S(n34) );
  ADDFXL U30 ( .A(n59), .B(n53), .CI(a[9]), .CO(n35), .S(n36) );
  ADDFXL U31 ( .A(n60), .B(n54), .CI(a[8]), .CO(n37), .S(n38) );
  ADDFXL U32 ( .A(n61), .B(n55), .CI(a[7]), .CO(n39), .S(n40) );
  ADDFXL U33 ( .A(n62), .B(n56), .CI(a[6]), .CO(n41), .S(n42) );
  ADDFXL U34 ( .A(n63), .B(n57), .CI(a[5]), .CO(n43), .S(n44) );
  ADDFXL U35 ( .A(n64), .B(n58), .CI(a[4]), .CO(n45), .S(n46) );
  ADDFXL U36 ( .A(n65), .B(n59), .CI(a[3]), .CO(n47), .S(n48) );
  XNOR2X1 U37 ( .A(n22), .B(n60), .Y(n50) );
  OR2X1 U38 ( .A(n22), .B(n60), .Y(n49) );
  CLKINVX1 U59 ( .A(a[15]), .Y(n51) );
  CLKINVX1 U60 ( .A(a[0]), .Y(n22) );
  CLKINVX1 U61 ( .A(a[6]), .Y(n60) );
  CLKINVX1 U62 ( .A(a[13]), .Y(n53) );
  CLKINVX1 U63 ( .A(a[1]), .Y(n65) );
  CLKINVX1 U64 ( .A(a[2]), .Y(n64) );
  CLKINVX1 U65 ( .A(a[3]), .Y(n63) );
  CLKINVX1 U66 ( .A(a[14]), .Y(n52) );
  CLKINVX1 U67 ( .A(a[4]), .Y(n62) );
  CLKINVX1 U68 ( .A(a[5]), .Y(n61) );
  CLKINVX1 U69 ( .A(a[7]), .Y(n59) );
  CLKINVX1 U70 ( .A(a[8]), .Y(n58) );
  CLKINVX1 U71 ( .A(a[9]), .Y(n57) );
  CLKINVX1 U72 ( .A(a[10]), .Y(n56) );
  CLKINVX1 U73 ( .A(a[11]), .Y(n55) );
  CLKINVX1 U74 ( .A(a[12]), .Y(n54) );
endmodule


module FAS_DW_mult_tc_33 ( a, product_28_, product_27_, product_26_, 
        product_25_, product_24_, product_23_, product_22_, product_21_, 
        product_20_, product_19_, product_18_, product_17_, product_16_, 
        product_15_, product_14_, product_13_, product_12_, product_11_, 
        product_10_, product_9_, product_8_, product_7_, product_6_, 
        product_5_, product_4_, product_3_, product_2_, product_1_ );
  input [15:0] a;
  output product_28_, product_27_, product_26_, product_25_, product_24_,
         product_23_, product_22_, product_21_, product_20_, product_19_,
         product_18_, product_17_, product_16_, product_15_, product_14_,
         product_13_, product_12_, product_11_, product_10_, product_9_,
         product_8_, product_7_, product_6_, product_5_, product_4_,
         product_3_, product_2_, product_1_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n114;

  CLKINVX1 U1 ( .A(n2), .Y(product_27_) );
  ADDFXL U3 ( .A(a[15]), .B(n98), .CI(n3), .CO(n2), .S(product_26_) );
  ADDFXL U4 ( .A(n99), .B(a[14]), .CI(n4), .CO(n3), .S(product_25_) );
  ADDFXL U5 ( .A(n28), .B(a[13]), .CI(n5), .CO(n4), .S(product_24_) );
  ADDFXL U6 ( .A(n29), .B(n30), .CI(n6), .CO(n5), .S(product_23_) );
  ADDFXL U7 ( .A(n33), .B(n31), .CI(n7), .CO(n6), .S(product_22_) );
  ADDFXL U8 ( .A(n36), .B(n34), .CI(n8), .CO(n7), .S(product_21_) );
  ADDFXL U9 ( .A(n37), .B(n39), .CI(n9), .CO(n8), .S(product_20_) );
  ADDFXL U10 ( .A(n40), .B(n44), .CI(n10), .CO(n9), .S(product_19_) );
  ADDFXL U11 ( .A(n45), .B(n49), .CI(n11), .CO(n10), .S(product_18_) );
  ADDFXL U12 ( .A(n50), .B(n54), .CI(n12), .CO(n11), .S(product_17_) );
  ADDFXL U13 ( .A(n55), .B(n59), .CI(n13), .CO(n12), .S(product_16_) );
  ADDFXL U14 ( .A(n60), .B(n64), .CI(n14), .CO(n13), .S(product_15_) );
  ADDFXL U15 ( .A(n65), .B(n69), .CI(n15), .CO(n14), .S(product_14_) );
  ADDFXL U16 ( .A(n70), .B(n74), .CI(n16), .CO(n15), .S(product_13_) );
  ADDFXL U17 ( .A(n75), .B(n79), .CI(n17), .CO(n16), .S(product_12_) );
  ADDFXL U18 ( .A(n80), .B(n84), .CI(n18), .CO(n17), .S(product_11_) );
  ADDFXL U19 ( .A(n85), .B(n87), .CI(n19), .CO(n18), .S(product_10_) );
  ADDFXL U20 ( .A(n88), .B(n89), .CI(n20), .CO(n19), .S(product_9_) );
  ADDFXL U21 ( .A(n90), .B(n93), .CI(n21), .CO(n20), .S(product_8_) );
  ADDFXL U22 ( .A(n94), .B(n95), .CI(n22), .CO(n21), .S(product_7_) );
  ADDFXL U23 ( .A(n96), .B(a[0]), .CI(n23), .CO(n22), .S(product_6_) );
  ADDFXL U24 ( .A(a[1]), .B(n108), .CI(n24), .CO(n23), .S(product_5_) );
  ADDFXL U25 ( .A(a[0]), .B(n109), .CI(n25), .CO(n24), .S(product_4_) );
  ADDHXL U26 ( .A(n110), .B(n26), .CO(n25), .S(product_3_) );
  ADDHXL U27 ( .A(n111), .B(n112), .CO(n26), .S(product_2_) );
  CLKINVX1 U28 ( .A(n112), .Y(product_1_) );
  ADDFXL U30 ( .A(n100), .B(n98), .CI(a[15]), .CO(n28), .S(n29) );
  ADDFXL U31 ( .A(n101), .B(a[14]), .CI(n32), .CO(n30), .S(n31) );
  CMPR42X1 U32 ( .A(n102), .B(n100), .C(n99), .D(n97), .ICI(n35), .S(n34), 
        .ICO(n32), .CO(n33) );
  CMPR42X1 U33 ( .A(a[12]), .B(n103), .C(n114), .D(n41), .ICI(n38), .S(n37), 
        .ICO(n35), .CO(n36) );
  CMPR42X1 U34 ( .A(n97), .B(n101), .C(n46), .D(n42), .ICI(n43), .S(n40), 
        .ICO(n38), .CO(n39) );
  ADDFXL U35 ( .A(n102), .B(n104), .CI(a[13]), .CO(n41), .S(n42) );
  CMPR42X1 U36 ( .A(n105), .B(n103), .C(n47), .D(n51), .ICI(n48), .S(n45), 
        .ICO(n43), .CO(n44) );
  ADDFXL U37 ( .A(a[12]), .B(a[10]), .CI(n114), .CO(n46), .S(n47) );
  CMPR42X1 U38 ( .A(n106), .B(n104), .C(n52), .D(n56), .ICI(n53), .S(n50), 
        .ICO(n48), .CO(n49) );
  ADDFXL U39 ( .A(a[11]), .B(a[9]), .CI(a[13]), .CO(n51), .S(n52) );
  CMPR42X1 U40 ( .A(n107), .B(a[15]), .C(n57), .D(n61), .ICI(n58), .S(n55), 
        .ICO(n53), .CO(n54) );
  ADDFXL U41 ( .A(a[12]), .B(a[8]), .CI(a[10]), .CO(n56), .S(n57) );
  CMPR42X1 U42 ( .A(n98), .B(n105), .C(n66), .D(n62), .ICI(n63), .S(n60), 
        .ICO(n58), .CO(n59) );
  ADDFXL U43 ( .A(a[11]), .B(n108), .CI(a[9]), .CO(n61), .S(n62) );
  CMPR42X1 U44 ( .A(n99), .B(n106), .C(n68), .D(n71), .ICI(n67), .S(n65), 
        .ICO(n63), .CO(n64) );
  ADDFXL U45 ( .A(a[10]), .B(n109), .CI(a[8]), .CO(n66), .S(n67) );
  CMPR42X1 U46 ( .A(n100), .B(n107), .C(n73), .D(n76), .ICI(n72), .S(n70), 
        .ICO(n68), .CO(n69) );
  ADDFXL U47 ( .A(a[9]), .B(n110), .CI(a[7]), .CO(n71), .S(n72) );
  CMPR42X1 U48 ( .A(n101), .B(n108), .C(a[6]), .D(n78), .ICI(n77), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFXL U49 ( .A(a[8]), .B(n111), .CI(n81), .CO(n76), .S(n77) );
  CMPR42X1 U50 ( .A(n112), .B(a[5]), .C(a[7]), .D(n82), .ICI(n83), .S(n80), 
        .ICO(n78), .CO(n79) );
  XNOR2X1 U51 ( .A(n102), .B(n109), .Y(n82) );
  OR2X1 U52 ( .A(n102), .B(n109), .Y(n81) );
  CMPR42X1 U53 ( .A(n103), .B(n110), .C(a[4]), .D(a[6]), .ICI(n86), .S(n85), 
        .ICO(n83), .CO(n84) );
  CMPR42X1 U54 ( .A(n104), .B(n111), .C(a[3]), .D(a[5]), .ICI(n91), .S(n88), 
        .ICO(n86), .CO(n87) );
  ADDFXL U55 ( .A(a[2]), .B(a[4]), .CI(n92), .CO(n89), .S(n90) );
  XNOR2X1 U56 ( .A(n105), .B(n112), .Y(n92) );
  OR2X1 U57 ( .A(n105), .B(n112), .Y(n91) );
  ADDFXL U58 ( .A(a[1]), .B(n106), .CI(a[3]), .CO(n93), .S(n94) );
  ADDHXL U59 ( .A(n107), .B(a[2]), .CO(n95), .S(n96) );
  CLKINVX1 U81 ( .A(n2), .Y(product_28_) );
  CLKINVX1 U82 ( .A(a[9]), .Y(n103) );
  CLKINVX1 U83 ( .A(a[0]), .Y(n112) );
  CLKINVX1 U84 ( .A(a[7]), .Y(n105) );
  CLKINVX1 U85 ( .A(a[5]), .Y(n107) );
  CLKINVX1 U86 ( .A(a[6]), .Y(n106) );
  CLKINVX1 U87 ( .A(a[8]), .Y(n104) );
  CLKINVX1 U88 ( .A(a[11]), .Y(n101) );
  CLKINVX1 U89 ( .A(a[12]), .Y(n100) );
  CLKBUFX3 U90 ( .A(a[14]), .Y(n114) );
  CLKINVX1 U91 ( .A(a[13]), .Y(n99) );
  CLKINVX1 U92 ( .A(a[10]), .Y(n102) );
  CLKINVX1 U93 ( .A(a[1]), .Y(n111) );
  CLKINVX1 U94 ( .A(a[2]), .Y(n110) );
  CLKINVX1 U95 ( .A(a[4]), .Y(n108) );
  CLKINVX1 U96 ( .A(a[15]), .Y(n97) );
  CLKINVX1 U97 ( .A(a[14]), .Y(n98) );
  CLKINVX1 U98 ( .A(a[3]), .Y(n109) );
endmodule


module FAS_DW_mult_tc_34 ( a, product );
  input [15:0] a;
  output [25:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103;

  CLKINVX1 U1 ( .A(n89), .Y(product[25]) );
  ADDFXL U3 ( .A(n90), .B(a[15]), .CI(n3), .CO(product[23]), .S(product[22])
         );
  ADDFXL U4 ( .A(n24), .B(n91), .CI(n4), .CO(n3), .S(product[21]) );
  ADDFXL U5 ( .A(n26), .B(n25), .CI(n5), .CO(n4), .S(product[20]) );
  ADDFXL U6 ( .A(n28), .B(n27), .CI(n6), .CO(n5), .S(product[19]) );
  ADDFXL U7 ( .A(n31), .B(n29), .CI(n7), .CO(n6), .S(product[18]) );
  ADDFXL U8 ( .A(n34), .B(n32), .CI(n8), .CO(n7), .S(product[17]) );
  ADDFXL U9 ( .A(n37), .B(n35), .CI(n9), .CO(n8), .S(product[16]) );
  ADDFXL U10 ( .A(n38), .B(n42), .CI(n10), .CO(n9), .S(product[15]) );
  ADDFXL U11 ( .A(n43), .B(n47), .CI(n11), .CO(n10), .S(product[14]) );
  ADDFXL U12 ( .A(n48), .B(n52), .CI(n12), .CO(n11), .S(product[13]) );
  ADDFXL U13 ( .A(n53), .B(n57), .CI(n13), .CO(n12), .S(product[12]) );
  ADDFXL U14 ( .A(n58), .B(n62), .CI(n14), .CO(n13), .S(product[11]) );
  ADDFXL U15 ( .A(n63), .B(n67), .CI(n15), .CO(n14), .S(product[10]) );
  ADDFXL U16 ( .A(n68), .B(n72), .CI(n16), .CO(n15), .S(product[9]) );
  ADDFXL U17 ( .A(n73), .B(n77), .CI(n17), .CO(n16), .S(product[8]) );
  ADDFXL U18 ( .A(n78), .B(n79), .CI(n18), .CO(n17), .S(product[7]) );
  ADDFXL U19 ( .A(n80), .B(n83), .CI(n19), .CO(n18), .S(product[6]) );
  ADDFXL U20 ( .A(n84), .B(n85), .CI(n20), .CO(n19), .S(product[5]) );
  ADDFXL U21 ( .A(n86), .B(n87), .CI(n21), .CO(n20), .S(product[4]) );
  ADDFXL U22 ( .A(n88), .B(product[0]), .CI(n22), .CO(n21), .S(product[3]) );
  ADDFXL U23 ( .A(n102), .B(n103), .CI(n23), .CO(n22), .S(product[2]) );
  ADDHXL U24 ( .A(product[0]), .B(n103), .CO(n23), .S(product[1]) );
  ADDFXL U25 ( .A(n92), .B(a[15]), .CI(n90), .CO(n24), .S(n25) );
  ADDFXL U26 ( .A(n93), .B(a[15]), .CI(n91), .CO(n26), .S(n27) );
  ADDFXL U27 ( .A(n94), .B(n92), .CI(n30), .CO(n28), .S(n29) );
  CMPR42X1 U28 ( .A(a[15]), .B(n90), .C(n95), .D(n93), .ICI(n33), .S(n32), 
        .ICO(n30), .CO(n31) );
  CMPR42X1 U29 ( .A(n91), .B(n96), .C(n94), .D(n39), .ICI(n36), .S(n35), .ICO(
        n33), .CO(n34) );
  CMPR42X1 U30 ( .A(n90), .B(n92), .C(n40), .D(n44), .ICI(n41), .S(n38), .ICO(
        n36), .CO(n37) );
  ADDFXL U31 ( .A(n97), .B(a[15]), .CI(n95), .CO(n39), .S(n40) );
  CMPR42X1 U32 ( .A(n90), .B(n91), .C(n49), .D(n45), .ICI(n46), .S(n43), .ICO(
        n41), .CO(n42) );
  ADDFXL U33 ( .A(n98), .B(n96), .CI(n93), .CO(n44), .S(n45) );
  CMPR42X1 U34 ( .A(n91), .B(n92), .C(n54), .D(n50), .ICI(n51), .S(n48), .ICO(
        n46), .CO(n47) );
  ADDFXL U35 ( .A(n99), .B(n97), .CI(n94), .CO(n49), .S(n50) );
  CMPR42X1 U36 ( .A(n92), .B(n93), .C(n59), .D(n55), .ICI(n56), .S(n53), .ICO(
        n51), .CO(n52) );
  ADDFXL U37 ( .A(n100), .B(n98), .CI(n95), .CO(n54), .S(n55) );
  CMPR42X1 U38 ( .A(n93), .B(n94), .C(n61), .D(n64), .ICI(n60), .S(n58), .ICO(
        n56), .CO(n57) );
  ADDFXL U39 ( .A(n101), .B(n99), .CI(n96), .CO(n59), .S(n60) );
  CMPR42X1 U40 ( .A(n94), .B(n95), .C(n66), .D(n69), .ICI(n65), .S(n63), .ICO(
        n61), .CO(n62) );
  ADDFXL U41 ( .A(n102), .B(n100), .CI(n97), .CO(n64), .S(n65) );
  CMPR42X1 U42 ( .A(n95), .B(n98), .C(n96), .D(n71), .ICI(n70), .S(n68), .ICO(
        n66), .CO(n67) );
  ADDFXL U43 ( .A(n103), .B(n101), .CI(n74), .CO(n69), .S(n70) );
  CMPR42X1 U44 ( .A(n96), .B(n99), .C(n97), .D(n75), .ICI(n76), .S(n73), .ICO(
        n71), .CO(n72) );
  ADDHXL U45 ( .A(n102), .B(product[0]), .CO(n74), .S(n75) );
  CMPR42X1 U46 ( .A(n100), .B(n103), .C(n98), .D(n97), .ICI(n81), .S(n78), 
        .ICO(n76), .CO(n77) );
  ADDFXL U47 ( .A(n99), .B(n98), .CI(n82), .CO(n79), .S(n80) );
  ADDHXL U48 ( .A(n101), .B(product[0]), .CO(n81), .S(n82) );
  ADDFXL U49 ( .A(n102), .B(n99), .CI(n100), .CO(n83), .S(n84) );
  ADDFXL U50 ( .A(n103), .B(n100), .CI(n101), .CO(n85), .S(n86) );
  ADDHXL U51 ( .A(n101), .B(n102), .CO(n87), .S(n88) );
  CLKINVX1 U72 ( .A(a[15]), .Y(n89) );
  CLKBUFX3 U73 ( .A(a[0]), .Y(product[0]) );
  CLKBUFX3 U74 ( .A(a[9]), .Y(n95) );
  CLKBUFX3 U75 ( .A(a[13]), .Y(n91) );
  CLKBUFX3 U76 ( .A(a[14]), .Y(n90) );
  CLKBUFX3 U77 ( .A(a[8]), .Y(n96) );
  CLKBUFX3 U78 ( .A(a[12]), .Y(n92) );
  CLKBUFX3 U79 ( .A(a[10]), .Y(n94) );
  CLKBUFX3 U80 ( .A(a[11]), .Y(n93) );
  CLKBUFX3 U81 ( .A(a[6]), .Y(n98) );
  CLKBUFX3 U82 ( .A(a[7]), .Y(n97) );
  CLKBUFX3 U83 ( .A(a[1]), .Y(n103) );
  CLKBUFX3 U84 ( .A(a[4]), .Y(n100) );
  CLKBUFX3 U85 ( .A(a[5]), .Y(n99) );
  CLKBUFX3 U86 ( .A(a[3]), .Y(n101) );
  CLKBUFX3 U87 ( .A(a[2]), .Y(n102) );
  BUFX2 U88 ( .A(product[25]), .Y(product[24]) );
endmodule


module FAS_DW_mult_tc_35 ( a, product );
  input [15:0] a;
  output [23:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83;

  CLKINVX1 U1 ( .A(n1), .Y(product[23]) );
  ADDFXL U2 ( .A(a[15]), .B(n70), .CI(n2), .CO(n1), .S(product[22]) );
  ADDFXL U3 ( .A(n24), .B(a[14]), .CI(n3), .CO(n2), .S(product[21]) );
  ADDFXL U4 ( .A(n25), .B(n26), .CI(n4), .CO(n3), .S(product[20]) );
  ADDFXL U5 ( .A(n29), .B(n27), .CI(n5), .CO(n4), .S(product[19]) );
  ADDFXL U6 ( .A(n30), .B(n32), .CI(n6), .CO(n5), .S(product[18]) );
  ADDFXL U7 ( .A(n33), .B(n35), .CI(n7), .CO(n6), .S(product[17]) );
  ADDFXL U8 ( .A(n36), .B(n38), .CI(n8), .CO(n7), .S(product[16]) );
  ADDFXL U9 ( .A(n39), .B(n41), .CI(n9), .CO(n8), .S(product[15]) );
  ADDFXL U10 ( .A(n42), .B(n44), .CI(n10), .CO(n9), .S(product[14]) );
  ADDFXL U11 ( .A(n45), .B(n47), .CI(n11), .CO(n10), .S(product[13]) );
  ADDFXL U12 ( .A(n48), .B(n50), .CI(n12), .CO(n11), .S(product[12]) );
  ADDFXL U13 ( .A(n51), .B(n53), .CI(n13), .CO(n12), .S(product[11]) );
  ADDFXL U14 ( .A(n54), .B(n56), .CI(n14), .CO(n13), .S(product[10]) );
  ADDFXL U15 ( .A(n57), .B(n59), .CI(n15), .CO(n14), .S(product[9]) );
  ADDFXL U16 ( .A(n60), .B(n61), .CI(n16), .CO(n15), .S(product[8]) );
  ADDFXL U17 ( .A(n62), .B(n65), .CI(n17), .CO(n16), .S(product[7]) );
  ADDFXL U18 ( .A(n66), .B(n67), .CI(n18), .CO(n17), .S(product[6]) );
  ADDFXL U19 ( .A(n68), .B(a[0]), .CI(n19), .CO(n18), .S(product[5]) );
  ADDFXL U20 ( .A(a[1]), .B(n80), .CI(n20), .CO(n19), .S(product[4]) );
  ADDFXL U21 ( .A(a[0]), .B(n81), .CI(n21), .CO(n20), .S(product[3]) );
  ADDHXL U22 ( .A(n82), .B(n22), .CO(n21), .S(product[2]) );
  ADDHXL U23 ( .A(n83), .B(n23), .CO(n22), .S(product[1]) );
  CLKINVX1 U24 ( .A(n23), .Y(product[0]) );
  ADDFXL U25 ( .A(n72), .B(n69), .CI(n71), .CO(n24), .S(n25) );
  ADDFXL U26 ( .A(a[14]), .B(a[12]), .CI(n28), .CO(n26), .S(n27) );
  CMPR42X1 U27 ( .A(n73), .B(n74), .C(n69), .D(a[13]), .ICI(n31), .S(n30), 
        .ICO(n28), .CO(n29) );
  CMPR42X1 U28 ( .A(a[10]), .B(n75), .C(a[12]), .D(a[14]), .ICI(n34), .S(n33), 
        .ICO(n31), .CO(n32) );
  CMPR42X1 U29 ( .A(a[9]), .B(n76), .C(a[11]), .D(a[13]), .ICI(n37), .S(n36), 
        .ICO(n34), .CO(n35) );
  CMPR42X1 U30 ( .A(a[8]), .B(a[15]), .C(a[10]), .D(a[12]), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U31 ( .A(n70), .B(n77), .C(a[9]), .D(a[11]), .ICI(n43), .S(n42), 
        .ICO(n40), .CO(n41) );
  CMPR42X1 U32 ( .A(n71), .B(n78), .C(a[8]), .D(a[10]), .ICI(n46), .S(n45), 
        .ICO(n43), .CO(n44) );
  CMPR42X1 U33 ( .A(n72), .B(n79), .C(a[7]), .D(a[9]), .ICI(n49), .S(n48), 
        .ICO(n46), .CO(n47) );
  CMPR42X1 U34 ( .A(n73), .B(n80), .C(a[6]), .D(a[8]), .ICI(n52), .S(n51), 
        .ICO(n49), .CO(n50) );
  CMPR42X1 U35 ( .A(n74), .B(n81), .C(a[5]), .D(a[7]), .ICI(n55), .S(n54), 
        .ICO(n52), .CO(n53) );
  CMPR42X1 U36 ( .A(n75), .B(n82), .C(a[4]), .D(a[6]), .ICI(n58), .S(n57), 
        .ICO(n55), .CO(n56) );
  CMPR42X1 U37 ( .A(n76), .B(n83), .C(a[3]), .D(a[5]), .ICI(n63), .S(n60), 
        .ICO(n58), .CO(n59) );
  ADDFXL U38 ( .A(a[2]), .B(a[4]), .CI(n64), .CO(n61), .S(n62) );
  XNOR2X1 U39 ( .A(n77), .B(n23), .Y(n64) );
  OR2X1 U40 ( .A(n77), .B(n23), .Y(n63) );
  ADDFXL U41 ( .A(a[1]), .B(n78), .CI(a[3]), .CO(n65), .S(n66) );
  ADDHXL U42 ( .A(n79), .B(a[2]), .CO(n67), .S(n68) );
  CLKINVX1 U63 ( .A(a[8]), .Y(n76) );
  CLKINVX1 U64 ( .A(a[9]), .Y(n75) );
  CLKINVX1 U65 ( .A(a[10]), .Y(n74) );
  CLKINVX1 U66 ( .A(a[11]), .Y(n73) );
  CLKINVX1 U67 ( .A(a[7]), .Y(n77) );
  CLKINVX1 U68 ( .A(a[0]), .Y(n23) );
  CLKINVX1 U69 ( .A(a[13]), .Y(n71) );
  CLKINVX1 U70 ( .A(a[1]), .Y(n83) );
  CLKINVX1 U71 ( .A(a[2]), .Y(n82) );
  CLKINVX1 U72 ( .A(a[5]), .Y(n79) );
  CLKINVX1 U73 ( .A(a[3]), .Y(n81) );
  CLKINVX1 U74 ( .A(a[4]), .Y(n80) );
  CLKINVX1 U75 ( .A(a[6]), .Y(n78) );
  CLKINVX1 U76 ( .A(a[14]), .Y(n70) );
  CLKINVX1 U77 ( .A(a[12]), .Y(n72) );
  CLKINVX1 U78 ( .A(a[15]), .Y(n69) );
endmodule


module FAS_DW_mult_tc_36 ( a, product_26_, product_25_, product_24_, 
        product_23_, product_22_, product_21_, product_20_, product_19_, 
        product_18_, product_17_, product_16_, product_15_, product_14_, 
        product_13_, product_12_, product_11_, product_10_, product_9_, 
        product_8_, product_7_, product_6_, product_5_, product_4_, product_3_, 
        product_2_ );
  input [15:0] a;
  output product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83;

  CLKINVX1 U3 ( .A(n2), .Y(product_25_) );
  ADDFXL U4 ( .A(n83), .B(n68), .CI(n3), .CO(n2), .S(product_24_) );
  ADDFXL U5 ( .A(n23), .B(a[14]), .CI(n4), .CO(n3), .S(product_23_) );
  ADDFXL U6 ( .A(n24), .B(n25), .CI(n5), .CO(n4), .S(product_22_) );
  ADDFXL U7 ( .A(n27), .B(n26), .CI(n6), .CO(n5), .S(product_21_) );
  ADDFXL U8 ( .A(n30), .B(n28), .CI(n7), .CO(n6), .S(product_20_) );
  ADDFXL U9 ( .A(n31), .B(n33), .CI(n8), .CO(n7), .S(product_19_) );
  ADDFXL U10 ( .A(n34), .B(n36), .CI(n9), .CO(n8), .S(product_18_) );
  ADDFXL U11 ( .A(n37), .B(n39), .CI(n10), .CO(n9), .S(product_17_) );
  ADDFXL U12 ( .A(n40), .B(n42), .CI(n11), .CO(n10), .S(product_16_) );
  ADDFXL U13 ( .A(n43), .B(n45), .CI(n12), .CO(n11), .S(product_15_) );
  ADDFXL U14 ( .A(n46), .B(n48), .CI(n13), .CO(n12), .S(product_14_) );
  ADDFXL U15 ( .A(n49), .B(n51), .CI(n14), .CO(n13), .S(product_13_) );
  ADDFXL U16 ( .A(n52), .B(n54), .CI(n15), .CO(n14), .S(product_12_) );
  ADDFXL U17 ( .A(n55), .B(n57), .CI(n16), .CO(n15), .S(product_11_) );
  ADDFXL U18 ( .A(n58), .B(n59), .CI(n17), .CO(n16), .S(product_10_) );
  ADDFXL U19 ( .A(n60), .B(n63), .CI(n18), .CO(n17), .S(product_9_) );
  ADDFXL U20 ( .A(n64), .B(n65), .CI(n19), .CO(n18), .S(product_8_) );
  ADDFXL U21 ( .A(n66), .B(a[5]), .CI(n20), .CO(n19), .S(product_7_) );
  ADDFXL U22 ( .A(a[4]), .B(n80), .CI(n21), .CO(n20), .S(product_6_) );
  ADDFXL U23 ( .A(a[3]), .B(n81), .CI(n22), .CO(n21), .S(product_5_) );
  XNOR2X1 U24 ( .A(a[2]), .B(n82), .Y(product_4_) );
  OR2X1 U25 ( .A(a[2]), .B(n82), .Y(n22) );
  ADDFXL U26 ( .A(n69), .B(n68), .CI(n83), .CO(n23), .S(n24) );
  ADDFXL U27 ( .A(n69), .B(a[14]), .CI(n70), .CO(n25), .S(n26) );
  ADDFXL U28 ( .A(n71), .B(a[13]), .CI(n29), .CO(n27), .S(n28) );
  CMPR42X1 U29 ( .A(n68), .B(n72), .C(n70), .D(n83), .ICI(n32), .S(n31), .ICO(
        n29), .CO(n30) );
  CMPR42X1 U30 ( .A(a[14]), .B(n67), .C(n73), .D(n71), .ICI(n35), .S(n34), 
        .ICO(n32), .CO(n33) );
  CMPR42X1 U31 ( .A(a[15]), .B(n74), .C(n72), .D(n69), .ICI(n38), .S(n37), 
        .ICO(n35), .CO(n36) );
  CMPR42X1 U32 ( .A(n75), .B(n73), .C(n70), .D(a[14]), .ICI(n41), .S(n40), 
        .ICO(n38), .CO(n39) );
  CMPR42X1 U33 ( .A(n76), .B(n74), .C(n71), .D(a[13]), .ICI(n44), .S(n43), 
        .ICO(n41), .CO(n42) );
  CMPR42X1 U34 ( .A(n77), .B(n75), .C(n72), .D(a[12]), .ICI(n47), .S(n46), 
        .ICO(n44), .CO(n45) );
  CMPR42X1 U35 ( .A(n78), .B(n76), .C(n73), .D(a[11]), .ICI(n50), .S(n49), 
        .ICO(n47), .CO(n48) );
  CMPR42X1 U36 ( .A(n79), .B(n77), .C(n74), .D(a[10]), .ICI(n53), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U37 ( .A(n80), .B(n78), .C(n75), .D(a[9]), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U38 ( .A(n81), .B(n79), .C(n76), .D(a[8]), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  ADDFXL U39 ( .A(a[7]), .B(n77), .CI(n62), .CO(n59), .S(n60) );
  XNOR2X1 U40 ( .A(n80), .B(n82), .Y(n62) );
  OR2X1 U41 ( .A(n80), .B(n82), .Y(n61) );
  ADDFXL U42 ( .A(n78), .B(n81), .CI(a[6]), .CO(n63), .S(n64) );
  XNOR2X1 U43 ( .A(n79), .B(n82), .Y(n66) );
  OR2X1 U44 ( .A(n79), .B(n82), .Y(n65) );
  CLKBUFX3 U69 ( .A(product_25_), .Y(product_26_) );
  CLKBUFX3 U70 ( .A(a[0]), .Y(product_2_) );
  CLKINVX1 U71 ( .A(a[15]), .Y(n67) );
  CLKBUFX3 U72 ( .A(a[1]), .Y(product_3_) );
  CLKINVX1 U73 ( .A(a[8]), .Y(n74) );
  CLKINVX1 U74 ( .A(a[6]), .Y(n76) );
  CLKINVX1 U75 ( .A(a[7]), .Y(n75) );
  CLKINVX1 U76 ( .A(a[9]), .Y(n73) );
  CLKINVX1 U77 ( .A(a[10]), .Y(n72) );
  CLKINVX1 U78 ( .A(a[3]), .Y(n79) );
  CLKINVX1 U79 ( .A(a[5]), .Y(n77) );
  CLKINVX1 U80 ( .A(a[4]), .Y(n78) );
  CLKBUFX3 U81 ( .A(a[15]), .Y(n83) );
  CLKINVX1 U82 ( .A(a[12]), .Y(n70) );
  CLKINVX1 U83 ( .A(a[0]), .Y(n82) );
  CLKINVX1 U84 ( .A(a[2]), .Y(n80) );
  CLKINVX1 U85 ( .A(a[11]), .Y(n71) );
  CLKINVX1 U86 ( .A(a[1]), .Y(n81) );
  CLKINVX1 U87 ( .A(a[14]), .Y(n68) );
  CLKINVX1 U88 ( .A(a[13]), .Y(n69) );
endmodule


module FAS_DW_mult_tc_37 ( a, product_30_, product_29_, product_28_, 
        product_27_, product_26_, product_25_, product_24_, product_23_, 
        product_22_, product_21_, product_20_, product_19_, product_18_, 
        product_17_, product_16_, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_, product_2_, 
        product_1_ );
  input [15:0] a;
  output product_30_, product_29_, product_28_, product_27_, product_26_,
         product_25_, product_24_, product_23_, product_22_, product_21_,
         product_20_, product_19_, product_18_, product_17_, product_16_,
         product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_, product_2_, product_1_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n33,
         n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n112, n114, n115, n116,
         n117;

  CLKINVX1 U1 ( .A(n2), .Y(product_29_) );
  ADDFXL U3 ( .A(n112), .B(n96), .CI(n3), .CO(n2), .S(product_28_) );
  ADDFXL U4 ( .A(a[13]), .B(n96), .CI(n4), .CO(n3), .S(product_27_) );
  ADDFXL U5 ( .A(n97), .B(n114), .CI(n5), .CO(n4), .S(product_26_) );
  ADDFXL U6 ( .A(n98), .B(n115), .CI(n6), .CO(n5), .S(product_25_) );
  ADDFXL U7 ( .A(n33), .B(n99), .CI(n7), .CO(n6), .S(product_24_) );
  ADDFXL U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product_23_) );
  ADDFXL U9 ( .A(n40), .B(n38), .CI(n9), .CO(n8), .S(product_22_) );
  ADDFXL U10 ( .A(n41), .B(n43), .CI(n10), .CO(n9), .S(product_21_) );
  ADDFXL U11 ( .A(n44), .B(n48), .CI(n11), .CO(n10), .S(product_20_) );
  ADDFXL U12 ( .A(n49), .B(n53), .CI(n12), .CO(n11), .S(product_19_) );
  ADDFXL U13 ( .A(n54), .B(n58), .CI(n13), .CO(n12), .S(product_18_) );
  ADDFXL U14 ( .A(n59), .B(n63), .CI(n14), .CO(n13), .S(product_17_) );
  ADDFXL U15 ( .A(n64), .B(n68), .CI(n15), .CO(n14), .S(product_16_) );
  ADDFXL U16 ( .A(n69), .B(n73), .CI(n16), .CO(n15), .S(product_15_) );
  ADDFXL U17 ( .A(n74), .B(n78), .CI(n17), .CO(n16), .S(product_14_) );
  ADDFXL U18 ( .A(n79), .B(n82), .CI(n18), .CO(n17), .S(product_13_) );
  ADDFXL U19 ( .A(n83), .B(n86), .CI(n19), .CO(n18), .S(product_12_) );
  ADDFXL U20 ( .A(n87), .B(n88), .CI(n20), .CO(n19), .S(product_11_) );
  ADDFXL U21 ( .A(n89), .B(n90), .CI(n21), .CO(n20), .S(product_10_) );
  ADDFXL U22 ( .A(n91), .B(n92), .CI(n22), .CO(n21), .S(product_9_) );
  ADDFXL U23 ( .A(n93), .B(n94), .CI(n23), .CO(n22), .S(product_8_) );
  ADDFXL U24 ( .A(n95), .B(a[2]), .CI(n24), .CO(n23), .S(product_7_) );
  ADDFXL U25 ( .A(a[1]), .B(n106), .CI(n25), .CO(n24), .S(product_6_) );
  ADDFXL U26 ( .A(a[0]), .B(n107), .CI(n26), .CO(n25), .S(product_5_) );
  ADDHXL U27 ( .A(n108), .B(n27), .CO(n26), .S(product_4_) );
  ADDHXL U28 ( .A(n109), .B(n28), .CO(n27), .S(product_3_) );
  ADDHXL U29 ( .A(n110), .B(n29), .CO(n28), .S(product_2_) );
  CLKINVX1 U30 ( .A(n29), .Y(product_1_) );
  ADDFXL U34 ( .A(n100), .B(n116), .CI(n36), .CO(n33), .S(n34) );
  CMPR42X1 U36 ( .A(n97), .B(n117), .C(n116), .D(a[15]), .ICI(n39), .S(n38), 
        .ICO(n36), .CO(n37) );
  CMPR42X1 U37 ( .A(a[14]), .B(n117), .C(a[8]), .D(n45), .ICI(n42), .S(n41), 
        .ICO(n39), .CO(n40) );
  CMPR42X1 U38 ( .A(n96), .B(n98), .C(n50), .D(n46), .ICI(n47), .S(n44), .ICO(
        n42), .CO(n43) );
  ADDFXL U39 ( .A(a[8]), .B(n99), .CI(a[7]), .CO(n45), .S(n46) );
  CMPR42X1 U40 ( .A(n100), .B(n112), .C(n51), .D(n55), .ICI(n52), .S(n49), 
        .ICO(n47), .CO(n48) );
  ADDFXL U41 ( .A(a[7]), .B(a[12]), .CI(a[6]), .CO(n50), .S(n51) );
  CMPR42X1 U42 ( .A(n101), .B(a[13]), .C(n56), .D(n60), .ICI(n57), .S(n54), 
        .ICO(n52), .CO(n53) );
  ADDFXL U43 ( .A(a[6]), .B(a[11]), .CI(a[5]), .CO(n55), .S(n56) );
  CMPR42X1 U44 ( .A(n102), .B(n114), .C(n61), .D(n65), .ICI(n62), .S(n59), 
        .ICO(n57), .CO(n58) );
  ADDFXL U45 ( .A(a[5]), .B(a[10]), .CI(a[4]), .CO(n60), .S(n61) );
  CMPR42X1 U46 ( .A(a[15]), .B(n115), .C(n67), .D(n66), .ICI(n70), .S(n64), 
        .ICO(n62), .CO(n63) );
  ADDFXL U47 ( .A(a[3]), .B(a[9]), .CI(a[4]), .CO(n65), .S(n66) );
  CMPR42X1 U48 ( .A(n103), .B(n116), .C(n72), .D(n75), .ICI(n71), .S(n69), 
        .ICO(n67), .CO(n68) );
  ADDFXL U49 ( .A(a[2]), .B(n97), .CI(a[3]), .CO(n70), .S(n71) );
  CMPR42X1 U50 ( .A(n104), .B(a[2]), .C(n117), .D(n77), .ICI(n76), .S(n74), 
        .ICO(n72), .CO(n73) );
  ADDFXL U51 ( .A(a[1]), .B(n98), .CI(n80), .CO(n75), .S(n76) );
  CMPR42X1 U52 ( .A(a[8]), .B(a[0]), .C(a[1]), .D(n84), .ICI(n81), .S(n79), 
        .ICO(n77), .CO(n78) );
  ADDHXL U53 ( .A(n99), .B(n105), .CO(n80), .S(n81) );
  ADDFXL U54 ( .A(a[0]), .B(a[7]), .CI(n85), .CO(n82), .S(n83) );
  ADDHXL U55 ( .A(n100), .B(n106), .CO(n84), .S(n85) );
  ADDFXL U56 ( .A(n107), .B(n101), .CI(a[6]), .CO(n86), .S(n87) );
  ADDFXL U57 ( .A(n108), .B(n102), .CI(a[5]), .CO(n88), .S(n89) );
  ADDFXL U58 ( .A(n109), .B(n103), .CI(a[4]), .CO(n90), .S(n91) );
  ADDFXL U59 ( .A(n110), .B(n104), .CI(a[3]), .CO(n92), .S(n93) );
  XNOR2X1 U60 ( .A(n29), .B(n105), .Y(n95) );
  OR2X1 U61 ( .A(n29), .B(n105), .Y(n94) );
  CLKINVX1 U87 ( .A(n2), .Y(product_30_) );
  CLKBUFX3 U88 ( .A(a[9]), .Y(n117) );
  CLKBUFX3 U89 ( .A(a[10]), .Y(n116) );
  CLKBUFX3 U90 ( .A(a[11]), .Y(n115) );
  CLKBUFX3 U91 ( .A(a[12]), .Y(n114) );
  CLKBUFX3 U92 ( .A(a[14]), .Y(n112) );
  CLKINVX1 U93 ( .A(a[13]), .Y(n98) );
  CLKINVX1 U94 ( .A(a[15]), .Y(n96) );
  CLKINVX1 U95 ( .A(a[0]), .Y(n29) );
  CLKINVX1 U96 ( .A(a[11]), .Y(n100) );
  CLKINVX1 U97 ( .A(a[7]), .Y(n104) );
  CLKINVX1 U98 ( .A(a[8]), .Y(n103) );
  CLKINVX1 U99 ( .A(a[9]), .Y(n102) );
  CLKINVX1 U100 ( .A(a[10]), .Y(n101) );
  CLKINVX1 U101 ( .A(a[14]), .Y(n97) );
  CLKINVX1 U102 ( .A(a[6]), .Y(n105) );
  CLKINVX1 U103 ( .A(a[5]), .Y(n106) );
  CLKINVX1 U104 ( .A(a[12]), .Y(n99) );
  CLKINVX1 U105 ( .A(a[1]), .Y(n110) );
  CLKINVX1 U106 ( .A(a[2]), .Y(n109) );
  CLKINVX1 U107 ( .A(a[3]), .Y(n108) );
  CLKINVX1 U108 ( .A(a[4]), .Y(n107) );
endmodule


module FAS_DW_mult_tc_38 ( a, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_ );
  input [15:0] a;
  output product_29_, product_28_, product_27_, product_26_, product_25_,
         product_24_, product_23_, product_22_, product_21_, product_20_,
         product_19_, product_18_, product_17_, product_16_, product_15_,
         product_14_, product_13_, product_12_, product_11_, product_10_,
         product_9_, product_8_, product_7_, product_6_, product_5_,
         product_4_, product_3_, product_2_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127;

  CLKINVX1 U1 ( .A(n1), .Y(product_29_) );
  ADDFXL U2 ( .A(a[14]), .B(n111), .CI(n2), .CO(n1), .S(product_28_) );
  ADDFXL U3 ( .A(n112), .B(a[13]), .CI(n3), .CO(n2), .S(product_27_) );
  ADDFXL U4 ( .A(n113), .B(a[12]), .CI(n4), .CO(n3), .S(product_26_) );
  ADDFXL U5 ( .A(n34), .B(n114), .CI(n5), .CO(n4), .S(product_25_) );
  ADDFXL U6 ( .A(n35), .B(n36), .CI(n6), .CO(n5), .S(product_24_) );
  ADDFXL U7 ( .A(n38), .B(n37), .CI(n7), .CO(n6), .S(product_23_) );
  ADDFXL U8 ( .A(n41), .B(n39), .CI(n8), .CO(n7), .S(product_22_) );
  ADDFXL U9 ( .A(n44), .B(n42), .CI(n9), .CO(n8), .S(product_21_) );
  ADDFXL U10 ( .A(n45), .B(n47), .CI(n10), .CO(n9), .S(product_20_) );
  ADDFXL U11 ( .A(n48), .B(n52), .CI(n11), .CO(n10), .S(product_19_) );
  ADDFXL U12 ( .A(n53), .B(n57), .CI(n12), .CO(n11), .S(product_18_) );
  ADDFXL U13 ( .A(n58), .B(n62), .CI(n13), .CO(n12), .S(product_17_) );
  ADDFXL U14 ( .A(n63), .B(n67), .CI(n14), .CO(n13), .S(product_16_) );
  ADDFXL U15 ( .A(n68), .B(n72), .CI(n15), .CO(n14), .S(product_15_) );
  ADDFXL U16 ( .A(n73), .B(n77), .CI(n16), .CO(n15), .S(product_14_) );
  ADDFXL U17 ( .A(n78), .B(n82), .CI(n17), .CO(n16), .S(product_13_) );
  ADDFXL U18 ( .A(n83), .B(n87), .CI(n18), .CO(n17), .S(product_12_) );
  ADDFXL U19 ( .A(n88), .B(n92), .CI(n19), .CO(n18), .S(product_11_) );
  ADDFXL U20 ( .A(n93), .B(n97), .CI(n20), .CO(n19), .S(product_10_) );
  ADDFXL U21 ( .A(n98), .B(n99), .CI(n21), .CO(n20), .S(product_9_) );
  ADDFXL U22 ( .A(n100), .B(n103), .CI(n22), .CO(n21), .S(product_8_) );
  ADDFXL U23 ( .A(n104), .B(n107), .CI(n23), .CO(n22), .S(product_7_) );
  ADDFXL U24 ( .A(n108), .B(n109), .CI(n24), .CO(n23), .S(product_6_) );
  ADDFXL U25 ( .A(n110), .B(n124), .CI(n25), .CO(n24), .S(product_5_) );
  ADDFXL U26 ( .A(n126), .B(a[2]), .CI(n26), .CO(n25), .S(product_4_) );
  ADDHXL U27 ( .A(n125), .B(n126), .CO(n26), .S(product_3_) );
  CLKINVX1 U28 ( .A(n126), .Y(product_2_) );
  ADDFXL U33 ( .A(a[11]), .B(n112), .CI(n127), .CO(n34), .S(n35) );
  ADDFXL U34 ( .A(n113), .B(a[14]), .CI(a[10]), .CO(n36), .S(n37) );
  ADDFXL U35 ( .A(a[9]), .B(a[13]), .CI(n40), .CO(n38), .S(n39) );
  CMPR42X1 U36 ( .A(n112), .B(n114), .C(a[8]), .D(n127), .ICI(n43), .S(n42), 
        .ICO(n40), .CO(n41) );
  CMPR42X1 U37 ( .A(a[14]), .B(n115), .C(a[7]), .D(n49), .ICI(n46), .S(n45), 
        .ICO(n43), .CO(n44) );
  CMPR42X1 U38 ( .A(n113), .B(n116), .C(n54), .D(n50), .ICI(n51), .S(n48), 
        .ICO(n46), .CO(n47) );
  ADDFXL U39 ( .A(a[6]), .B(n112), .CI(n127), .CO(n49), .S(n50) );
  CMPR42X1 U40 ( .A(n114), .B(n117), .C(n55), .D(n59), .ICI(n56), .S(n53), 
        .ICO(n51), .CO(n52) );
  ADDFXL U41 ( .A(n113), .B(a[14]), .CI(a[5]), .CO(n54), .S(n55) );
  CMPR42X1 U42 ( .A(n115), .B(n118), .C(n60), .D(n64), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  ADDFXL U43 ( .A(a[4]), .B(a[13]), .CI(n127), .CO(n59), .S(n60) );
  CMPR42X1 U44 ( .A(n114), .B(n116), .C(n69), .D(n65), .ICI(n66), .S(n63), 
        .ICO(n61), .CO(n62) );
  ADDFXL U45 ( .A(n119), .B(n112), .CI(a[3]), .CO(n64), .S(n65) );
  CMPR42X1 U46 ( .A(n115), .B(n117), .C(n71), .D(n74), .ICI(n70), .S(n68), 
        .ICO(n66), .CO(n67) );
  ADDFXL U47 ( .A(n120), .B(n113), .CI(a[2]), .CO(n69), .S(n70) );
  CMPR42X1 U48 ( .A(n116), .B(n118), .C(n76), .D(n79), .ICI(n75), .S(n73), 
        .ICO(n71), .CO(n72) );
  ADDFXL U49 ( .A(n121), .B(n114), .CI(a[1]), .CO(n74), .S(n75) );
  CMPR42X1 U50 ( .A(n117), .B(n122), .C(n119), .D(n81), .ICI(n80), .S(n78), 
        .ICO(n76), .CO(n77) );
  ADDFXL U51 ( .A(a[0]), .B(n115), .CI(n84), .CO(n79), .S(n80) );
  CMPR42X1 U52 ( .A(n116), .B(n118), .C(n89), .D(n85), .ICI(n86), .S(n83), 
        .ICO(n81), .CO(n82) );
  ADDHXL U53 ( .A(n120), .B(n123), .CO(n84), .S(n85) );
  CMPR42X1 U54 ( .A(n117), .B(n119), .C(n94), .D(n90), .ICI(n91), .S(n88), 
        .ICO(n86), .CO(n87) );
  ADDHXL U55 ( .A(n121), .B(n124), .CO(n89), .S(n90) );
  CMPR42X1 U56 ( .A(n118), .B(n122), .C(n120), .D(n96), .ICI(n95), .S(n93), 
        .ICO(n91), .CO(n92) );
  ADDHXL U57 ( .A(n125), .B(n119), .CO(n94), .S(n95) );
  CMPR42X1 U58 ( .A(a[7]), .B(n126), .C(n123), .D(n121), .ICI(n101), .S(n98), 
        .ICO(n96), .CO(n97) );
  ADDFXL U59 ( .A(n105), .B(n122), .CI(n102), .CO(n99), .S(n100) );
  ADDHXL U60 ( .A(n120), .B(n124), .CO(n101), .S(n102) );
  ADDFXL U61 ( .A(n123), .B(n121), .CI(n106), .CO(n103), .S(n104) );
  ADDHXL U62 ( .A(n125), .B(n122), .CO(n105), .S(n106) );
  ADDFXL U63 ( .A(n126), .B(a[4]), .CI(n124), .CO(n107), .S(n108) );
  ADDHXL U64 ( .A(n123), .B(n125), .CO(n109), .S(n110) );
  CLKINVX1 U88 ( .A(a[15]), .Y(n111) );
  CLKINVX1 U89 ( .A(a[8]), .Y(n118) );
  CLKINVX1 U90 ( .A(a[9]), .Y(n117) );
  CLKINVX1 U91 ( .A(a[10]), .Y(n116) );
  CLKINVX1 U92 ( .A(a[12]), .Y(n114) );
  CLKINVX1 U93 ( .A(a[11]), .Y(n115) );
  CLKINVX1 U94 ( .A(a[0]), .Y(n126) );
  CLKINVX1 U95 ( .A(a[4]), .Y(n122) );
  CLKBUFX3 U96 ( .A(a[15]), .Y(n127) );
  CLKINVX1 U97 ( .A(a[7]), .Y(n119) );
  CLKINVX1 U98 ( .A(a[3]), .Y(n123) );
  CLKINVX1 U99 ( .A(a[14]), .Y(n112) );
  CLKINVX1 U100 ( .A(a[2]), .Y(n124) );
  CLKINVX1 U101 ( .A(a[13]), .Y(n113) );
  CLKINVX1 U102 ( .A(a[6]), .Y(n120) );
  CLKINVX1 U103 ( .A(a[5]), .Y(n121) );
  CLKINVX1 U104 ( .A(a[1]), .Y(n125) );
endmodule


module FAS_DW_mult_tc_39 ( a, product );
  input [15:0] a;
  output [22:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73;

  CLKINVX1 U1 ( .A(n1), .Y(product[22]) );
  ADDFXL U2 ( .A(a[14]), .B(n59), .CI(n2), .CO(n1), .S(product[21]) );
  ADDFXL U3 ( .A(n60), .B(a[13]), .CI(n3), .CO(n2), .S(product[20]) );
  ADDFXL U4 ( .A(n61), .B(a[12]), .CI(n4), .CO(n3), .S(product[19]) );
  ADDFXL U5 ( .A(n29), .B(n62), .CI(n5), .CO(n4), .S(product[18]) );
  ADDFXL U6 ( .A(n30), .B(n31), .CI(n6), .CO(n5), .S(product[17]) );
  ADDFXL U7 ( .A(n32), .B(n33), .CI(n7), .CO(n6), .S(product[16]) );
  ADDFXL U8 ( .A(n35), .B(n34), .CI(n8), .CO(n7), .S(product[15]) );
  ADDFXL U9 ( .A(n36), .B(n37), .CI(n9), .CO(n8), .S(product[14]) );
  ADDFXL U10 ( .A(n38), .B(n39), .CI(n10), .CO(n9), .S(product[13]) );
  ADDFXL U11 ( .A(n40), .B(n41), .CI(n11), .CO(n10), .S(product[12]) );
  ADDFXL U12 ( .A(n42), .B(n43), .CI(n12), .CO(n11), .S(product[11]) );
  ADDFXL U13 ( .A(n44), .B(n45), .CI(n13), .CO(n12), .S(product[10]) );
  ADDFXL U14 ( .A(n46), .B(n47), .CI(n14), .CO(n13), .S(product[9]) );
  ADDFXL U15 ( .A(n48), .B(n49), .CI(n15), .CO(n14), .S(product[8]) );
  ADDFXL U16 ( .A(n50), .B(n51), .CI(n16), .CO(n15), .S(product[7]) );
  ADDFXL U17 ( .A(n52), .B(n53), .CI(n17), .CO(n16), .S(product[6]) );
  ADDFXL U18 ( .A(n54), .B(n55), .CI(n18), .CO(n17), .S(product[5]) );
  ADDFXL U19 ( .A(n56), .B(n57), .CI(n19), .CO(n18), .S(product[4]) );
  ADDFXL U20 ( .A(n58), .B(n72), .CI(n20), .CO(n19), .S(product[3]) );
  ADDFXL U21 ( .A(n22), .B(a[2]), .CI(n21), .CO(n20), .S(product[2]) );
  ADDHXL U22 ( .A(n73), .B(n22), .CO(n21), .S(product[1]) );
  CLKINVX1 U23 ( .A(n22), .Y(product[0]) );
  ADDFXL U27 ( .A(a[11]), .B(n60), .CI(a[15]), .CO(n29), .S(n30) );
  ADDFXL U28 ( .A(n61), .B(a[14]), .CI(a[10]), .CO(n31), .S(n32) );
  ADDFXL U29 ( .A(a[9]), .B(a[13]), .CI(a[15]), .CO(n33), .S(n34) );
  ADDFXL U30 ( .A(n62), .B(n60), .CI(a[8]), .CO(n35), .S(n36) );
  ADDFXL U31 ( .A(n63), .B(n61), .CI(a[7]), .CO(n37), .S(n38) );
  ADDFXL U32 ( .A(n64), .B(n62), .CI(a[6]), .CO(n39), .S(n40) );
  ADDFXL U33 ( .A(n65), .B(n63), .CI(a[5]), .CO(n41), .S(n42) );
  ADDFXL U34 ( .A(n66), .B(n64), .CI(a[4]), .CO(n43), .S(n44) );
  ADDFXL U35 ( .A(n67), .B(n65), .CI(a[3]), .CO(n45), .S(n46) );
  ADDFXL U36 ( .A(n68), .B(n66), .CI(a[2]), .CO(n47), .S(n48) );
  ADDFXL U37 ( .A(n69), .B(n67), .CI(a[1]), .CO(n49), .S(n50) );
  ADDFXL U38 ( .A(n70), .B(n68), .CI(a[0]), .CO(n51), .S(n52) );
  ADDHXL U39 ( .A(n69), .B(n71), .CO(n53), .S(n54) );
  ADDHXL U40 ( .A(n70), .B(n72), .CO(n55), .S(n56) );
  ADDHXL U41 ( .A(n71), .B(n73), .CO(n57), .S(n58) );
  CLKINVX1 U62 ( .A(a[15]), .Y(n59) );
  CLKINVX1 U63 ( .A(a[0]), .Y(n22) );
  CLKINVX1 U64 ( .A(a[12]), .Y(n62) );
  CLKINVX1 U65 ( .A(a[14]), .Y(n60) );
  CLKINVX1 U66 ( .A(a[1]), .Y(n73) );
  CLKINVX1 U67 ( .A(a[3]), .Y(n71) );
  CLKINVX1 U68 ( .A(a[13]), .Y(n61) );
  CLKINVX1 U69 ( .A(a[2]), .Y(n72) );
  CLKINVX1 U70 ( .A(a[4]), .Y(n70) );
  CLKINVX1 U71 ( .A(a[5]), .Y(n69) );
  CLKINVX1 U72 ( .A(a[6]), .Y(n68) );
  CLKINVX1 U73 ( .A(a[7]), .Y(n67) );
  CLKINVX1 U74 ( .A(a[8]), .Y(n66) );
  CLKINVX1 U75 ( .A(a[9]), .Y(n65) );
  CLKINVX1 U76 ( .A(a[10]), .Y(n64) );
  CLKINVX1 U77 ( .A(a[11]), .Y(n63) );
endmodule


module FAS_DW_mult_tc_40 ( a, product );
  input [15:0] a;
  output [30:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n29, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172;

  CLKINVX1 U1 ( .A(n1), .Y(product[30]) );
  ADDFXL U2 ( .A(n161), .B(n144), .CI(n2), .CO(n1), .S(product[29]) );
  ADDFXL U3 ( .A(n29), .B(n162), .CI(n3), .CO(n2), .S(product[28]) );
  ADDFXL U4 ( .A(n32), .B(n146), .CI(n4), .CO(n3), .S(product[27]) );
  ADDFXL U5 ( .A(n33), .B(n34), .CI(n5), .CO(n4), .S(product[26]) );
  ADDFXL U6 ( .A(n37), .B(n35), .CI(n6), .CO(n5), .S(product[25]) );
  ADDFXL U7 ( .A(n40), .B(n38), .CI(n7), .CO(n6), .S(product[24]) );
  ADDFXL U8 ( .A(n41), .B(n43), .CI(n8), .CO(n7), .S(product[23]) );
  ADDFXL U9 ( .A(n44), .B(n48), .CI(n9), .CO(n8), .S(product[22]) );
  ADDFXL U10 ( .A(n49), .B(n53), .CI(n10), .CO(n9), .S(product[21]) );
  ADDFXL U11 ( .A(n54), .B(n59), .CI(n11), .CO(n10), .S(product[20]) );
  ADDFXL U12 ( .A(n60), .B(n65), .CI(n12), .CO(n11), .S(product[19]) );
  ADDFXL U13 ( .A(n66), .B(n73), .CI(n13), .CO(n12), .S(product[18]) );
  ADDFXL U14 ( .A(n74), .B(n81), .CI(n14), .CO(n13), .S(product[17]) );
  ADDFXL U15 ( .A(n82), .B(n89), .CI(n15), .CO(n14), .S(product[16]) );
  ADDFXL U16 ( .A(n90), .B(n97), .CI(n16), .CO(n15), .S(product[15]) );
  ADDFXL U17 ( .A(n98), .B(n105), .CI(n17), .CO(n16), .S(product[14]) );
  ADDFXL U18 ( .A(n106), .B(n111), .CI(n18), .CO(n17), .S(product[13]) );
  ADDFXL U19 ( .A(n112), .B(n117), .CI(n19), .CO(n18), .S(product[12]) );
  ADDFXL U20 ( .A(n118), .B(n124), .CI(n20), .CO(n19), .S(product[11]) );
  ADDFXL U21 ( .A(n125), .B(n129), .CI(n21), .CO(n20), .S(product[10]) );
  ADDFXL U22 ( .A(n130), .B(n134), .CI(n22), .CO(n21), .S(product[9]) );
  ADDFXL U23 ( .A(n135), .B(n136), .CI(n23), .CO(n22), .S(product[8]) );
  ADDFXL U24 ( .A(n137), .B(n140), .CI(n24), .CO(n23), .S(product[7]) );
  ADDFXL U25 ( .A(n141), .B(n142), .CI(n25), .CO(n24), .S(product[6]) );
  ADDFXL U26 ( .A(n143), .B(product[0]), .CI(n26), .CO(n25), .S(product[5]) );
  ADDFXL U27 ( .A(n171), .B(product[1]), .CI(n27), .CO(n26), .S(product[4]) );
  ADDHXL U28 ( .A(product[0]), .B(n172), .CO(n27), .S(product[3]) );
  CLKINVX1 U29 ( .A(n161), .Y(n29) );
  ADDFXL U33 ( .A(n163), .B(n29), .CI(a[15]), .CO(n32), .S(n33) );
  ADDFXL U34 ( .A(n164), .B(a[14]), .CI(n36), .CO(n34), .S(n35) );
  CMPR42X1 U35 ( .A(n144), .B(n147), .C(n146), .D(n165), .ICI(n39), .S(n38), 
        .ICO(n36), .CO(n37) );
  CMPR42X1 U36 ( .A(a[12]), .B(n161), .C(n166), .D(n45), .ICI(n42), .S(n41), 
        .ICO(n39), .CO(n40) );
  CMPR42X1 U37 ( .A(n144), .B(n148), .C(n50), .D(n46), .ICI(n47), .S(n44), 
        .ICO(n42), .CO(n43) );
  ADDFXL U38 ( .A(n162), .B(n149), .CI(n167), .CO(n45), .S(n46) );
  CMPR42X1 U39 ( .A(n163), .B(n55), .C(n51), .D(n56), .ICI(n52), .S(n49), 
        .ICO(n47), .CO(n48) );
  ADDFXL U40 ( .A(n161), .B(a[10]), .CI(n168), .CO(n50), .S(n51) );
  CMPR42X1 U41 ( .A(n144), .B(n150), .C(n62), .D(n57), .ICI(n58), .S(n54), 
        .ICO(n52), .CO(n53) );
  CMPR42X1 U42 ( .A(n151), .B(n169), .C(n164), .D(n162), .ICI(n61), .S(n57), 
        .ICO(n55), .CO(n56) );
  CMPR42X1 U43 ( .A(n170), .B(n70), .C(n68), .D(n63), .ICI(n64), .S(n60), 
        .ICO(n58), .CO(n59) );
  CMPR42X1 U44 ( .A(a[8]), .B(n165), .C(n161), .D(n163), .ICI(n67), .S(n63), 
        .ICO(n61), .CO(n62) );
  CMPR42X1 U45 ( .A(n78), .B(n71), .C(n76), .D(n69), .ICI(n72), .S(n66), .ICO(
        n64), .CO(n65) );
  CMPR42X1 U46 ( .A(n144), .B(n152), .C(n162), .D(n164), .ICI(n75), .S(n69), 
        .ICO(n67), .CO(n68) );
  ADDFXL U47 ( .A(n171), .B(n153), .CI(n166), .CO(n70), .S(n71) );
  CMPR42X1 U48 ( .A(n79), .B(n86), .C(n84), .D(n77), .ICI(n80), .S(n74), .ICO(
        n72), .CO(n73) );
  CMPR42X1 U49 ( .A(n154), .B(n165), .C(n167), .D(n172), .ICI(n83), .S(n77), 
        .ICO(n75), .CO(n76) );
  ADDFXL U50 ( .A(n163), .B(a[6]), .CI(n161), .CO(n78), .S(n79) );
  CMPR42X1 U51 ( .A(n87), .B(n94), .C(n92), .D(n85), .ICI(n88), .S(n82), .ICO(
        n80), .CO(n81) );
  CMPR42X1 U52 ( .A(n144), .B(n166), .C(n168), .D(product[2]), .ICI(n91), .S(
        n85), .ICO(n83), .CO(n84) );
  ADDFXL U53 ( .A(n164), .B(a[5]), .CI(n162), .CO(n86), .S(n87) );
  CMPR42X1 U54 ( .A(n165), .B(n95), .C(n93), .D(n100), .ICI(n96), .S(n90), 
        .ICO(n88), .CO(n89) );
  CMPR42X1 U55 ( .A(n155), .B(n169), .C(n163), .D(n102), .ICI(n99), .S(n93), 
        .ICO(n91), .CO(n92) );
  ADDFXL U56 ( .A(product[1]), .B(a[15]), .CI(n167), .CO(n94), .S(n95) );
  CMPR42X1 U57 ( .A(n168), .B(product[0]), .C(n108), .D(n101), .ICI(n104), .S(
        n98), .ICO(n96), .CO(n97) );
  CMPR42X1 U58 ( .A(n166), .B(n161), .C(n164), .D(n103), .ICI(n107), .S(n101), 
        .ICO(n99), .CO(n100) );
  ADDHXL U59 ( .A(n156), .B(n170), .CO(n102), .S(n103) );
  CMPR42X1 U60 ( .A(n165), .B(n167), .C(n114), .D(n109), .ICI(n110), .S(n106), 
        .ICO(n104), .CO(n105) );
  CMPR42X1 U61 ( .A(n157), .B(n171), .C(n169), .D(n162), .ICI(n113), .S(n109), 
        .ICO(n107), .CO(n108) );
  CMPR42X1 U62 ( .A(n163), .B(n166), .C(n116), .D(n119), .ICI(n115), .S(n112), 
        .ICO(n110), .CO(n111) );
  CMPR42X1 U63 ( .A(n158), .B(n172), .C(n170), .D(n168), .ICI(n121), .S(n115), 
        .ICO(n113), .CO(n114) );
  CMPR42X1 U64 ( .A(n164), .B(n167), .C(n123), .D(n126), .ICI(n120), .S(n118), 
        .ICO(n116), .CO(n117) );
  ADDFXL U65 ( .A(product[2]), .B(n169), .CI(n122), .CO(n119), .S(n120) );
  XNOR2X1 U66 ( .A(n171), .B(n159), .Y(n122) );
  OR2X1 U67 ( .A(n171), .B(n159), .Y(n121) );
  CMPR42X1 U68 ( .A(n165), .B(n170), .C(n168), .D(n128), .ICI(n127), .S(n125), 
        .ICO(n123), .CO(n124) );
  ADDFXL U69 ( .A(product[1]), .B(n172), .CI(n138), .CO(n126), .S(n127) );
  CMPR42X1 U70 ( .A(n166), .B(n171), .C(n169), .D(n139), .ICI(n133), .S(n130), 
        .ICO(n128), .CO(n129) );
  CMPR42X1 U72 ( .A(n172), .B(product[1]), .C(n170), .D(n167), .ICI(n138), .S(
        n135), .ICO(n133), .CO(n134) );
  ADDFXL U73 ( .A(n171), .B(n168), .CI(n139), .CO(n136), .S(n137) );
  ADDHXL U74 ( .A(product[2]), .B(product[0]), .CO(n138), .S(n139) );
  ADDFXL U75 ( .A(product[1]), .B(n169), .CI(n172), .CO(n140), .S(n141) );
  ADDHXL U76 ( .A(n170), .B(product[2]), .CO(n142), .S(n143) );
  CLKINVX1 U112 ( .A(a[6]), .Y(n153) );
  CLKINVX1 U113 ( .A(a[10]), .Y(n149) );
  CLKINVX1 U114 ( .A(a[3]), .Y(n156) );
  CLKBUFX3 U115 ( .A(a[0]), .Y(product[0]) );
  CLKINVX1 U116 ( .A(a[4]), .Y(n155) );
  CLKINVX1 U117 ( .A(a[2]), .Y(n157) );
  CLKINVX1 U118 ( .A(a[5]), .Y(n154) );
  CLKINVX1 U119 ( .A(a[8]), .Y(n151) );
  CLKINVX1 U120 ( .A(a[7]), .Y(n152) );
  CLKINVX1 U121 ( .A(a[1]), .Y(n158) );
  CLKBUFX3 U122 ( .A(a[1]), .Y(product[1]) );
  CLKBUFX3 U123 ( .A(a[10]), .Y(n165) );
  CLKBUFX3 U124 ( .A(a[9]), .Y(n166) );
  CLKBUFX3 U125 ( .A(a[2]), .Y(product[2]) );
  CLKINVX1 U126 ( .A(a[13]), .Y(n146) );
  CLKINVX1 U127 ( .A(a[12]), .Y(n147) );
  CLKINVX1 U128 ( .A(a[15]), .Y(n144) );
  CLKBUFX3 U129 ( .A(a[14]), .Y(n161) );
  CLKINVX1 U130 ( .A(a[11]), .Y(n148) );
  CLKINVX1 U131 ( .A(a[9]), .Y(n150) );
  CLKBUFX3 U132 ( .A(a[5]), .Y(n170) );
  CLKBUFX3 U133 ( .A(a[8]), .Y(n167) );
  CLKBUFX3 U134 ( .A(a[6]), .Y(n169) );
  CLKBUFX3 U135 ( .A(a[13]), .Y(n162) );
  CLKBUFX3 U136 ( .A(a[7]), .Y(n168) );
  CLKBUFX3 U137 ( .A(a[12]), .Y(n163) );
  CLKBUFX3 U138 ( .A(a[3]), .Y(n172) );
  CLKBUFX3 U139 ( .A(a[11]), .Y(n164) );
  CLKBUFX3 U140 ( .A(a[4]), .Y(n171) );
  CLKINVX1 U141 ( .A(a[0]), .Y(n159) );
endmodule


module FAS_DW_mult_tc_41 ( a, product_28_, product_27_, product_26_, 
        product_25_, product_24_, product_23_, product_22_, product_21_, 
        product_20_, product_19_, product_18_, product_17_, product_16_, 
        product_15_, product_14_, product_13_, product_12_, product_11_, 
        product_10_, product_9_, product_8_, product_7_, product_6_, 
        product_5_, product_4_, product_3_, product_2_, product_1_ );
  input [15:0] a;
  output product_28_, product_27_, product_26_, product_25_, product_24_,
         product_23_, product_22_, product_21_, product_20_, product_19_,
         product_18_, product_17_, product_16_, product_15_, product_14_,
         product_13_, product_12_, product_11_, product_10_, product_9_,
         product_8_, product_7_, product_6_, product_5_, product_4_,
         product_3_, product_2_, product_1_;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122;

  CLKINVX1 U2 ( .A(n109), .Y(product_27_) );
  ADDFXL U4 ( .A(n110), .B(a[15]), .CI(n3), .CO(product_26_), .S(product_25_)
         );
  ADDFXL U5 ( .A(n25), .B(n111), .CI(n4), .CO(n3), .S(product_24_) );
  ADDFXL U6 ( .A(n28), .B(n26), .CI(n5), .CO(n4), .S(product_23_) );
  ADDFXL U7 ( .A(n29), .B(n31), .CI(n6), .CO(n5), .S(product_22_) );
  ADDFXL U8 ( .A(n32), .B(n34), .CI(n7), .CO(n6), .S(product_21_) );
  ADDFXL U9 ( .A(n37), .B(n35), .CI(n8), .CO(n7), .S(product_20_) );
  ADDFXL U10 ( .A(n40), .B(n38), .CI(n9), .CO(n8), .S(product_19_) );
  ADDFXL U11 ( .A(n41), .B(n45), .CI(n10), .CO(n9), .S(product_18_) );
  ADDFXL U12 ( .A(n46), .B(n51), .CI(n11), .CO(n10), .S(product_17_) );
  ADDFXL U13 ( .A(n52), .B(n57), .CI(n12), .CO(n11), .S(product_16_) );
  ADDFXL U14 ( .A(n58), .B(n63), .CI(n13), .CO(n12), .S(product_15_) );
  ADDFXL U15 ( .A(n64), .B(n69), .CI(n14), .CO(n13), .S(product_14_) );
  ADDFXL U16 ( .A(n70), .B(n75), .CI(n15), .CO(n14), .S(product_13_) );
  ADDFXL U17 ( .A(n76), .B(n81), .CI(n16), .CO(n15), .S(product_12_) );
  ADDFXL U18 ( .A(n82), .B(n88), .CI(n17), .CO(n16), .S(product_11_) );
  ADDFXL U19 ( .A(n89), .B(n93), .CI(n18), .CO(n17), .S(product_10_) );
  ADDFXL U20 ( .A(n94), .B(n97), .CI(n19), .CO(n18), .S(product_9_) );
  ADDFXL U21 ( .A(n98), .B(n101), .CI(n20), .CO(n19), .S(product_8_) );
  ADDFXL U22 ( .A(n102), .B(n103), .CI(n21), .CO(n20), .S(product_7_) );
  ADDFXL U23 ( .A(n104), .B(n105), .CI(n22), .CO(n21), .S(product_6_) );
  ADDFXL U24 ( .A(n106), .B(n107), .CI(n23), .CO(n22), .S(product_5_) );
  ADDFXL U25 ( .A(n85), .B(product_1_), .CI(n108), .CO(n23), .S(product_4_) );
  ADDFXL U27 ( .A(n112), .B(n110), .CI(n27), .CO(n25), .S(n26) );
  CMPR42X1 U28 ( .A(a[15]), .B(n110), .C(n113), .D(n111), .ICI(n30), .S(n29), 
        .ICO(n27), .CO(n28) );
  CMPR42X1 U29 ( .A(a[15]), .B(n111), .C(n114), .D(n112), .ICI(n33), .S(n32), 
        .ICO(n30), .CO(n31) );
  CMPR42X1 U30 ( .A(a[15]), .B(n112), .C(n115), .D(n113), .ICI(n36), .S(n35), 
        .ICO(n33), .CO(n34) );
  CMPR42X1 U31 ( .A(n113), .B(n116), .C(n114), .D(n42), .ICI(n39), .S(n38), 
        .ICO(n36), .CO(n37) );
  CMPR42X1 U32 ( .A(n115), .B(n47), .C(n43), .D(n48), .ICI(n44), .S(n41), 
        .ICO(n39), .CO(n40) );
  ADDFXL U33 ( .A(n114), .B(n110), .CI(n117), .CO(n42), .S(n43) );
  CMPR42X1 U34 ( .A(n111), .B(n115), .C(n54), .D(n49), .ICI(n50), .S(n46), 
        .ICO(n44), .CO(n45) );
  CMPR42X1 U35 ( .A(a[15]), .B(n116), .C(n118), .D(n110), .ICI(n53), .S(n49), 
        .ICO(n47), .CO(n48) );
  CMPR42X1 U36 ( .A(n112), .B(n116), .C(n55), .D(n60), .ICI(n56), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U37 ( .A(a[15]), .B(n117), .C(n119), .D(n111), .ICI(n59), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U38 ( .A(n112), .B(n113), .C(n66), .D(n61), .ICI(n62), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U39 ( .A(n118), .B(n120), .C(n117), .D(n110), .ICI(n65), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U40 ( .A(n113), .B(n114), .C(n72), .D(n67), .ICI(n68), .S(n64), 
        .ICO(n62), .CO(n63) );
  CMPR42X1 U41 ( .A(n119), .B(n121), .C(n118), .D(n111), .ICI(n71), .S(n67), 
        .ICO(n65), .CO(n66) );
  CMPR42X1 U42 ( .A(n114), .B(n115), .C(n78), .D(n74), .ICI(n73), .S(n70), 
        .ICO(n68), .CO(n69) );
  CMPR42X1 U43 ( .A(n120), .B(n122), .C(n119), .D(n112), .ICI(n77), .S(n73), 
        .ICO(n71), .CO(n72) );
  CMPR42X1 U44 ( .A(n113), .B(n115), .C(n80), .D(n83), .ICI(n79), .S(n76), 
        .ICO(n74), .CO(n75) );
  CMPR42X1 U45 ( .A(n121), .B(product_2_), .C(n120), .D(n116), .ICI(n85), .S(
        n79), .ICO(n77), .CO(n78) );
  CMPR42X1 U46 ( .A(n114), .B(product_3_), .C(n87), .D(n90), .ICI(n84), .S(n82), .ICO(n80), .CO(n81) );
  ADDFXL U47 ( .A(n121), .B(n117), .CI(n116), .CO(n83), .S(n84) );
  ADDHXL U48 ( .A(n122), .B(product_1_), .CO(n85), .S(product_3_) );
  CMPR42X1 U49 ( .A(n115), .B(n118), .C(n117), .D(n92), .ICI(n91), .S(n89), 
        .ICO(n87), .CO(n88) );
  ADDFXL U50 ( .A(product_2_), .B(n122), .CI(n95), .CO(n90), .S(n91) );
  CMPR42X1 U51 ( .A(n116), .B(n119), .C(n118), .D(n99), .ICI(n96), .S(n94), 
        .ICO(n92), .CO(n93) );
  ADDHXL U52 ( .A(product_2_), .B(product_1_), .CO(n95), .S(n96) );
  ADDFXL U53 ( .A(n119), .B(n117), .CI(n100), .CO(n97), .S(n98) );
  ADDHXL U54 ( .A(n120), .B(product_1_), .CO(n99), .S(n100) );
  ADDFXL U55 ( .A(n121), .B(n118), .CI(n120), .CO(n101), .S(n102) );
  ADDFXL U56 ( .A(n122), .B(n119), .CI(n121), .CO(n103), .S(n104) );
  ADDFXL U57 ( .A(product_2_), .B(n120), .CI(n122), .CO(n105), .S(n106) );
  ADDHXL U58 ( .A(n121), .B(product_2_), .CO(n107), .S(n108) );
  CLKBUFX3 U79 ( .A(product_27_), .Y(product_28_) );
  CLKINVX1 U80 ( .A(a[15]), .Y(n109) );
  CLKBUFX3 U81 ( .A(a[0]), .Y(product_1_) );
  CLKBUFX3 U82 ( .A(a[1]), .Y(product_2_) );
  CLKBUFX3 U83 ( .A(a[9]), .Y(n115) );
  CLKBUFX3 U84 ( .A(a[11]), .Y(n113) );
  CLKBUFX3 U85 ( .A(a[8]), .Y(n116) );
  CLKBUFX3 U86 ( .A(a[10]), .Y(n114) );
  CLKBUFX3 U87 ( .A(a[6]), .Y(n118) );
  CLKBUFX3 U88 ( .A(a[12]), .Y(n112) );
  CLKBUFX3 U89 ( .A(a[5]), .Y(n119) );
  CLKBUFX3 U90 ( .A(a[13]), .Y(n111) );
  CLKBUFX3 U91 ( .A(a[4]), .Y(n120) );
  CLKBUFX3 U92 ( .A(a[7]), .Y(n117) );
  CLKBUFX3 U93 ( .A(a[3]), .Y(n121) );
  CLKBUFX3 U94 ( .A(a[14]), .Y(n110) );
  CLKBUFX3 U95 ( .A(a[2]), .Y(n122) );
endmodule


module FAS_DW_mult_tc_42 ( a, product_28_, product_27_, product_26_, 
        product_25_, product_24_, product_23_, product_22_, product_21_, 
        product_20_, product_19_, product_18_, product_17_, product_16_, 
        product_15_, product_14_, product_13_, product_12_, product_11_, 
        product_10_, product_9_, product_8_, product_7_, product_6_, 
        product_5_, product_4_, product_3_, product_2_, product_1_ );
  input [15:0] a;
  output product_28_, product_27_, product_26_, product_25_, product_24_,
         product_23_, product_22_, product_21_, product_20_, product_19_,
         product_18_, product_17_, product_16_, product_15_, product_14_,
         product_13_, product_12_, product_11_, product_10_, product_9_,
         product_8_, product_7_, product_6_, product_5_, product_4_,
         product_3_, product_2_, product_1_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84, n85, n87;

  CLKINVX1 U3 ( .A(n2), .Y(product_27_) );
  ADDFXL U4 ( .A(a[15]), .B(n68), .CI(n3), .CO(n2), .S(product_26_) );
  ADDFXL U5 ( .A(n69), .B(a[14]), .CI(n4), .CO(n3), .S(product_25_) );
  ADDFXL U6 ( .A(n70), .B(a[13]), .CI(n5), .CO(n4), .S(product_24_) );
  ADDFXL U7 ( .A(n71), .B(a[12]), .CI(n6), .CO(n5), .S(product_23_) );
  ADDFXL U8 ( .A(n26), .B(a[11]), .CI(n7), .CO(n6), .S(product_22_) );
  ADDFXL U9 ( .A(n27), .B(n28), .CI(n8), .CO(n7), .S(product_21_) );
  ADDFXL U10 ( .A(n30), .B(n29), .CI(n9), .CO(n8), .S(product_20_) );
  ADDFXL U11 ( .A(n33), .B(n31), .CI(n10), .CO(n9), .S(product_19_) );
  ADDFXL U12 ( .A(n34), .B(n36), .CI(n11), .CO(n10), .S(product_18_) );
  ADDFXL U13 ( .A(n37), .B(n39), .CI(n12), .CO(n11), .S(product_17_) );
  ADDFXL U14 ( .A(n40), .B(n42), .CI(n13), .CO(n12), .S(product_16_) );
  ADDFXL U15 ( .A(n43), .B(n45), .CI(n14), .CO(n13), .S(product_15_) );
  ADDFXL U16 ( .A(n46), .B(n48), .CI(n15), .CO(n14), .S(product_14_) );
  ADDFXL U17 ( .A(n49), .B(n51), .CI(n16), .CO(n15), .S(product_13_) );
  ADDFXL U18 ( .A(n52), .B(n53), .CI(n17), .CO(n16), .S(product_12_) );
  ADDFXL U19 ( .A(n54), .B(n57), .CI(n18), .CO(n17), .S(product_11_) );
  ADDFXL U20 ( .A(n58), .B(n59), .CI(n19), .CO(n18), .S(product_10_) );
  ADDFXL U21 ( .A(n60), .B(n61), .CI(n20), .CO(n19), .S(product_9_) );
  ADDFXL U22 ( .A(n62), .B(n63), .CI(n21), .CO(n20), .S(product_8_) );
  ADDFXL U23 ( .A(n64), .B(n65), .CI(n22), .CO(n21), .S(product_7_) );
  ADDFXL U24 ( .A(n66), .B(a[3]), .CI(n23), .CO(n22), .S(product_6_) );
  ADDFXL U25 ( .A(a[4]), .B(a[2]), .CI(n24), .CO(n23), .S(product_5_) );
  ADDFXL U26 ( .A(a[3]), .B(a[1]), .CI(n25), .CO(n24), .S(product_4_) );
  ADDHXL U27 ( .A(a[0]), .B(a[2]), .CO(n25), .S(product_3_) );
  ADDFXL U28 ( .A(n72), .B(n68), .CI(a[15]), .CO(n26), .S(n27) );
  ADDFXL U29 ( .A(n69), .B(a[14]), .CI(n73), .CO(n28), .S(n29) );
  ADDFXL U30 ( .A(n74), .B(a[13]), .CI(n32), .CO(n30), .S(n31) );
  CMPR42X1 U31 ( .A(n75), .B(n71), .C(n70), .D(n67), .ICI(n35), .S(n34), .ICO(
        n32), .CO(n33) );
  CMPR42X1 U32 ( .A(a[11]), .B(n76), .C(n67), .D(n84), .ICI(n38), .S(n37), 
        .ICO(n35), .CO(n36) );
  CMPR42X1 U33 ( .A(a[15]), .B(n72), .C(n77), .D(n85), .ICI(n41), .S(n40), 
        .ICO(n38), .CO(n39) );
  CMPR42X1 U34 ( .A(n78), .B(n73), .C(a[12]), .D(n84), .ICI(n44), .S(n43), 
        .ICO(n41), .CO(n42) );
  CMPR42X1 U35 ( .A(n79), .B(n74), .C(n87), .D(n85), .ICI(n47), .S(n46), .ICO(
        n44), .CO(n45) );
  CMPR42X1 U36 ( .A(n80), .B(n75), .C(a[10]), .D(a[12]), .ICI(n50), .S(n49), 
        .ICO(n47), .CO(n48) );
  CMPR42X1 U37 ( .A(n81), .B(n76), .C(a[9]), .D(n87), .ICI(n55), .S(n52), 
        .ICO(n50), .CO(n51) );
  ADDFXL U38 ( .A(a[8]), .B(a[10]), .CI(n56), .CO(n53), .S(n54) );
  XNOR2X1 U39 ( .A(n77), .B(n82), .Y(n56) );
  OR2X1 U40 ( .A(n77), .B(n82), .Y(n55) );
  ADDFXL U41 ( .A(a[7]), .B(n78), .CI(a[9]), .CO(n57), .S(n58) );
  ADDFXL U42 ( .A(a[6]), .B(n79), .CI(a[8]), .CO(n59), .S(n60) );
  ADDFXL U43 ( .A(a[5]), .B(n80), .CI(a[7]), .CO(n61), .S(n62) );
  ADDFXL U44 ( .A(a[4]), .B(n81), .CI(a[6]), .CO(n63), .S(n64) );
  XNOR2X1 U45 ( .A(a[5]), .B(n82), .Y(n66) );
  OR2X1 U46 ( .A(a[5]), .B(n82), .Y(n65) );
  CLKBUFX3 U70 ( .A(product_27_), .Y(product_28_) );
  CLKBUFX3 U71 ( .A(a[11]), .Y(n87) );
  CLKBUFX3 U72 ( .A(a[13]), .Y(n85) );
  CLKBUFX3 U73 ( .A(a[14]), .Y(n84) );
  CLKINVX1 U74 ( .A(a[6]), .Y(n76) );
  CLKINVX1 U75 ( .A(a[7]), .Y(n75) );
  CLKINVX1 U76 ( .A(a[9]), .Y(n73) );
  CLKINVX1 U77 ( .A(a[5]), .Y(n77) );
  CLKINVX1 U78 ( .A(a[15]), .Y(n67) );
  CLKINVX1 U79 ( .A(a[8]), .Y(n74) );
  CLKINVX1 U80 ( .A(a[10]), .Y(n72) );
  CLKINVX1 U81 ( .A(a[11]), .Y(n71) );
  CLKINVX1 U82 ( .A(a[0]), .Y(n82) );
  CLKINVX1 U83 ( .A(a[1]), .Y(n81) );
  CLKINVX1 U84 ( .A(a[2]), .Y(n80) );
  CLKINVX1 U85 ( .A(a[3]), .Y(n79) );
  CLKINVX1 U86 ( .A(a[4]), .Y(n78) );
  CLKINVX1 U87 ( .A(a[12]), .Y(n70) );
  CLKINVX1 U88 ( .A(a[14]), .Y(n68) );
  CLKINVX1 U89 ( .A(a[13]), .Y(n69) );
  BUFX2 U90 ( .A(a[0]), .Y(product_1_) );
  BUFX2 U91 ( .A(a[1]), .Y(product_2_) );
endmodule


module FAS ( data_valid, data, clk, rst, fir_d, fir_valid, fft_valid, done, 
        freq, fft_d1, fft_d2, fft_d3, fft_d4, fft_d5, fft_d6, fft_d7, fft_d8, 
        fft_d9, fft_d10, fft_d11, fft_d12, fft_d13, fft_d14, fft_d15, fft_d0, 
        test_si, test_se );
  input [15:0] data;
  output [15:0] fir_d;
  output [3:0] freq;
  output [31:0] fft_d1;
  output [31:0] fft_d2;
  output [31:0] fft_d3;
  output [31:0] fft_d4;
  output [31:0] fft_d5;
  output [31:0] fft_d6;
  output [31:0] fft_d7;
  output [31:0] fft_d8;
  output [31:0] fft_d9;
  output [31:0] fft_d10;
  output [31:0] fft_d11;
  output [31:0] fft_d12;
  output [31:0] fft_d13;
  output [31:0] fft_d14;
  output [31:0] fft_d15;
  output [31:0] fft_d0;
  input data_valid, clk, rst, test_si, test_se;
  output fir_valid, fft_valid, done;
  wire   hd01_35, hd02_35, hd03_35, hd04_35, hd05_35, hd06_35, hd07_35,
         hd08_35, hd08_20_, hd08_19_, hd08_18_, hd08_17_, hd08_16_, hd08_15_,
         hd08_14_, hd08_13_, hd08_12_, hd08_11_, hd08_10_, hd08_9_, hd08_8_,
         hd08_7_, hd08_6_, hd08_5_, hd09_35, hd10_35, hd11_35, hd12_35,
         hd13_35, hd14_35, hd15_35, hd16_35, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, multiplier_r_31, multiplier_r_8, multiplier_r_6, N162, N163,
         N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174,
         N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185,
         N186, N187, N188, N189, N190, N191, N192, N193, multiplier_i_31,
         multiplier_i_9, multiplier_i_8, multiplier_i_6, multiplier_i_0, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, BF2I_b_s, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N359, N360, N361, N362, N363, N368, N369, N370, N371, N372,
         N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
         N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394,
         N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
         N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416,
         N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427,
         N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N569, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582,
         N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593,
         N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604,
         N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615,
         N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626,
         N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648,
         N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659,
         N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670,
         N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681,
         N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692,
         N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703,
         N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714,
         N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725,
         N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736,
         N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747,
         N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758,
         N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769,
         N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813,
         N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824,
         N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835,
         N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846,
         N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857,
         N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868,
         N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879,
         N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890,
         N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901,
         N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912,
         N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923,
         N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934,
         N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945,
         N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956,
         N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967,
         N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978,
         N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989,
         N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000,
         N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010,
         N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020,
         N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030,
         N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040,
         N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050,
         N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060,
         N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070,
         N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080,
         N1081, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091,
         N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101,
         N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111,
         N1112, N1113, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122,
         N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132,
         N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142,
         N1143, N1144, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196,
         N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206,
         N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216,
         N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1230, N1231,
         N1232, N1233, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354,
         N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364,
         N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374,
         N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384,
         N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394,
         N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403, N1404,
         N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413, N1414,
         N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423, N1424,
         N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433, N1434,
         N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443, N1444,
         N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453, N1454,
         N1455, N1456, N1457, N1458, U3_U3_Z_0, U3_U3_Z_1, U3_U3_Z_2,
         U3_U3_Z_3, U3_U3_Z_4, U3_U3_Z_5, U3_U3_Z_6, U3_U3_Z_7, U3_U3_Z_8,
         U3_U3_Z_9, U3_U3_Z_10, U3_U3_Z_11, U3_U3_Z_12, U3_U3_Z_13, U3_U3_Z_14,
         U3_U3_Z_15, U3_U5_Z_0, U3_U5_Z_1, U3_U5_Z_2, U3_U5_Z_3, U3_U5_Z_4,
         U3_U5_Z_5, U3_U5_Z_6, U3_U5_Z_7, U3_U5_Z_8, U3_U5_Z_9, U3_U5_Z_10,
         U3_U5_Z_11, U3_U5_Z_12, U3_U5_Z_13, U3_U5_Z_14, U3_U5_Z_15,
         U3_U5_Z_16, U3_U5_Z_17, U3_U5_Z_18, U3_U5_Z_19, U3_U5_Z_20,
         U3_U5_Z_21, U3_U5_Z_22, U3_U5_Z_23, U3_U5_Z_24, U3_U5_Z_25,
         U3_U5_Z_26, U3_U5_Z_27, U3_U5_Z_28, U3_U5_Z_29, U3_U5_Z_30,
         U3_U5_Z_31, U3_U6_Z_0, U3_U6_Z_1, U3_U6_Z_2, U3_U6_Z_3, U3_U6_Z_4,
         U3_U6_Z_5, U3_U6_Z_6, U3_U6_Z_7, U3_U6_Z_8, U3_U6_Z_9, U3_U6_Z_10,
         U3_U6_Z_11, U3_U6_Z_12, U3_U6_Z_13, U3_U6_Z_14, U3_U6_Z_15,
         U3_U6_Z_16, U3_U6_Z_17, U3_U6_Z_18, U3_U6_Z_19, U3_U6_Z_20,
         U3_U6_Z_21, U3_U6_Z_22, U3_U6_Z_23, U3_U6_Z_24, U3_U6_Z_25,
         U3_U6_Z_26, U3_U6_Z_27, U3_U6_Z_28, U3_U6_Z_29, U3_U6_Z_30,
         U3_U6_Z_31, U3_U7_Z_0, U3_U7_Z_1, U3_U7_Z_2, U3_U7_Z_3, U3_U7_Z_4,
         U3_U7_Z_5, U3_U7_Z_6, U3_U7_Z_7, U3_U7_Z_8, U3_U7_Z_9, U3_U7_Z_10,
         U3_U7_Z_11, U3_U7_Z_12, U3_U7_Z_13, U3_U7_Z_14, U3_U7_Z_15,
         U3_U7_Z_16, U3_U7_Z_17, U3_U7_Z_18, U3_U7_Z_19, U3_U7_Z_20,
         U3_U7_Z_21, U3_U7_Z_22, U3_U7_Z_23, U3_U7_Z_24, U3_U7_Z_25,
         U3_U7_Z_26, U3_U7_Z_27, U3_U7_Z_28, U3_U7_Z_29, U3_U7_Z_30,
         U3_U7_Z_31, U3_U8_Z_0, U3_U8_Z_1, U3_U8_Z_2, U3_U8_Z_3, U3_U8_Z_4,
         U3_U8_Z_5, U3_U8_Z_6, U3_U8_Z_7, U3_U8_Z_8, U3_U8_Z_9, U3_U8_Z_10,
         U3_U8_Z_11, U3_U8_Z_12, U3_U8_Z_13, U3_U8_Z_14, U3_U8_Z_15,
         U3_U8_Z_16, U3_U8_Z_17, U3_U8_Z_18, U3_U8_Z_19, U3_U8_Z_20,
         U3_U8_Z_21, U3_U8_Z_22, U3_U8_Z_23, U3_U8_Z_24, U3_U8_Z_25,
         U3_U8_Z_26, U3_U8_Z_27, U3_U8_Z_28, U3_U8_Z_29, U3_U8_Z_30,
         U3_U8_Z_31, n2850, n2860, n2870, n2880, n2890, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n3000, n3010, n3020, n3030, n3040,
         n3050, n3060, n30700, n3080, n3090, n3100, n3110, n3120, n3130, n3140,
         n3150, n3160, n1599, n1601, n1603, n1605, n1607, n1609, n1611, n1613,
         n1615, n1617, n1619, n1621, n1623, n1625, n1627, n1629, n1631, n1633,
         n1635, n1637, n1639, n1641, n1643, n1645, n1647, n1649, n1651, n1653,
         n1655, n1657, n1659, n1661, n1663, n1665, n1667, n1669, n1671, n1673,
         n1675, n1677, n1679, n1681, n1683, n1685, n1687, n1689, n1691, n1693,
         n1695, n1697, n1699, n1701, n1703, n1705, n1707, n1709, n1711, n1713,
         n1715, n1717, n1719, n1721, n1723, n1725, n1824, n1832, n1840, n1848,
         n1856, n1864, n1872, n1880, n1888, n1896, n1904, n1912, n1920, n1928,
         n1936, n1944, n3067, n3068, n3069, n30701, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3461, n3462, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n40101, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6064, n6067, n6068, n6071, n6072, n6073, n6074,
         n6075, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         mult_add_355_aco_b, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n101101, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224;
  wire   [22:0] hd01;
  wire   [22:0] hd02;
  wire   [22:0] hd03;
  wire   [21:0] hd04;
  wire   [24:0] hd05;
  wire   [25:0] hd06;
  wire   [25:0] hd07;
  wire   [26:0] hd09;
  wire   [27:0] hd10;
  wire   [27:0] hd11;
  wire   [25:0] hd12;
  wire   [27:0] hd13;
  wire   [28:0] hd14;
  wire   [29:0] hd15;
  wire   [29:0] hd16;
  wire   [35:0] d01;
  wire   [35:1] hd_a02;
  wire   [35:0] d02;
  wire   [35:0] hd_a03;
  wire   [35:0] d03;
  wire   [35:0] hd_a04;
  wire   [35:0] d04;
  wire   [35:0] hd_a05;
  wire   [35:0] d05;
  wire   [35:0] hd_a06;
  wire   [35:0] d06;
  wire   [35:0] hd_a07;
  wire   [35:0] d07;
  wire   [35:0] hd_a08;
  wire   [35:0] d08;
  wire   [35:0] hd_a09;
  wire   [35:0] d09;
  wire   [35:0] hd_a10;
  wire   [35:0] d10;
  wire   [35:0] hd_a11;
  wire   [35:0] d11;
  wire   [35:0] hd_a12;
  wire   [35:0] d12;
  wire   [35:0] hd_a13;
  wire   [35:0] d13;
  wire   [35:0] hd_a14;
  wire   [35:0] d14;
  wire   [35:0] hd_a15;
  wire   [35:0] d15;
  wire   [35:0] hd_a16;
  wire   [35:0] d16;
  wire   [35:0] hd_a17;
  wire   [35:0] d17;
  wire   [35:0] hd_a18;
  wire   [35:0] d18;
  wire   [35:0] hd_a19;
  wire   [35:0] d19;
  wire   [35:0] hd_a20;
  wire   [35:0] d20;
  wire   [35:0] hd_a21;
  wire   [35:0] d21;
  wire   [35:0] hd_a22;
  wire   [35:0] d22;
  wire   [35:0] hd_a23;
  wire   [35:0] d23;
  wire   [35:0] hd_a24;
  wire   [35:0] d24;
  wire   [35:0] hd_a25;
  wire   [35:0] d25;
  wire   [35:0] hd_a26;
  wire   [35:0] d26;
  wire   [35:0] hd_a27;
  wire   [35:0] d27;
  wire   [35:0] hd_a28;
  wire   [35:0] d28;
  wire   [35:0] hd_a29;
  wire   [35:0] d29;
  wire   [35:0] hd_a30;
  wire   [35:0] d30;
  wire   [31:0] hd_a31;
  wire   [31:0] d31;
  wire   [31:16] hd_a32;
  wire   [31:16] d32;
  wire   [3:0] counter;
  wire   [15:0] BF2I_a_xr_n;
  wire   [15:0] BF2I_a_er_n;
  wire   [15:0] BF2II_a_er_n;
  wire   [15:0] BF2II_a_ei_n;
  wire   [16:11] multiplier_r;
  wire   [14:11] multiplier_i;
  wire   [31:0] result_r;
  wire   [31:0] result_i;
  wire   [31:0] BF2I_b_xr_n;
  wire   [31:0] BF2I_b_xi_n;
  wire   [31:0] BF2I_b_er_n;
  wire   [31:0] BF2I_b_ei_n;
  wire   [31:0] BF2II_b_xr_n;
  wire   [31:0] BF2II_b_xi_n;
  wire   [31:0] fft_d15_q;
  wire   [31:0] fft_d;

  FAS_DW01_add_0 r1319 ( .A({U3_U8_Z_31, U3_U8_Z_30, U3_U8_Z_29, U3_U8_Z_28, 
        U3_U8_Z_27, U3_U8_Z_26, U3_U8_Z_25, U3_U8_Z_24, U3_U8_Z_23, U3_U8_Z_22, 
        U3_U8_Z_21, U3_U8_Z_20, U3_U8_Z_19, U3_U8_Z_18, U3_U8_Z_17, U3_U8_Z_16, 
        U3_U8_Z_15, U3_U8_Z_14, U3_U8_Z_13, U3_U8_Z_12, U3_U8_Z_11, U3_U8_Z_10, 
        U3_U8_Z_9, U3_U8_Z_8, U3_U8_Z_7, U3_U8_Z_6, U3_U8_Z_5, U3_U8_Z_4, 
        U3_U8_Z_3, U3_U8_Z_2, U3_U8_Z_1, U3_U8_Z_0}), .B(BF2I_b_er_n), .SUM({
        N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, 
        N371, N370, N369, N368, N543, N542, N541, N540, N539, N538, N537, N536, 
        N535, N534, N533, N532, N531, N530, N529, N528}) );
  FAS_DW01_add_1 add_72 ( .B(d07), .SUM(hd_a08), .A_35_(hd08_35), .A_34_(
        hd08_35), .A_33_(hd08_35), .A_32_(hd08_35), .A_31_(hd08_35), .A_30_(
        hd08_35), .A_29_(hd08_35), .A_28_(hd08_35), .A_27_(hd08_35), .A_26_(
        hd08_35), .A_25_(hd08_35), .A_24_(hd08_35), .A_23_(hd08_35), .A_22_(
        hd08_35), .A_21_(hd08_35), .A_20_(hd08_20_), .A_19_(hd08_19_), .A_18_(
        hd08_18_), .A_17_(hd08_17_), .A_16_(hd08_16_), .A_15_(hd08_15_), 
        .A_14_(hd08_14_), .A_13_(hd08_13_), .A_12_(hd08_12_), .A_11_(hd08_11_), 
        .A_10_(hd08_10_), .A_9_(hd08_9_), .A_8_(hd08_8_), .A_7_(hd08_7_), 
        .A_6_(hd08_6_), .A_5_(hd08_5_), .A_4_(data[2]), .A_3_(data[1]), .A_2_(
        data[0]) );
  FAS_DW01_add_2 add_75 ( .B(d10), .SUM(hd_a11), .A_35_(hd11_35), .A_34_(
        hd11_35), .A_33_(hd11_35), .A_32_(hd11_35), .A_31_(hd11_35), .A_30_(
        hd11_35), .A_29_(hd11_35), .A_28_(hd11_35), .A_27_(hd11[27]), .A_26_(
        hd11[26]), .A_25_(hd11[25]), .A_24_(hd11[24]), .A_23_(hd11[23]), 
        .A_22_(hd11[22]), .A_21_(hd11[21]), .A_20_(hd11[20]), .A_19_(hd11[19]), 
        .A_18_(hd11[18]), .A_17_(hd11[17]), .A_16_(hd11[16]), .A_15_(hd11[15]), 
        .A_14_(hd11[14]), .A_13_(hd11[13]), .A_12_(hd11[12]), .A_11_(hd11[11]), 
        .A_10_(hd11[10]), .A_9_(hd11[9]), .A_8_(hd11[8]), .A_7_(hd11[7]), 
        .A_6_(hd11[6]), .A_5_(hd11[5]), .A_4_(hd11[4]), .A_3_(hd11[3]), .A_2_(
        hd11[2]), .A_1_(hd11[1]) );
  FAS_DW01_add_3 add_89 ( .B(d24), .SUM(hd_a25), .A_35_(hd08_35), .A_34_(
        hd08_35), .A_33_(hd08_35), .A_32_(hd08_35), .A_31_(hd08_35), .A_30_(
        hd08_35), .A_29_(hd08_35), .A_28_(hd08_35), .A_27_(hd08_35), .A_26_(
        hd08_35), .A_25_(hd08_35), .A_24_(hd08_35), .A_23_(hd08_35), .A_22_(
        hd08_35), .A_21_(hd08_35), .A_20_(hd08_20_), .A_19_(hd08_19_), .A_18_(
        hd08_18_), .A_17_(hd08_17_), .A_16_(hd08_16_), .A_15_(hd08_15_), 
        .A_14_(hd08_14_), .A_13_(hd08_13_), .A_12_(hd08_12_), .A_11_(hd08_11_), 
        .A_10_(hd08_10_), .A_9_(hd08_9_), .A_8_(hd08_8_), .A_7_(hd08_7_), 
        .A_6_(hd08_6_), .A_5_(hd08_5_), .A_4_(data[2]), .A_3_(data[1]), .A_2_(
        data[0]) );
  FAS_DW01_add_4 add_84 ( .B(d19), .SUM(hd_a20), .A_35_(hd13_35), .A_34_(
        hd13_35), .A_33_(hd13_35), .A_32_(hd13_35), .A_31_(hd13_35), .A_30_(
        hd13_35), .A_29_(hd13_35), .A_28_(hd13_35), .A_27_(hd13[27]), .A_26_(
        hd13[26]), .A_25_(hd13[25]), .A_24_(hd13[24]), .A_23_(hd13[23]), 
        .A_22_(hd13[22]), .A_21_(hd13[21]), .A_20_(hd13[20]), .A_19_(hd13[19]), 
        .A_18_(hd13[18]), .A_17_(hd13[17]), .A_16_(hd13[16]), .A_15_(hd13[15]), 
        .A_14_(hd13[14]), .A_13_(hd13[13]), .A_12_(hd13[12]), .A_11_(hd13[11]), 
        .A_10_(hd13[10]), .A_9_(hd13[9]), .A_8_(hd13[8]), .A_7_(hd13[7]), 
        .A_6_(hd13[6]), .A_5_(hd13[5]), .A_4_(hd13[4]), .A_3_(hd13[3]), .A_2_(
        hd13[2]), .A_1_(hd13[1]) );
  FAS_DW01_add_5 add_92 ( .A({hd05_35, hd05_35, hd05_35, hd05_35, hd05_35, 
        hd05_35, hd05_35, hd05_35, hd05_35, hd05_35, hd05_35, hd05}), .B(d27), 
        .SUM(hd_a28) );
  FAS_DW01_add_6 add_95 ( .A_31_(hd02_35), .A_30_(hd02_35), .A_29_(hd02_35), 
        .A_28_(hd02_35), .A_27_(hd02_35), .A_26_(hd02_35), .A_25_(hd02_35), 
        .A_24_(hd02_35), .A_23_(hd02_35), .A_22_(hd02[22]), .A_21_(hd02[21]), 
        .A_20_(hd02[20]), .A_19_(hd02[19]), .A_18_(hd02[18]), .A_17_(hd02[17]), 
        .A_16_(hd02[16]), .A_15_(hd02[15]), .A_14_(hd02[14]), .A_13_(hd02[13]), 
        .A_12_(hd02[12]), .A_11_(hd02[11]), .A_10_(hd02[10]), .A_9_(hd02[9]), 
        .A_8_(hd02[8]), .A_7_(hd02[7]), .A_6_(hd02[6]), .A_5_(hd02[5]), .A_4_(
        hd02[4]), .A_3_(hd02[3]), .A_2_(hd02[2]), .A_1_(hd02[1]), .B_31_(
        d30[31]), .B_30_(d30[30]), .B_29_(d30[29]), .B_28_(d30[28]), .B_27_(
        d30[27]), .B_26_(d30[26]), .B_25_(d30[25]), .B_24_(d30[24]), .B_23_(
        d30[23]), .B_22_(d30[22]), .B_21_(d30[21]), .B_20_(d30[20]), .B_19_(
        d30[19]), .B_18_(d30[18]), .B_17_(d30[17]), .B_16_(d30[16]), .B_15_(
        d30[15]), .B_14_(d30[14]), .B_13_(d30[13]), .B_12_(d30[12]), .B_11_(
        d30[11]), .B_10_(d30[10]), .B_9_(d30[9]), .B_8_(d30[8]), .B_7_(d30[7]), 
        .B_6_(d30[6]), .B_5_(d30[5]), .B_4_(d30[4]), .B_3_(d30[3]), .B_2_(
        d30[2]), .B_1_(d30[1]), .B_0_(d30[0]), .SUM_31_(hd_a31[31]), .SUM_30_(
        hd_a31[30]), .SUM_29_(hd_a31[29]), .SUM_28_(hd_a31[28]), .SUM_27_(
        hd_a31[27]), .SUM_26_(hd_a31[26]), .SUM_25_(hd_a31[25]), .SUM_24_(
        hd_a31[24]), .SUM_23_(hd_a31[23]), .SUM_22_(hd_a31[22]), .SUM_21_(
        hd_a31[21]), .SUM_20_(hd_a31[20]), .SUM_19_(hd_a31[19]), .SUM_18_(
        hd_a31[18]), .SUM_17_(hd_a31[17]), .SUM_16_(hd_a31[16]), .SUM_15_(
        hd_a31[15]), .SUM_14_(hd_a31[14]), .SUM_13_(hd_a31[13]), .SUM_12_(
        hd_a31[12]), .SUM_11_(hd_a31[11]), .SUM_10_(hd_a31[10]), .SUM_9_(
        hd_a31[9]), .SUM_8_(hd_a31[8]), .SUM_7_(hd_a31[7]), .SUM_6_(hd_a31[6]), 
        .SUM_5_(hd_a31[5]), .SUM_4_(hd_a31[4]), .SUM_3_(hd_a31[3]), .SUM_2_(
        hd_a31[2]), .SUM_1_(hd_a31[1]), .SUM_0_(hd_a31[0]) );
  FAS_DW01_add_7 add_80 ( .A({hd16_35, hd16_35, hd16_35, hd16_35, hd16_35, 
        hd16_35, hd16}), .B(d15), .SUM(hd_a16) );
  FAS_DW01_addsub_2 r1284 ( .A({U3_U3_Z_15, U3_U3_Z_14, U3_U3_Z_13, U3_U3_Z_12, 
        U3_U3_Z_11, U3_U3_Z_10, U3_U3_Z_9, U3_U3_Z_8, U3_U3_Z_7, U3_U3_Z_6, 
        U3_U3_Z_5, U3_U3_Z_4, U3_U3_Z_3, U3_U3_Z_2, U3_U3_Z_1, U3_U3_Z_0}), 
        .B(BF2I_a_er_n), .ADD_SUB(mult_add_355_aco_b), .SUM({N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97}) );
  FAS_DW01_add_8 add_74 ( .B(d09), .SUM(hd_a10), .A_35_(hd10_35), .A_34_(
        hd10_35), .A_33_(hd10_35), .A_32_(hd10_35), .A_31_(hd10_35), .A_30_(
        hd10_35), .A_29_(hd10_35), .A_28_(hd10_35), .A_27_(hd10[27]), .A_26_(
        hd10[26]), .A_25_(hd10[25]), .A_24_(hd10[24]), .A_23_(hd10[23]), 
        .A_22_(hd10[22]), .A_21_(hd10[21]), .A_20_(hd10[20]), .A_19_(hd10[19]), 
        .A_18_(hd10[18]), .A_17_(hd10[17]), .A_16_(hd10[16]), .A_15_(hd10[15]), 
        .A_14_(hd10[14]), .A_13_(hd10[13]), .A_12_(hd10[12]), .A_11_(hd10[11]), 
        .A_10_(hd10[10]), .A_9_(hd10[9]), .A_8_(hd10[8]), .A_7_(hd10[7]), 
        .A_6_(hd10[6]), .A_5_(hd10[5]), .A_4_(hd10[4]), .A_3_(hd10[3]), .A_2_(
        hd10[2]), .A_1_(hd10[1]) );
  FAS_DW01_add_9 add_87 ( .B(d22), .SUM(hd_a23), .A_35_(hd10_35), .A_34_(
        hd10_35), .A_33_(hd10_35), .A_32_(hd10_35), .A_31_(hd10_35), .A_30_(
        hd10_35), .A_29_(hd10_35), .A_28_(hd10_35), .A_27_(hd10[27]), .A_26_(
        hd10[26]), .A_25_(hd10[25]), .A_24_(hd10[24]), .A_23_(hd10[23]), 
        .A_22_(hd10[22]), .A_21_(hd10[21]), .A_20_(hd10[20]), .A_19_(hd10[19]), 
        .A_18_(hd10[18]), .A_17_(hd10[17]), .A_16_(hd10[16]), .A_15_(hd10[15]), 
        .A_14_(hd10[14]), .A_13_(hd10[13]), .A_12_(hd10[12]), .A_11_(hd10[11]), 
        .A_10_(hd10[10]), .A_9_(hd10[9]), .A_8_(hd10[8]), .A_7_(hd10[7]), 
        .A_6_(hd10[6]), .A_5_(hd10[5]), .A_4_(hd10[4]), .A_3_(hd10[3]), .A_2_(
        hd10[2]), .A_1_(hd10[1]) );
  FAS_DW01_add_10 add_67 ( .A({hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, 
        hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, 
        hd03}), .B(d02), .SUM(hd_a03) );
  FAS_DW01_add_11 add_82 ( .B(d17), .SUM(hd_a18), .A_35_(hd15_35), .A_34_(
        hd15_35), .A_33_(hd15_35), .A_32_(hd15_35), .A_31_(hd15_35), .A_30_(
        hd15_35), .A_29_(hd15[29]), .A_28_(hd15[28]), .A_27_(hd15[27]), 
        .A_26_(hd15[26]), .A_25_(hd15[25]), .A_24_(hd15[24]), .A_23_(hd15[23]), 
        .A_22_(hd15[22]), .A_21_(hd15[21]), .A_20_(hd15[20]), .A_19_(hd15[19]), 
        .A_18_(hd15[18]), .A_17_(hd15[17]), .A_16_(hd15[16]), .A_15_(hd15[15]), 
        .A_14_(hd15[14]), .A_13_(hd15[13]), .A_12_(hd15[12]), .A_11_(hd15[11]), 
        .A_10_(hd15[10]), .A_9_(hd15[9]), .A_8_(hd15[8]), .A_7_(hd15[7]), 
        .A_6_(hd15[6]), .A_5_(hd15[5]), .A_4_(hd15[4]), .A_3_(hd15[3]), .A_2_(
        hd15[2]), .A_1_(hd15[1]) );
  FAS_DW01_add_12 add_69 ( .A({hd05_35, hd05_35, hd05_35, hd05_35, hd05_35, 
        hd05_35, hd05_35, hd05_35, hd05_35, hd05_35, hd05_35, hd05}), .B(d04), 
        .SUM(hd_a05) );
  FAS_DW01_add_13 add_68 ( .A({hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, 
        hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, 
        hd04_35, hd04}), .B(d03), .SUM(hd_a04) );
  FAS_DW01_add_14 add_79 ( .B(d14), .SUM(hd_a15), .A_35_(hd15_35), .A_34_(
        hd15_35), .A_33_(hd15_35), .A_32_(hd15_35), .A_31_(hd15_35), .A_30_(
        hd15_35), .A_29_(hd15[29]), .A_28_(hd15[28]), .A_27_(hd15[27]), 
        .A_26_(hd15[26]), .A_25_(hd15[25]), .A_24_(hd15[24]), .A_23_(hd15[23]), 
        .A_22_(hd15[22]), .A_21_(hd15[21]), .A_20_(hd15[20]), .A_19_(hd15[19]), 
        .A_18_(hd15[18]), .A_17_(hd15[17]), .A_16_(hd15[16]), .A_15_(hd15[15]), 
        .A_14_(hd15[14]), .A_13_(hd15[13]), .A_12_(hd15[12]), .A_11_(hd15[11]), 
        .A_10_(hd15[10]), .A_9_(hd15[9]), .A_8_(hd15[8]), .A_7_(hd15[7]), 
        .A_6_(hd15[6]), .A_5_(hd15[5]), .A_4_(hd15[4]), .A_3_(hd15[3]), .A_2_(
        hd15[2]), .A_1_(hd15[1]) );
  FAS_DW01_add_15 add_77 ( .B(d12), .SUM(hd_a13), .A_35_(hd13_35), .A_34_(
        hd13_35), .A_33_(hd13_35), .A_32_(hd13_35), .A_31_(hd13_35), .A_30_(
        hd13_35), .A_29_(hd13_35), .A_28_(hd13_35), .A_27_(hd13[27]), .A_26_(
        hd13[26]), .A_25_(hd13[25]), .A_24_(hd13[24]), .A_23_(hd13[23]), 
        .A_22_(hd13[22]), .A_21_(hd13[21]), .A_20_(hd13[20]), .A_19_(hd13[19]), 
        .A_18_(hd13[18]), .A_17_(hd13[17]), .A_16_(hd13[16]), .A_15_(hd13[15]), 
        .A_14_(hd13[14]), .A_13_(hd13[13]), .A_12_(hd13[12]), .A_11_(hd13[11]), 
        .A_10_(hd13[10]), .A_9_(hd13[9]), .A_8_(hd13[8]), .A_7_(hd13[7]), 
        .A_6_(hd13[6]), .A_5_(hd13[5]), .A_4_(hd13[4]), .A_3_(hd13[3]), .A_2_(
        hd13[2]), .A_1_(hd13[1]) );
  FAS_DW01_sub_0 sub_507 ( .A(BF2I_b_xi_n), .B(result_i), .DIFF({N363, N362, 
        N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, 
        N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, 
        N337, N336, N335, N334, N333, N332}) );
  FAS_DW01_sub_1 r1248 ( .A(BF2II_b_xi_n), .B({U3_U7_Z_31, U3_U7_Z_30, 
        U3_U7_Z_29, U3_U7_Z_28, U3_U7_Z_27, U3_U7_Z_26, U3_U7_Z_25, U3_U7_Z_24, 
        U3_U7_Z_23, U3_U7_Z_22, U3_U7_Z_21, U3_U7_Z_20, U3_U7_Z_19, U3_U7_Z_18, 
        U3_U7_Z_17, U3_U7_Z_16, U3_U7_Z_15, U3_U7_Z_14, U3_U7_Z_13, U3_U7_Z_12, 
        U3_U7_Z_11, U3_U7_Z_10, U3_U7_Z_9, U3_U7_Z_8, U3_U7_Z_7, U3_U7_Z_6, 
        U3_U7_Z_5, U3_U7_Z_4, U3_U7_Z_3, U3_U7_Z_2, U3_U7_Z_1, U3_U7_Z_0}), 
        .DIFF({N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, 
        N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, 
        N441, N440, N439, N438, N437, N436, N435, N434, N433, N432}) );
  FAS_DW01_addsub_3 r1277 ( .A({U3_U6_Z_31, U3_U6_Z_30, U3_U6_Z_29, U3_U6_Z_28, 
        U3_U6_Z_27, U3_U6_Z_26, U3_U6_Z_25, U3_U6_Z_24, U3_U6_Z_23, U3_U6_Z_22, 
        U3_U6_Z_21, U3_U6_Z_20, U3_U6_Z_19, U3_U6_Z_18, U3_U6_Z_17, U3_U6_Z_16, 
        U3_U6_Z_15, U3_U6_Z_14, U3_U6_Z_13, U3_U6_Z_12, U3_U6_Z_11, U3_U6_Z_10, 
        U3_U6_Z_9, U3_U6_Z_8, U3_U6_Z_7, U3_U6_Z_6, U3_U6_Z_5, U3_U6_Z_4, 
        U3_U6_Z_3, U3_U6_Z_2, U3_U6_Z_1, U3_U6_Z_0}), .B(BF2I_b_ei_n), 
        .SUM_31_(N399), .SUM_30_(N398), .SUM_29_(N397), .SUM_28_(N396), 
        .SUM_27_(N395), .SUM_26_(N394), .SUM_25_(N393), .SUM_24_(N392), 
        .SUM_23_(N391), .SUM_22_(N390), .SUM_21_(N389), .SUM_20_(N388), 
        .SUM_19_(N387), .SUM_18_(N386), .SUM_17_(N385), .SUM_16_(N384) );
  FAS_DW01_add_16 add_81 ( .A({hd16_35, hd16_35, hd16_35, hd16_35, hd16_35, 
        hd16_35, hd16}), .B(d16), .SUM(hd_a17) );
  FAS_DW01_add_17 add_93 ( .A({hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, 
        hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, hd04_35, 
        hd04_35, hd04}), .B(d28), .SUM(hd_a29) );
  FAS_DW01_add_18 add_78 ( .B(d13), .SUM(hd_a14), .A_35_(hd14_35), .A_34_(
        hd14_35), .A_33_(hd14_35), .A_32_(hd14_35), .A_31_(hd14_35), .A_30_(
        hd14_35), .A_29_(hd14_35), .A_28_(hd14[28]), .A_27_(hd14[27]), .A_26_(
        hd14[26]), .A_25_(hd14[25]), .A_24_(hd14[24]), .A_23_(hd14[23]), 
        .A_22_(hd14[22]), .A_21_(hd14[21]), .A_20_(hd14[20]), .A_19_(hd14[19]), 
        .A_18_(hd14[18]), .A_17_(hd14[17]), .A_16_(hd14[16]), .A_15_(hd14[15]), 
        .A_14_(hd14[14]), .A_13_(hd14[13]), .A_12_(hd14[12]), .A_11_(hd14[11]), 
        .A_10_(hd14[10]), .A_9_(hd14[9]), .A_8_(hd14[8]), .A_7_(hd14[7]), 
        .A_6_(hd14[6]), .A_5_(hd14[5]), .A_4_(hd14[4]), .A_3_(hd14[3]), .A_2_(
        hd14[2]) );
  FAS_DW01_add_19 add_91 ( .B(d26), .SUM(hd_a27), .A_35_(hd06_35), .A_34_(
        hd06_35), .A_33_(hd06_35), .A_32_(hd06_35), .A_31_(hd06_35), .A_30_(
        hd06_35), .A_29_(hd06_35), .A_28_(hd06_35), .A_27_(hd06_35), .A_26_(
        hd06_35), .A_25_(hd06[25]), .A_24_(hd06[24]), .A_23_(hd06[23]), 
        .A_22_(hd06[22]), .A_21_(hd06[21]), .A_20_(hd06[20]), .A_19_(hd06[19]), 
        .A_18_(hd06[18]), .A_17_(hd06[17]), .A_16_(hd06[16]), .A_15_(hd06[15]), 
        .A_14_(hd06[14]), .A_13_(hd06[13]), .A_12_(hd06[12]), .A_11_(hd06[11]), 
        .A_10_(hd06[10]), .A_9_(hd06[9]), .A_8_(hd06[8]), .A_7_(hd06[7]), 
        .A_6_(hd06[6]), .A_5_(hd06[5]), .A_4_(hd06[4]), .A_3_(hd06[3]), .A_2_(
        hd06[2]), .A_1_(hd06[1]) );
  FAS_DW01_add_20 add_66 ( .A_35_(hd02_35), .A_34_(hd02_35), .A_33_(hd02_35), 
        .A_32_(hd02_35), .A_31_(hd02_35), .A_30_(hd02_35), .A_29_(hd02_35), 
        .A_28_(hd02_35), .A_27_(hd02_35), .A_26_(hd02_35), .A_25_(hd02_35), 
        .A_24_(hd02_35), .A_23_(hd02_35), .A_22_(hd02[22]), .A_21_(hd02[21]), 
        .A_20_(hd02[20]), .A_19_(hd02[19]), .A_18_(hd02[18]), .A_17_(hd02[17]), 
        .A_16_(hd02[16]), .A_15_(hd02[15]), .A_14_(hd02[14]), .A_13_(hd02[13]), 
        .A_12_(hd02[12]), .A_11_(hd02[11]), .A_10_(hd02[10]), .A_9_(hd02[9]), 
        .A_8_(hd02[8]), .A_7_(hd02[7]), .A_6_(hd02[6]), .A_5_(hd02[5]), .A_4_(
        hd02[4]), .A_3_(hd02[3]), .A_2_(hd02[2]), .A_1_(hd02[1]), .B_35_(
        d01[35]), .B_34_(d01[34]), .B_33_(d01[33]), .B_32_(d01[32]), .B_31_(
        d01[31]), .B_30_(d01[30]), .B_29_(d01[29]), .B_28_(d01[28]), .B_27_(
        d01[27]), .B_26_(d01[26]), .B_25_(d01[25]), .B_24_(d01[24]), .B_23_(
        d01[23]), .B_22_(d01[22]), .B_21_(d01[21]), .B_20_(d01[20]), .B_19_(
        d01[19]), .B_18_(d01[18]), .B_17_(d01[17]), .B_16_(d01[16]), .B_15_(
        d01[15]), .B_14_(d01[14]), .B_13_(d01[13]), .B_12_(d01[12]), .B_11_(
        d01[11]), .B_10_(d01[10]), .B_9_(d01[9]), .B_8_(d01[8]), .B_7_(d01[7]), 
        .B_6_(d01[6]), .B_5_(d01[5]), .B_4_(d01[4]), .B_3_(d01[3]), .B_2_(
        d01[2]), .B_1_(d01[1]), .SUM_35_(hd_a02[35]), .SUM_34_(hd_a02[34]), 
        .SUM_33_(hd_a02[33]), .SUM_32_(hd_a02[32]), .SUM_31_(hd_a02[31]), 
        .SUM_30_(hd_a02[30]), .SUM_29_(hd_a02[29]), .SUM_28_(hd_a02[28]), 
        .SUM_27_(hd_a02[27]), .SUM_26_(hd_a02[26]), .SUM_25_(hd_a02[25]), 
        .SUM_24_(hd_a02[24]), .SUM_23_(hd_a02[23]), .SUM_22_(hd_a02[22]), 
        .SUM_21_(hd_a02[21]), .SUM_20_(hd_a02[20]), .SUM_19_(hd_a02[19]), 
        .SUM_18_(hd_a02[18]), .SUM_17_(hd_a02[17]), .SUM_16_(hd_a02[16]), 
        .SUM_15_(hd_a02[15]), .SUM_14_(hd_a02[14]), .SUM_13_(hd_a02[13]), 
        .SUM_12_(hd_a02[12]), .SUM_11_(hd_a02[11]), .SUM_10_(hd_a02[10]), 
        .SUM_9_(hd_a02[9]), .SUM_8_(hd_a02[8]), .SUM_7_(hd_a02[7]), .SUM_6_(
        hd_a02[6]), .SUM_5_(hd_a02[5]), .SUM_4_(hd_a02[4]), .SUM_3_(hd_a02[3]), 
        .SUM_2_(hd_a02[2]), .SUM_1_(hd_a02[1]) );
  FAS_DW01_add_21 add_83 ( .B(d18), .SUM(hd_a19), .A_35_(hd14_35), .A_34_(
        hd14_35), .A_33_(hd14_35), .A_32_(hd14_35), .A_31_(hd14_35), .A_30_(
        hd14_35), .A_29_(hd14_35), .A_28_(hd14[28]), .A_27_(hd14[27]), .A_26_(
        hd14[26]), .A_25_(hd14[25]), .A_24_(hd14[24]), .A_23_(hd14[23]), 
        .A_22_(hd14[22]), .A_21_(hd14[21]), .A_20_(hd14[20]), .A_19_(hd14[19]), 
        .A_18_(hd14[18]), .A_17_(hd14[17]), .A_16_(hd14[16]), .A_15_(hd14[15]), 
        .A_14_(hd14[14]), .A_13_(hd14[13]), .A_12_(hd14[12]), .A_11_(hd14[11]), 
        .A_10_(hd14[10]), .A_9_(hd14[9]), .A_8_(hd14[8]), .A_7_(hd14[7]), 
        .A_6_(hd14[6]), .A_5_(hd14[5]), .A_4_(hd14[4]), .A_3_(hd14[3]), .A_2_(
        hd14[2]) );
  FAS_DW01_add_22 add_76 ( .B(d11), .SUM(hd_a12), .A_35_(hd12_35), .A_34_(
        hd12_35), .A_33_(hd12_35), .A_32_(hd12_35), .A_31_(hd12_35), .A_30_(
        hd12_35), .A_29_(hd12_35), .A_28_(hd12_35), .A_27_(hd12_35), .A_26_(
        hd12_35), .A_25_(hd12[25]), .A_24_(hd12[24]), .A_23_(hd12[23]), 
        .A_22_(hd12[22]), .A_21_(hd12[21]), .A_20_(hd12[20]), .A_19_(hd12[19]), 
        .A_18_(hd12[18]), .A_17_(hd12[17]), .A_16_(hd12[16]), .A_15_(hd12[15]), 
        .A_14_(hd12[14]), .A_13_(hd12[13]), .A_12_(hd12[12]), .A_11_(hd12[11]), 
        .A_10_(hd12[10]), .A_9_(hd12[9]), .A_8_(hd12[8]), .A_7_(hd12[7]), 
        .A_6_(hd12[6]), .A_5_(hd12[5]), .A_4_(hd12[4]), .A_3_(hd12[3]), .A_2_(
        hd12[2]) );
  FAS_DW01_add_23 add_85 ( .B(d20), .SUM(hd_a21), .A_35_(hd12_35), .A_34_(
        hd12_35), .A_33_(hd12_35), .A_32_(hd12_35), .A_31_(hd12_35), .A_30_(
        hd12_35), .A_29_(hd12_35), .A_28_(hd12_35), .A_27_(hd12_35), .A_26_(
        hd12_35), .A_25_(hd12[25]), .A_24_(hd12[24]), .A_23_(hd12[23]), 
        .A_22_(hd12[22]), .A_21_(hd12[21]), .A_20_(hd12[20]), .A_19_(hd12[19]), 
        .A_18_(hd12[18]), .A_17_(hd12[17]), .A_16_(hd12[16]), .A_15_(hd12[15]), 
        .A_14_(hd12[14]), .A_13_(hd12[13]), .A_12_(hd12[12]), .A_11_(hd12[11]), 
        .A_10_(hd12[10]), .A_9_(hd12[9]), .A_8_(hd12[8]), .A_7_(hd12[7]), 
        .A_6_(hd12[6]), .A_5_(hd12[5]), .A_4_(hd12[4]), .A_3_(hd12[3]), .A_2_(
        hd12[2]) );
  FAS_DW01_add_24 add_94 ( .A({hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, 
        hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, hd03_35, 
        hd03}), .B(d29), .SUM(hd_a30) );
  FAS_DW01_add_25 add_88 ( .A({hd09_35, hd09_35, hd09_35, hd09_35, hd09_35, 
        hd09_35, hd09_35, hd09_35, hd09_35, hd09}), .B(d23), .SUM(hd_a24) );
  FAS_DW01_add_26 add_71 ( .B(d06), .SUM(hd_a07), .A_35_(hd07_35), .A_34_(
        hd07_35), .A_33_(hd07_35), .A_32_(hd07_35), .A_31_(hd07_35), .A_30_(
        hd07_35), .A_29_(hd07_35), .A_28_(hd07_35), .A_27_(hd07_35), .A_26_(
        hd07_35), .A_25_(hd07[25]), .A_24_(hd07[24]), .A_23_(hd07[23]), 
        .A_22_(hd07[22]), .A_21_(hd07[21]), .A_20_(hd07[20]), .A_19_(hd07[19]), 
        .A_18_(hd07[18]), .A_17_(hd07[17]), .A_16_(hd07[16]), .A_15_(hd07[15]), 
        .A_14_(hd07[14]), .A_13_(hd07[13]), .A_12_(hd07[12]), .A_11_(hd07[11]), 
        .A_10_(hd07[10]), .A_9_(hd07[9]), .A_8_(hd07[8]), .A_7_(hd07[7]), 
        .A_6_(hd07[6]), .A_5_(hd07[5]), .A_4_(hd07[4]), .A_3_(hd07[3]), .A_2_(
        hd07[2]), .A_1_(hd07[1]) );
  FAS_DW01_add_27 add_86 ( .B(d21), .SUM(hd_a22), .A_35_(hd11_35), .A_34_(
        hd11_35), .A_33_(hd11_35), .A_32_(hd11_35), .A_31_(hd11_35), .A_30_(
        hd11_35), .A_29_(hd11_35), .A_28_(hd11_35), .A_27_(hd11[27]), .A_26_(
        hd11[26]), .A_25_(hd11[25]), .A_24_(hd11[24]), .A_23_(hd11[23]), 
        .A_22_(hd11[22]), .A_21_(hd11[21]), .A_20_(hd11[20]), .A_19_(hd11[19]), 
        .A_18_(hd11[18]), .A_17_(hd11[17]), .A_16_(hd11[16]), .A_15_(hd11[15]), 
        .A_14_(hd11[14]), .A_13_(hd11[13]), .A_12_(hd11[12]), .A_11_(hd11[11]), 
        .A_10_(hd11[10]), .A_9_(hd11[9]), .A_8_(hd11[8]), .A_7_(hd11[7]), 
        .A_6_(hd11[6]), .A_5_(hd11[5]), .A_4_(hd11[4]), .A_3_(hd11[3]), .A_2_(
        hd11[2]), .A_1_(hd11[1]) );
  FAS_DW01_sub_2 sub_281 ( .A(BF2I_a_xr_n), .B(fir_d), .DIFF({N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76}) );
  FAS_DW01_add_28 add_96 ( .A_31_(hd01_35), .A_30_(hd01_35), .A_29_(hd01_35), 
        .A_28_(hd01_35), .A_27_(hd01_35), .A_26_(hd01_35), .A_25_(hd01_35), 
        .A_24_(hd01_35), .A_23_(hd01_35), .A_22_(hd01[22]), .A_21_(hd01[21]), 
        .A_20_(hd01[20]), .A_19_(hd01[19]), .A_18_(hd01[18]), .A_17_(hd01[17]), 
        .A_16_(hd01[16]), .A_15_(hd01[15]), .A_14_(hd01[14]), .A_13_(hd01[13]), 
        .A_12_(hd01[12]), .A_11_(hd01[11]), .A_10_(hd01[10]), .A_9_(hd01[9]), 
        .A_8_(hd01[8]), .A_7_(hd01[7]), .A_6_(hd01[6]), .A_5_(hd01[5]), .A_4_(
        hd01[4]), .A_3_(hd01[3]), .A_2_(hd01[2]), .A_1_(hd01[1]), .B_31_(
        d31[31]), .B_30_(d31[30]), .B_29_(d31[29]), .B_28_(d31[28]), .B_27_(
        d31[27]), .B_26_(d31[26]), .B_25_(d31[25]), .B_24_(d31[24]), .B_23_(
        d31[23]), .B_22_(d31[22]), .B_21_(d31[21]), .B_20_(d31[20]), .B_19_(
        d31[19]), .B_18_(d31[18]), .B_17_(d31[17]), .B_16_(d31[16]), .B_15_(
        d31[15]), .B_14_(d31[14]), .B_13_(d31[13]), .B_12_(d31[12]), .B_11_(
        d31[11]), .B_10_(d31[10]), .B_9_(d31[9]), .B_8_(d31[8]), .B_7_(d31[7]), 
        .B_6_(d31[6]), .B_5_(d31[5]), .B_4_(d31[4]), .B_3_(d31[3]), .B_2_(
        d31[2]), .B_1_(d31[1]), .SUM_31_(hd_a32[31]), .SUM_30_(hd_a32[30]), 
        .SUM_29_(hd_a32[29]), .SUM_28_(hd_a32[28]), .SUM_27_(hd_a32[27]), 
        .SUM_26_(hd_a32[26]), .SUM_25_(hd_a32[25]), .SUM_24_(hd_a32[24]), 
        .SUM_23_(hd_a32[23]), .SUM_22_(hd_a32[22]), .SUM_21_(hd_a32[21]), 
        .SUM_20_(hd_a32[20]), .SUM_19_(hd_a32[19]), .SUM_18_(hd_a32[18]), 
        .SUM_17_(hd_a32[17]), .SUM_16_(hd_a32[16]) );
  FAS_DW01_add_29 add_90 ( .B(d25), .SUM(hd_a26), .A_35_(hd07_35), .A_34_(
        hd07_35), .A_33_(hd07_35), .A_32_(hd07_35), .A_31_(hd07_35), .A_30_(
        hd07_35), .A_29_(hd07_35), .A_28_(hd07_35), .A_27_(hd07_35), .A_26_(
        hd07_35), .A_25_(hd07[25]), .A_24_(hd07[24]), .A_23_(hd07[23]), 
        .A_22_(hd07[22]), .A_21_(hd07[21]), .A_20_(hd07[20]), .A_19_(hd07[19]), 
        .A_18_(hd07[18]), .A_17_(hd07[17]), .A_16_(hd07[16]), .A_15_(hd07[15]), 
        .A_14_(hd07[14]), .A_13_(hd07[13]), .A_12_(hd07[12]), .A_11_(hd07[11]), 
        .A_10_(hd07[10]), .A_9_(hd07[9]), .A_8_(hd07[8]), .A_7_(hd07[7]), 
        .A_6_(hd07[6]), .A_5_(hd07[5]), .A_4_(hd07[4]), .A_3_(hd07[3]), .A_2_(
        hd07[2]), .A_1_(hd07[1]) );
  FAS_DW01_add_30 add_73 ( .A({hd09_35, hd09_35, hd09_35, hd09_35, hd09_35, 
        hd09_35, hd09_35, hd09_35, hd09_35, hd09}), .B(d08), .SUM(hd_a09) );
  FAS_DW01_sub_3 sub_506 ( .A(BF2I_b_xr_n), .B(result_r), .DIFF({N331, N330, 
        N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, 
        N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, 
        N305, N304, N303, N302, N301, N300}) );
  FAS_DW01_sub_4 r59 ( .A(BF2II_b_xr_n), .B({U3_U5_Z_31, U3_U5_Z_30, 
        U3_U5_Z_29, U3_U5_Z_28, U3_U5_Z_27, U3_U5_Z_26, U3_U5_Z_25, U3_U5_Z_24, 
        U3_U5_Z_23, U3_U5_Z_22, U3_U5_Z_21, U3_U5_Z_20, U3_U5_Z_19, U3_U5_Z_18, 
        U3_U5_Z_17, U3_U5_Z_16, U3_U5_Z_15, U3_U5_Z_14, U3_U5_Z_13, U3_U5_Z_12, 
        U3_U5_Z_11, U3_U5_Z_10, U3_U5_Z_9, U3_U5_Z_8, U3_U5_Z_7, U3_U5_Z_6, 
        U3_U5_Z_5, U3_U5_Z_4, U3_U5_Z_3, U3_U5_Z_2, U3_U5_Z_1, U3_U5_Z_0}), 
        .DIFF({N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, 
        N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, 
        N409, N408, N407, N406, N405, N404, N403, N402, N401, N400}) );
  FAS_DW01_add_31 add_505_aco ( .A(BF2I_b_xi_n), .B({N1426, N1425, N1424, 
        N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, 
        N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, 
        N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395}), .SUM(
        BF2I_b_ei_n) );
  FAS_DW01_add_32 add_433 ( .A({N257, N256, N255, N254, N253, N252, N251, N250, 
        N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, 
        N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226}), .B({N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, 
        N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, 
        N265, N264, N263, N262, N261, N260, N259, N258}), .SUM(result_i) );
  FAS_DW01_add_33 add_504_aco ( .A(BF2I_b_xr_n), .B({N1458, N1457, N1456, 
        N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, 
        N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, 
        N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427}), .SUM(
        BF2I_b_er_n) );
  FAS_DW01_sub_5 sub_432 ( .A({N193, N192, N191, N190, N189, N188, N187, N186, 
        N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, 
        N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162}), .B({N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, 
        N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, 
        N201, N200, N199, N198, N197, N196, N195, N194}), .DIFF(result_r) );
  FAS_DW01_sub_6 sub_363_aco ( .A({N128, N127, N126, N125, N124, N123, N122, 
        N121, N120, N119, N118, N117, N116, N115, N114, N113}), .B({N1394, 
        N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, 
        N1383, N1382, N1381, N1380, N1379}), .DIFF(BF2II_a_ei_n) );
  FAS_DW01_add_34 add_355_aco ( .A({N145, N144, N143, N142, N141, N140, N139, 
        N138, N137, N136, N135, N134, N133, N132, N131, N130}), .B({N1378, 
        N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, 
        N1367, N1366, N1365, N1364, N1363}), .SUM(BF2II_a_er_n) );
  FAS_DW01_add_35 add_280_aco ( .A(BF2I_a_xr_n), .B({N1362, N1361, N1360, 
        N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, 
        N1349, N1348, N1347}), .SUM(BF2I_a_er_n) );
  FAS_DW01_inc_1 add_100_S2 ( .A({n11218, d32[30:16]}), .SUM({N43, N42, N41, 
        N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28}) );
  FAS_DW01_add_36 add_70 ( .B(d05), .SUM(hd_a06), .A_35_(hd06_35), .A_34_(
        hd06_35), .A_33_(hd06_35), .A_32_(hd06_35), .A_31_(hd06_35), .A_30_(
        hd06_35), .A_29_(hd06_35), .A_28_(hd06_35), .A_27_(hd06_35), .A_26_(
        hd06_35), .A_25_(hd06[25]), .A_24_(hd06[24]), .A_23_(hd06[23]), 
        .A_22_(hd06[22]), .A_21_(hd06[21]), .A_20_(hd06[20]), .A_19_(hd06[19]), 
        .A_18_(hd06[18]), .A_17_(hd06[17]), .A_16_(hd06[16]), .A_15_(hd06[15]), 
        .A_14_(hd06[14]), .A_13_(hd06[13]), .A_12_(hd06[12]), .A_11_(hd06[11]), 
        .A_10_(hd06[10]), .A_9_(hd06[9]), .A_8_(hd06[8]), .A_7_(hd06[7]), 
        .A_6_(hd06[6]), .A_5_(hd06[5]), .A_4_(hd06[4]), .A_3_(hd06[3]), .A_2_(
        hd06[2]), .A_1_(hd06[1]) );
  FAS_DW01_add_37 add_790 ( .SUM(fft_d), .A_31_(N1112), .A_30_(N1111), .A_29_(
        N1110), .A_28_(N1109), .A_27_(N1108), .A_26_(N1107), .A_25_(N1106), 
        .A_24_(N1105), .A_23_(N1104), .A_22_(N1103), .A_21_(N1102), .A_20_(
        N1101), .A_19_(N1100), .A_18_(N1099), .A_17_(N1098), .A_16_(N1097), 
        .A_15_(N1096), .A_14_(N1095), .A_13_(N1094), .A_12_(N1093), .A_11_(
        N1092), .A_10_(N1091), .A_9_(N1090), .A_8_(N1089), .A_7_(N1088), 
        .A_6_(N1087), .A_5_(N1086), .A_4_(N1085), .A_3_(N1084), .A_2_(N1083), 
        .A_0_(N1081), .B_31_(N1144), .B_30_(N1143), .B_29_(N1142), .B_28_(
        N1141), .B_27_(N1140), .B_26_(N1139), .B_25_(N1138), .B_24_(N1137), 
        .B_23_(N1136), .B_22_(N1135), .B_21_(N1134), .B_20_(N1133), .B_19_(
        N1132), .B_18_(N1131), .B_17_(N1130), .B_16_(N1129), .B_15_(N1128), 
        .B_14_(N1127), .B_13_(N1126), .B_12_(N1125), .B_11_(N1124), .B_10_(
        N1123), .B_9_(N1122), .B_8_(N1121), .B_7_(N1120), .B_6_(N1119), .B_5_(
        N1118), .B_4_(N1117), .B_3_(N1116), .B_2_(N1115), .B_0_(N1113) );
  FAS_DW_mult_tc_22 mult_790 ( .a(fft_d15_q[31:16]), .product_31_(N1112), 
        .product_30_(N1111), .product_29_(N1110), .product_28_(N1109), 
        .product_27_(N1108), .product_26_(N1107), .product_25_(N1106), 
        .product_24_(N1105), .product_23_(N1104), .product_22_(N1103), 
        .product_21_(N1102), .product_20_(N1101), .product_19_(N1100), 
        .product_18_(N1099), .product_17_(N1098), .product_16_(N1097), 
        .product_15_(N1096), .product_14_(N1095), .product_13_(N1094), 
        .product_12_(N1093), .product_11_(N1092), .product_10_(N1091), 
        .product_9_(N1090), .product_8_(N1089), .product_7_(N1088), 
        .product_6_(N1087), .product_5_(N1086), .product_4_(N1085), 
        .product_3_(N1084), .product_2_(N1083), .product_0_(N1081) );
  FAS_DW_mult_tc_23 mult_790_2 ( .a(fft_d15_q[15:0]), .product_31_(N1144), 
        .product_30_(N1143), .product_29_(N1142), .product_28_(N1141), 
        .product_27_(N1140), .product_26_(N1139), .product_25_(N1138), 
        .product_24_(N1137), .product_23_(N1136), .product_22_(N1135), 
        .product_21_(N1134), .product_20_(N1133), .product_19_(N1132), 
        .product_18_(N1131), .product_17_(N1130), .product_16_(N1129), 
        .product_15_(N1128), .product_14_(N1127), .product_13_(N1126), 
        .product_12_(N1125), .product_11_(N1124), .product_10_(N1123), 
        .product_9_(N1122), .product_8_(N1121), .product_7_(N1120), 
        .product_6_(N1119), .product_5_(N1118), .product_4_(N1117), 
        .product_3_(N1116), .product_2_(N1115), .product_0_(N1113) );
  FAS_DW_mult_tc_24 mult_37 ( .a(data), .product_26_(hd06_35), .product_25_(
        hd06[25]), .product_24_(hd06[24]), .product_23_(hd06[23]), 
        .product_22_(hd06[22]), .product_21_(hd06[21]), .product_20_(hd06[20]), 
        .product_19_(hd06[19]), .product_18_(hd06[18]), .product_17_(hd06[17]), 
        .product_16_(hd06[16]), .product_15_(hd06[15]), .product_14_(hd06[14]), 
        .product_13_(hd06[13]), .product_12_(hd06[12]), .product_11_(hd06[11]), 
        .product_10_(hd06[10]), .product_9_(hd06[9]), .product_8_(hd06[8]), 
        .product_7_(hd06[7]), .product_6_(hd06[6]), .product_5_(hd06[5]), 
        .product_4_(hd06[4]), .product_3_(hd06[3]), .product_2_(hd06[2]), 
        .product_1_(hd06[1]) );
  FAS_DW_mult_tc_25 mult_432 ( .a(BF2II_a_er_n), .b_17_(multiplier_r_31), 
        .b_16_(multiplier_r[16]), .b_15_(multiplier_r[15]), .b_14_(
        multiplier_r[14]), .b_13_(multiplier_r[13]), .b_12_(multiplier_r[12]), 
        .b_11_(multiplier_r[11]), .b_10_(multiplier_r[15]), .b_9_(
        multiplier_r_31), .b_8_(multiplier_r_8), .b_7_(multiplier_r[14]), 
        .b_6_(multiplier_r_6), .b_5_(multiplier_r_6), .b_4_(multiplier_r_6), 
        .b_3_(multiplier_r_31), .b_2_(multiplier_i_6), .b_1_(multiplier_i[12]), 
        .b_0_(multiplier_i_0), .product_31_(N193), .product_30_(N192), 
        .product_29_(N191), .product_28_(N190), .product_27_(N189), 
        .product_26_(N188), .product_25_(N187), .product_24_(N186), 
        .product_23_(N185), .product_22_(N184), .product_21_(N183), 
        .product_20_(N182), .product_19_(N181), .product_18_(N180), 
        .product_17_(N179), .product_16_(N178), .product_15_(N177), 
        .product_14_(N176), .product_13_(N175), .product_12_(N174), 
        .product_11_(N173), .product_10_(N172), .product_9_(N171), 
        .product_8_(N170), .product_7_(N169), .product_6_(N168), .product_5_(
        N167), .product_4_(N166), .product_3_(N165), .product_2_(N164), 
        .product_1_(N163), .product_0_(N162) );
  FAS_DW_mult_tc_26 mult_432_2 ( .a(BF2II_a_ei_n), .b_16_(multiplier_i_31), 
        .b_15_(n10479), .b_14_(multiplier_i[14]), .b_13_(n10480), .b_12_(
        multiplier_i[12]), .b_11_(multiplier_i[11]), .b_10_(n10479), .b_9_(
        multiplier_i_9), .b_8_(multiplier_i_8), .b_7_(multiplier_i[14]), 
        .b_6_(multiplier_i_6), .b_5_(multiplier_i_6), .b_4_(multiplier_i_6), 
        .b_3_(multiplier_i_9), .b_2_(multiplier_i_6), .b_1_(n10480), .b_0_(
        multiplier_i_0), .product_31_(N225), .product_30_(N224), .product_29_(
        N223), .product_28_(N222), .product_27_(N221), .product_26_(N220), 
        .product_25_(N219), .product_24_(N218), .product_23_(N217), 
        .product_22_(N216), .product_21_(N215), .product_20_(N214), 
        .product_19_(N213), .product_18_(N212), .product_17_(N211), 
        .product_16_(N210), .product_15_(N209), .product_14_(N208), 
        .product_13_(N207), .product_12_(N206), .product_11_(N205), 
        .product_10_(N204), .product_9_(N203), .product_8_(N202), .product_7_(
        N201), .product_6_(N200), .product_5_(N199), .product_4_(N198), 
        .product_3_(N197), .product_2_(N196), .product_1_(N195), .product_0_(
        N194) );
  FAS_DW_mult_uns_5 mult_add_504_aco ( .a(result_r), .b(BF2I_b_s), 
        .product_31_(N1458), .product_30_(N1457), .product_29_(N1456), 
        .product_28_(N1455), .product_27_(N1454), .product_26_(N1453), 
        .product_25_(N1452), .product_24_(N1451), .product_23_(N1450), 
        .product_22_(N1449), .product_21_(N1448), .product_20_(N1447), 
        .product_19_(N1446), .product_18_(N1445), .product_17_(N1444), 
        .product_16_(N1443), .product_15_(N1442), .product_14_(N1441), 
        .product_13_(N1440), .product_12_(N1439), .product_11_(N1438), 
        .product_10_(N1437), .product_9_(N1436), .product_8_(N1435), 
        .product_7_(N1434), .product_6_(N1433), .product_5_(N1432), 
        .product_4_(N1431), .product_3_(N1430), .product_2_(N1429), 
        .product_1_(N1428), .product_0_(N1427) );
  FAS_DW_mult_tc_27 mult_433 ( .a(BF2II_a_ei_n), .b_17_(multiplier_r_31), 
        .b_16_(multiplier_r[16]), .b_15_(multiplier_r[15]), .b_14_(
        multiplier_r[14]), .b_13_(multiplier_r[13]), .b_12_(multiplier_r[12]), 
        .b_11_(multiplier_r[11]), .b_10_(multiplier_r[15]), .b_9_(
        multiplier_r_31), .b_8_(multiplier_r_8), .b_7_(multiplier_r[14]), 
        .b_6_(multiplier_r_6), .b_5_(multiplier_r_6), .b_4_(multiplier_r_6), 
        .b_3_(multiplier_r_31), .b_2_(multiplier_i_6), .b_1_(multiplier_i[12]), 
        .b_0_(multiplier_i_0), .product_31_(N257), .product_30_(N256), 
        .product_29_(N255), .product_28_(N254), .product_27_(N253), 
        .product_26_(N252), .product_25_(N251), .product_24_(N250), 
        .product_23_(N249), .product_22_(N248), .product_21_(N247), 
        .product_20_(N246), .product_19_(N245), .product_18_(N244), 
        .product_17_(N243), .product_16_(N242), .product_15_(N241), 
        .product_14_(N240), .product_13_(N239), .product_12_(N238), 
        .product_11_(N237), .product_10_(N236), .product_9_(N235), 
        .product_8_(N234), .product_7_(N233), .product_6_(N232), .product_5_(
        N231), .product_4_(N230), .product_3_(N229), .product_2_(N228), 
        .product_1_(N227), .product_0_(N226) );
  FAS_DW_mult_tc_28 mult_433_2 ( .a(BF2II_a_er_n), .b_16_(multiplier_i_31), 
        .b_15_(n10479), .b_14_(multiplier_i[14]), .b_13_(n10480), .b_12_(
        multiplier_i[12]), .b_11_(multiplier_i[11]), .b_10_(n10479), .b_9_(
        multiplier_i_9), .b_8_(multiplier_i_8), .b_7_(multiplier_i[14]), 
        .b_6_(multiplier_i_6), .b_5_(multiplier_i_6), .b_4_(multiplier_i_6), 
        .b_3_(multiplier_i_9), .b_2_(multiplier_i_6), .b_1_(n10480), .b_0_(
        multiplier_i_0), .product_31_(N289), .product_30_(N288), .product_29_(
        N287), .product_28_(N286), .product_27_(N285), .product_26_(N284), 
        .product_25_(N283), .product_24_(N282), .product_23_(N281), 
        .product_22_(N280), .product_21_(N279), .product_20_(N278), 
        .product_19_(N277), .product_18_(N276), .product_17_(N275), 
        .product_16_(N274), .product_15_(N273), .product_14_(N272), 
        .product_13_(N271), .product_12_(N270), .product_11_(N269), 
        .product_10_(N268), .product_9_(N267), .product_8_(N266), .product_7_(
        N265), .product_6_(N264), .product_5_(N263), .product_4_(N262), 
        .product_3_(N261), .product_2_(N260), .product_1_(N259), .product_0_(
        N258) );
  FAS_DW_mult_uns_6 mult_add_505_aco ( .a(result_i), .b(BF2I_b_s), 
        .product_31_(N1426), .product_30_(N1425), .product_29_(N1424), 
        .product_28_(N1423), .product_27_(N1422), .product_26_(N1421), 
        .product_25_(N1420), .product_24_(N1419), .product_23_(N1418), 
        .product_22_(N1417), .product_21_(N1416), .product_20_(N1415), 
        .product_19_(N1414), .product_18_(N1413), .product_17_(N1412), 
        .product_16_(N1411), .product_15_(N1410), .product_14_(N1409), 
        .product_13_(N1408), .product_12_(N1407), .product_11_(N1406), 
        .product_10_(N1405), .product_9_(N1404), .product_8_(N1403), 
        .product_7_(N1402), .product_6_(N1401), .product_5_(N1400), 
        .product_4_(N1399), .product_3_(N1398), .product_2_(N1397), 
        .product_1_(N1396), .product_0_(N1395) );
  FAS_DW_mult_tc_29 mult_33 ( .a(data), .product_23_(hd02_35), .product_22_(
        hd02[22]), .product_21_(hd02[21]), .product_20_(hd02[20]), 
        .product_19_(hd02[19]), .product_18_(hd02[18]), .product_17_(hd02[17]), 
        .product_16_(hd02[16]), .product_15_(hd02[15]), .product_14_(hd02[14]), 
        .product_13_(hd02[13]), .product_12_(hd02[12]), .product_11_(hd02[11]), 
        .product_10_(hd02[10]), .product_9_(hd02[9]), .product_8_(hd02[8]), 
        .product_7_(hd02[7]), .product_6_(hd02[6]), .product_5_(hd02[5]), 
        .product_4_(hd02[4]), .product_3_(hd02[3]), .product_2_(hd02[2]), 
        .product_1_(hd02[1]) );
  FAS_DW_mult_tc_30 mult_40 ( .a(data), .product({hd09_35, hd09}) );
  FAS_DW_mult_tc_31 mult_38 ( .a(data), .product_26_(hd07_35), .product_25_(
        hd07[25]), .product_24_(hd07[24]), .product_23_(hd07[23]), 
        .product_22_(hd07[22]), .product_21_(hd07[21]), .product_20_(hd07[20]), 
        .product_19_(hd07[19]), .product_18_(hd07[18]), .product_17_(hd07[17]), 
        .product_16_(hd07[16]), .product_15_(hd07[15]), .product_14_(hd07[14]), 
        .product_13_(hd07[13]), .product_12_(hd07[12]), .product_11_(hd07[11]), 
        .product_10_(hd07[10]), .product_9_(hd07[9]), .product_8_(hd07[8]), 
        .product_7_(hd07[7]), .product_6_(hd07[6]), .product_5_(hd07[5]), 
        .product_4_(hd07[4]), .product_3_(hd07[3]), .product_2_(hd07[2]), 
        .product_1_(hd07[1]) );
  FAS_DW_mult_tc_32 mult_32 ( .a(data), .product_23_(hd01_35), .product_22_(
        hd01[22]), .product_21_(hd01[21]), .product_20_(hd01[20]), 
        .product_19_(hd01[19]), .product_18_(hd01[18]), .product_17_(hd01[17]), 
        .product_16_(hd01[16]), .product_15_(hd01[15]), .product_14_(hd01[14]), 
        .product_13_(hd01[13]), .product_12_(hd01[12]), .product_11_(hd01[11]), 
        .product_10_(hd01[10]), .product_9_(hd01[9]), .product_8_(hd01[8]), 
        .product_7_(hd01[7]), .product_6_(hd01[6]), .product_5_(hd01[5]), 
        .product_4_(hd01[4]), .product_3_(hd01[3]), .product_2_(hd01[2]), 
        .product_1_(hd01[1]) );
  FAS_DW_mult_tc_33 mult_42 ( .a(data), .product_28_(hd11_35), .product_27_(
        hd11[27]), .product_26_(hd11[26]), .product_25_(hd11[25]), 
        .product_24_(hd11[24]), .product_23_(hd11[23]), .product_22_(hd11[22]), 
        .product_21_(hd11[21]), .product_20_(hd11[20]), .product_19_(hd11[19]), 
        .product_18_(hd11[18]), .product_17_(hd11[17]), .product_16_(hd11[16]), 
        .product_15_(hd11[15]), .product_14_(hd11[14]), .product_13_(hd11[13]), 
        .product_12_(hd11[12]), .product_11_(hd11[11]), .product_10_(hd11[10]), 
        .product_9_(hd11[9]), .product_8_(hd11[8]), .product_7_(hd11[7]), 
        .product_6_(hd11[6]), .product_5_(hd11[5]), .product_4_(hd11[4]), 
        .product_3_(hd11[3]), .product_2_(hd11[2]), .product_1_(hd11[1]) );
  FAS_DW_mult_tc_34 mult_36 ( .a(data), .product({hd05_35, hd05}) );
  FAS_DW_mult_tc_35 mult_34 ( .a(data), .product({hd03_35, hd03}) );
  FAS_DW_mult_tc_36 mult_43 ( .a(data), .product_26_(hd12_35), .product_25_(
        hd12[25]), .product_24_(hd12[24]), .product_23_(hd12[23]), 
        .product_22_(hd12[22]), .product_21_(hd12[21]), .product_20_(hd12[20]), 
        .product_19_(hd12[19]), .product_18_(hd12[18]), .product_17_(hd12[17]), 
        .product_16_(hd12[16]), .product_15_(hd12[15]), .product_14_(hd12[14]), 
        .product_13_(hd12[13]), .product_12_(hd12[12]), .product_11_(hd12[11]), 
        .product_10_(hd12[10]), .product_9_(hd12[9]), .product_8_(hd12[8]), 
        .product_7_(hd12[7]), .product_6_(hd12[6]), .product_5_(hd12[5]), 
        .product_4_(hd12[4]), .product_3_(hd12[3]), .product_2_(hd12[2]) );
  FAS_DW_mult_tc_37 mult_46 ( .a(data), .product_30_(hd15_35), .product_29_(
        hd15[29]), .product_28_(hd15[28]), .product_27_(hd15[27]), 
        .product_26_(hd15[26]), .product_25_(hd15[25]), .product_24_(hd15[24]), 
        .product_23_(hd15[23]), .product_22_(hd15[22]), .product_21_(hd15[21]), 
        .product_20_(hd15[20]), .product_19_(hd15[19]), .product_18_(hd15[18]), 
        .product_17_(hd15[17]), .product_16_(hd15[16]), .product_15_(hd15[15]), 
        .product_14_(hd15[14]), .product_13_(hd15[13]), .product_12_(hd15[12]), 
        .product_11_(hd15[11]), .product_10_(hd15[10]), .product_9_(hd15[9]), 
        .product_8_(hd15[8]), .product_7_(hd15[7]), .product_6_(hd15[6]), 
        .product_5_(hd15[5]), .product_4_(hd15[4]), .product_3_(hd15[3]), 
        .product_2_(hd15[2]), .product_1_(hd15[1]) );
  FAS_DW_mult_tc_38 mult_45 ( .a(data), .product_29_(hd14_35), .product_28_(
        hd14[28]), .product_27_(hd14[27]), .product_26_(hd14[26]), 
        .product_25_(hd14[25]), .product_24_(hd14[24]), .product_23_(hd14[23]), 
        .product_22_(hd14[22]), .product_21_(hd14[21]), .product_20_(hd14[20]), 
        .product_19_(hd14[19]), .product_18_(hd14[18]), .product_17_(hd14[17]), 
        .product_16_(hd14[16]), .product_15_(hd14[15]), .product_14_(hd14[14]), 
        .product_13_(hd14[13]), .product_12_(hd14[12]), .product_11_(hd14[11]), 
        .product_10_(hd14[10]), .product_9_(hd14[9]), .product_8_(hd14[8]), 
        .product_7_(hd14[7]), .product_6_(hd14[6]), .product_5_(hd14[5]), 
        .product_4_(hd14[4]), .product_3_(hd14[3]), .product_2_(hd14[2]) );
  FAS_DW_mult_tc_39 mult_35 ( .a(data), .product({hd04_35, hd04}) );
  FAS_DW_mult_tc_40 mult_47 ( .a(data), .product({hd16_35, hd16}) );
  FAS_DW_mult_tc_41 mult_44 ( .a(data), .product_28_(hd13_35), .product_27_(
        hd13[27]), .product_26_(hd13[26]), .product_25_(hd13[25]), 
        .product_24_(hd13[24]), .product_23_(hd13[23]), .product_22_(hd13[22]), 
        .product_21_(hd13[21]), .product_20_(hd13[20]), .product_19_(hd13[19]), 
        .product_18_(hd13[18]), .product_17_(hd13[17]), .product_16_(hd13[16]), 
        .product_15_(hd13[15]), .product_14_(hd13[14]), .product_13_(hd13[13]), 
        .product_12_(hd13[12]), .product_11_(hd13[11]), .product_10_(hd13[10]), 
        .product_9_(hd13[9]), .product_8_(hd13[8]), .product_7_(hd13[7]), 
        .product_6_(hd13[6]), .product_5_(hd13[5]), .product_4_(hd13[4]), 
        .product_3_(hd13[3]), .product_2_(hd13[2]), .product_1_(hd13[1]) );
  FAS_DW_mult_tc_42 mult_41 ( .a(data), .product_28_(hd10_35), .product_27_(
        hd10[27]), .product_26_(hd10[26]), .product_25_(hd10[25]), 
        .product_24_(hd10[24]), .product_23_(hd10[23]), .product_22_(hd10[22]), 
        .product_21_(hd10[21]), .product_20_(hd10[20]), .product_19_(hd10[19]), 
        .product_18_(hd10[18]), .product_17_(hd10[17]), .product_16_(hd10[16]), 
        .product_15_(hd10[15]), .product_14_(hd10[14]), .product_13_(hd10[13]), 
        .product_12_(hd10[12]), .product_11_(hd10[11]), .product_10_(hd10[10]), 
        .product_9_(hd10[9]), .product_8_(hd10[8]), .product_7_(hd10[7]), 
        .product_6_(hd10[6]), .product_5_(hd10[5]), .product_4_(hd10[4]), 
        .product_3_(hd10[3]), .product_2_(hd10[2]), .product_1_(hd10[1]) );
  CLKMX2X2 U4025 ( .A(1'b0), .B(d02[0]), .S0(n8631), .Y(n5992) );
  OA21XL U4027 ( .A0(n8689), .A1(n6194), .B0(n6190), .Y(n6195) );
  NAND3X2 U4028 ( .A(n8781), .B(n8755), .C(n8792), .Y(n9317) );
  NOR2X2 U4029 ( .A(n6111), .B(n11224), .Y(n9250) );
  NOR2X2 U4030 ( .A(BF2I_b_s), .B(n11223), .Y(n9249) );
  INVX3 U4031 ( .A(mult_add_355_aco_b), .Y(n9245) );
  OA21X2 U4032 ( .A0(n10475), .A1(n9582), .B0(n9617), .Y(n9584) );
  NAND2XL U4033 ( .A(n6193), .B(n9623), .Y(n9617) );
  OAI21X1 U4034 ( .A0(n9380), .A1(n9381), .B0(fir_valid), .Y(n9315) );
  NOR2XL U4035 ( .A(n9245), .B(n9198), .Y(N1363) );
  AOI22XL U4036 ( .A0(N446), .A1(n9383), .B0(N542), .B1(n9384), .Y(n9419) );
  AOI22XL U4037 ( .A0(N445), .A1(n9383), .B0(N541), .B1(n9384), .Y(n9417) );
  AOI22XL U4038 ( .A0(N444), .A1(n9383), .B0(N540), .B1(n9384), .Y(n9415) );
  AOI22XL U4039 ( .A0(N443), .A1(n9383), .B0(N539), .B1(n9384), .Y(n9413) );
  AOI22XL U4040 ( .A0(N442), .A1(n9383), .B0(N538), .B1(n9384), .Y(n9411) );
  AOI22XL U4041 ( .A0(N441), .A1(n9383), .B0(N537), .B1(n9384), .Y(n9409) );
  AOI22XL U4042 ( .A0(N440), .A1(n9383), .B0(N536), .B1(n9384), .Y(n9407) );
  AOI22XL U4043 ( .A0(N439), .A1(n9383), .B0(N535), .B1(n9384), .Y(n9405) );
  AOI22XL U4044 ( .A0(N438), .A1(n9383), .B0(N534), .B1(n9384), .Y(n9403) );
  AOI22XL U4045 ( .A0(N437), .A1(n9383), .B0(N533), .B1(n9384), .Y(n9401) );
  AOI22XL U4046 ( .A0(N436), .A1(n9383), .B0(N532), .B1(n9384), .Y(n9399) );
  AOI22XL U4047 ( .A0(N435), .A1(n9383), .B0(N531), .B1(n9384), .Y(n9397) );
  AOI22XL U4048 ( .A0(N434), .A1(n9383), .B0(N530), .B1(n9384), .Y(n9395) );
  AOI22XL U4049 ( .A0(N433), .A1(n9383), .B0(N529), .B1(n9384), .Y(n9393) );
  AOI22XL U4050 ( .A0(n9468), .A1(N452), .B0(N388), .B1(n9469), .Y(n9496) );
  AOI22XL U4051 ( .A0(n9468), .A1(N453), .B0(N389), .B1(n9469), .Y(n9495) );
  AOI22XL U4052 ( .A0(n9468), .A1(N454), .B0(N390), .B1(n9469), .Y(n9494) );
  AOI22XL U4053 ( .A0(n9468), .A1(N455), .B0(N391), .B1(n9469), .Y(n9493) );
  AOI22XL U4054 ( .A0(n9468), .A1(N456), .B0(N392), .B1(n9469), .Y(n9492) );
  AOI22XL U4055 ( .A0(n9468), .A1(N457), .B0(N393), .B1(n9469), .Y(n9491) );
  AOI22XL U4056 ( .A0(n9468), .A1(N458), .B0(N394), .B1(n9469), .Y(n9490) );
  AOI22XL U4057 ( .A0(n9468), .A1(N459), .B0(N395), .B1(n9469), .Y(n9489) );
  AOI22XL U4058 ( .A0(n9468), .A1(N460), .B0(N396), .B1(n9469), .Y(n9488) );
  AOI22XL U4059 ( .A0(n9468), .A1(N461), .B0(N397), .B1(n9469), .Y(n9487) );
  AOI22XL U4060 ( .A0(n9468), .A1(N462), .B0(N398), .B1(n9469), .Y(n9486) );
  AOI22XL U4061 ( .A0(n9468), .A1(N463), .B0(n9469), .B1(N399), .Y(n9485) );
  AOI22XL U4062 ( .A0(N384), .A1(n9468), .B0(n9469), .B1(N368), .Y(n9484) );
  AOI22XL U4063 ( .A0(N385), .A1(n9468), .B0(n9469), .B1(N369), .Y(n9483) );
  AOI22XL U4064 ( .A0(N386), .A1(n9468), .B0(n9469), .B1(N370), .Y(n9482) );
  AOI22XL U4065 ( .A0(N387), .A1(n9468), .B0(n9469), .B1(N371), .Y(n9481) );
  AOI22XL U4066 ( .A0(N388), .A1(n9468), .B0(n9469), .B1(N372), .Y(n9480) );
  AOI22XL U4067 ( .A0(N389), .A1(n9468), .B0(n9469), .B1(N373), .Y(n9479) );
  AOI22XL U4068 ( .A0(N390), .A1(n9468), .B0(n9469), .B1(N374), .Y(n9478) );
  AOI22XL U4069 ( .A0(N391), .A1(n9468), .B0(n9469), .B1(N375), .Y(n9477) );
  AOI22XL U4070 ( .A0(N392), .A1(n9468), .B0(n9469), .B1(N376), .Y(n9476) );
  AOI22XL U4071 ( .A0(N393), .A1(n9468), .B0(n9469), .B1(N377), .Y(n9475) );
  AOI22XL U4072 ( .A0(N394), .A1(n9468), .B0(n9469), .B1(N378), .Y(n9474) );
  AOI22XL U4073 ( .A0(N395), .A1(n9468), .B0(n9469), .B1(N379), .Y(n9473) );
  AOI22XL U4074 ( .A0(N396), .A1(n9468), .B0(n9469), .B1(N380), .Y(n9472) );
  AOI22XL U4075 ( .A0(N397), .A1(n9468), .B0(n9469), .B1(N381), .Y(n9471) );
  AOI22XL U4076 ( .A0(N398), .A1(n9468), .B0(n9469), .B1(N382), .Y(n9470) );
  AOI22XL U4077 ( .A0(N399), .A1(n9468), .B0(n9469), .B1(N383), .Y(n9467) );
  CLKBUFX3 U4078 ( .A(n8891), .Y(n8886) );
  CLKBUFX3 U4079 ( .A(n8891), .Y(n8887) );
  CLKBUFX3 U4080 ( .A(n8890), .Y(n8888) );
  CLKBUFX3 U4081 ( .A(n8892), .Y(n8884) );
  CLKBUFX3 U4082 ( .A(n8892), .Y(n8885) );
  CLKBUFX3 U4083 ( .A(n8894), .Y(n8881) );
  CLKBUFX3 U4084 ( .A(n8893), .Y(n8882) );
  CLKBUFX3 U4085 ( .A(n8893), .Y(n8883) );
  CLKBUFX3 U4086 ( .A(n8895), .Y(n8879) );
  CLKBUFX3 U4087 ( .A(n8894), .Y(n8880) );
  CLKBUFX3 U4088 ( .A(n8896), .Y(n8876) );
  CLKBUFX3 U4089 ( .A(n8896), .Y(n8877) );
  CLKBUFX3 U4090 ( .A(n8895), .Y(n8878) );
  CLKBUFX3 U4091 ( .A(n8897), .Y(n8874) );
  CLKBUFX3 U4092 ( .A(n8897), .Y(n8875) );
  CLKBUFX3 U4093 ( .A(n8899), .Y(n8871) );
  CLKBUFX3 U4094 ( .A(n8898), .Y(n8872) );
  CLKBUFX3 U4095 ( .A(n8898), .Y(n8873) );
  CLKBUFX3 U4096 ( .A(n8900), .Y(n8869) );
  CLKBUFX3 U4097 ( .A(n8899), .Y(n8870) );
  CLKBUFX3 U4098 ( .A(n8901), .Y(n8867) );
  CLKBUFX3 U4099 ( .A(n8900), .Y(n8868) );
  CLKBUFX3 U4100 ( .A(n8902), .Y(n8864) );
  CLKBUFX3 U4101 ( .A(n8902), .Y(n8865) );
  CLKBUFX3 U4102 ( .A(n8901), .Y(n8866) );
  CLKBUFX3 U4103 ( .A(n8903), .Y(n8862) );
  CLKBUFX3 U4104 ( .A(n8903), .Y(n8863) );
  CLKBUFX3 U4105 ( .A(n8905), .Y(n8859) );
  CLKBUFX3 U4106 ( .A(n8904), .Y(n8860) );
  CLKBUFX3 U4107 ( .A(n8904), .Y(n8861) );
  CLKBUFX3 U4108 ( .A(n8906), .Y(n8857) );
  CLKBUFX3 U4109 ( .A(n8905), .Y(n8858) );
  CLKBUFX3 U4110 ( .A(n8907), .Y(n8854) );
  CLKBUFX3 U4111 ( .A(n8907), .Y(n8855) );
  CLKBUFX3 U4112 ( .A(n8906), .Y(n8856) );
  CLKBUFX3 U4113 ( .A(n8890), .Y(n8889) );
  CLKBUFX3 U4114 ( .A(n9143), .Y(n8937) );
  CLKBUFX3 U4115 ( .A(n9143), .Y(n8936) );
  CLKBUFX3 U4116 ( .A(n9137), .Y(n9015) );
  CLKBUFX3 U4117 ( .A(n9139), .Y(n8994) );
  CLKBUFX3 U4118 ( .A(n9142), .Y(n8956) );
  CLKBUFX3 U4119 ( .A(n9141), .Y(n8961) );
  CLKBUFX3 U4120 ( .A(n9141), .Y(n8966) );
  CLKBUFX3 U4121 ( .A(n9141), .Y(n8971) );
  CLKBUFX3 U4122 ( .A(n9137), .Y(n9012) );
  CLKBUFX3 U4123 ( .A(n9138), .Y(n9007) );
  CLKBUFX3 U4124 ( .A(n9143), .Y(n8939) );
  CLKBUFX3 U4125 ( .A(n9140), .Y(n8976) );
  CLKBUFX3 U4126 ( .A(n9143), .Y(n8944) );
  CLKBUFX3 U4127 ( .A(n9139), .Y(n8989) );
  CLKBUFX3 U4128 ( .A(n9140), .Y(n8981) );
  CLKBUFX3 U4129 ( .A(n9142), .Y(n8949) );
  CLKBUFX3 U4130 ( .A(n9138), .Y(n9010) );
  CLKBUFX3 U4131 ( .A(n9138), .Y(n9002) );
  CLKBUFX3 U4132 ( .A(n9142), .Y(n8954) );
  CLKBUFX3 U4133 ( .A(n9142), .Y(n8959) );
  CLKBUFX3 U4134 ( .A(n9141), .Y(n8964) );
  CLKBUFX3 U4135 ( .A(n9138), .Y(n9005) );
  CLKBUFX3 U4136 ( .A(n9139), .Y(n8997) );
  CLKBUFX3 U4137 ( .A(n9141), .Y(n8969) );
  CLKBUFX3 U4138 ( .A(n9143), .Y(n8934) );
  CLKBUFX3 U4139 ( .A(n9143), .Y(n8942) );
  CLKBUFX3 U4140 ( .A(n9137), .Y(n9018) );
  CLKBUFX3 U4141 ( .A(n9140), .Y(n8974) );
  CLKBUFX3 U4142 ( .A(n9142), .Y(n8947) );
  CLKBUFX3 U4143 ( .A(n9140), .Y(n8979) );
  CLKBUFX3 U4144 ( .A(n9138), .Y(n9000) );
  CLKBUFX3 U4145 ( .A(n9142), .Y(n8952) );
  CLKBUFX3 U4146 ( .A(n9139), .Y(n8992) );
  CLKBUFX3 U4147 ( .A(n9140), .Y(n8984) );
  CLKBUFX3 U4148 ( .A(n9142), .Y(n8957) );
  CLKBUFX3 U4149 ( .A(n9137), .Y(n9013) );
  CLKBUFX3 U4150 ( .A(n9141), .Y(n8962) );
  CLKBUFX3 U4151 ( .A(n9139), .Y(n8995) );
  CLKBUFX3 U4152 ( .A(n9141), .Y(n8967) );
  CLKBUFX3 U4153 ( .A(n9137), .Y(n9016) );
  CLKBUFX3 U4154 ( .A(n9141), .Y(n8972) );
  CLKBUFX3 U4155 ( .A(n9138), .Y(n9008) );
  CLKBUFX3 U4156 ( .A(n9143), .Y(n8940) );
  CLKBUFX3 U4157 ( .A(n9140), .Y(n8977) );
  CLKBUFX3 U4158 ( .A(n9143), .Y(n8945) );
  CLKBUFX3 U4159 ( .A(n9139), .Y(n8990) );
  CLKBUFX3 U4160 ( .A(n9143), .Y(n8935) );
  CLKBUFX3 U4161 ( .A(n9140), .Y(n8982) );
  CLKBUFX3 U4162 ( .A(n9142), .Y(n8950) );
  CLKBUFX3 U4163 ( .A(n9137), .Y(n9017) );
  CLKBUFX3 U4164 ( .A(n9138), .Y(n9011) );
  CLKBUFX3 U4165 ( .A(n9138), .Y(n9006) );
  CLKBUFX3 U4166 ( .A(n9138), .Y(n9001) );
  CLKBUFX3 U4167 ( .A(n9139), .Y(n8996) );
  CLKBUFX3 U4168 ( .A(n9139), .Y(n8991) );
  CLKBUFX3 U4169 ( .A(n9143), .Y(n8938) );
  CLKBUFX3 U4170 ( .A(n9143), .Y(n8943) );
  CLKBUFX3 U4171 ( .A(n9142), .Y(n8948) );
  CLKBUFX3 U4172 ( .A(n9142), .Y(n8953) );
  CLKBUFX3 U4173 ( .A(n9142), .Y(n8958) );
  CLKBUFX3 U4174 ( .A(n9141), .Y(n8963) );
  CLKBUFX3 U4175 ( .A(n9141), .Y(n8968) );
  CLKBUFX3 U4176 ( .A(n9140), .Y(n8973) );
  CLKBUFX3 U4177 ( .A(n9140), .Y(n8978) );
  CLKBUFX3 U4178 ( .A(n9140), .Y(n8983) );
  CLKBUFX3 U4179 ( .A(n9138), .Y(n9003) );
  CLKBUFX3 U4180 ( .A(n9143), .Y(n8941) );
  CLKBUFX3 U4181 ( .A(n9143), .Y(n8946) );
  CLKBUFX3 U4182 ( .A(n9142), .Y(n8951) );
  CLKBUFX3 U4183 ( .A(n9142), .Y(n8955) );
  CLKBUFX3 U4184 ( .A(n9141), .Y(n8960) );
  CLKBUFX3 U4185 ( .A(n9141), .Y(n8965) );
  CLKBUFX3 U4186 ( .A(n9141), .Y(n8970) );
  CLKBUFX3 U4187 ( .A(n9140), .Y(n8975) );
  CLKBUFX3 U4188 ( .A(n9140), .Y(n8980) );
  CLKBUFX3 U4189 ( .A(n9140), .Y(n8985) );
  CLKBUFX3 U4190 ( .A(n9139), .Y(n8986) );
  CLKBUFX3 U4191 ( .A(n9137), .Y(n9021) );
  CLKBUFX3 U4192 ( .A(n9139), .Y(n8988) );
  CLKBUFX3 U4193 ( .A(n9139), .Y(n8987) );
  CLKBUFX3 U4194 ( .A(n9139), .Y(n8993) );
  CLKBUFX3 U4195 ( .A(n9139), .Y(n8998) );
  CLKBUFX3 U4196 ( .A(n9138), .Y(n8999) );
  CLKBUFX3 U4197 ( .A(n9138), .Y(n9004) );
  CLKBUFX3 U4198 ( .A(n9138), .Y(n9009) );
  CLKBUFX3 U4199 ( .A(n9137), .Y(n9014) );
  CLKBUFX3 U4200 ( .A(n9137), .Y(n9019) );
  CLKBUFX3 U4201 ( .A(n9137), .Y(n9020) );
  CLKBUFX3 U4202 ( .A(n9137), .Y(n9022) );
  CLKBUFX3 U4203 ( .A(n9136), .Y(n9031) );
  CLKBUFX3 U4204 ( .A(n9136), .Y(n9036) );
  CLKBUFX3 U4205 ( .A(n9137), .Y(n9023) );
  CLKBUFX3 U4206 ( .A(n9137), .Y(n9024) );
  CLKBUFX3 U4207 ( .A(n9136), .Y(n9025) );
  CLKBUFX3 U4208 ( .A(n9136), .Y(n9026) );
  CLKBUFX3 U4209 ( .A(n9136), .Y(n9027) );
  CLKBUFX3 U4210 ( .A(n9136), .Y(n9028) );
  CLKBUFX3 U4211 ( .A(n9136), .Y(n9029) );
  CLKBUFX3 U4212 ( .A(n9136), .Y(n9030) );
  CLKBUFX3 U4213 ( .A(n9136), .Y(n9032) );
  CLKBUFX3 U4214 ( .A(n9136), .Y(n9033) );
  CLKBUFX3 U4215 ( .A(n9136), .Y(n9034) );
  CLKBUFX3 U4216 ( .A(n9136), .Y(n9035) );
  CLKBUFX3 U4217 ( .A(n9136), .Y(n9037) );
  CLKBUFX3 U4218 ( .A(n9135), .Y(n9038) );
  CLKBUFX3 U4219 ( .A(n9135), .Y(n9039) );
  CLKBUFX3 U4220 ( .A(n9135), .Y(n9040) );
  CLKBUFX3 U4221 ( .A(n9135), .Y(n9041) );
  CLKBUFX3 U4222 ( .A(n9135), .Y(n9042) );
  CLKBUFX3 U4223 ( .A(n9135), .Y(n9043) );
  CLKBUFX3 U4224 ( .A(n9135), .Y(n9044) );
  CLKBUFX3 U4225 ( .A(n9135), .Y(n9045) );
  CLKBUFX3 U4226 ( .A(n9135), .Y(n9046) );
  CLKBUFX3 U4227 ( .A(n9135), .Y(n9047) );
  CLKBUFX3 U4228 ( .A(n9135), .Y(n9048) );
  CLKBUFX3 U4229 ( .A(n9129), .Y(n9127) );
  CLKBUFX3 U4230 ( .A(n9135), .Y(n9049) );
  CLKBUFX3 U4231 ( .A(n9132), .Y(n9084) );
  CLKBUFX3 U4232 ( .A(n9134), .Y(n9052) );
  CLKBUFX3 U4233 ( .A(n9130), .Y(n9108) );
  CLKBUFX3 U4234 ( .A(n9134), .Y(n9057) );
  CLKBUFX3 U4235 ( .A(n9129), .Y(n9120) );
  CLKBUFX3 U4236 ( .A(n9132), .Y(n9089) );
  CLKBUFX3 U4237 ( .A(n9134), .Y(n9062) );
  CLKBUFX3 U4238 ( .A(n9144), .Y(n8924) );
  CLKBUFX3 U4239 ( .A(n9131), .Y(n9101) );
  CLKBUFX3 U4240 ( .A(n9133), .Y(n9067) );
  CLKBUFX3 U4241 ( .A(n9144), .Y(n8931) );
  CLKBUFX3 U4242 ( .A(n9130), .Y(n9113) );
  CLKBUFX3 U4243 ( .A(n9133), .Y(n9072) );
  CLKBUFX3 U4244 ( .A(n9129), .Y(n9125) );
  CLKBUFX3 U4245 ( .A(n9131), .Y(n9094) );
  CLKBUFX3 U4246 ( .A(n9132), .Y(n9077) );
  CLKBUFX3 U4247 ( .A(n9130), .Y(n9106) );
  CLKBUFX3 U4248 ( .A(n9132), .Y(n9082) );
  CLKBUFX3 U4249 ( .A(n9135), .Y(n9050) );
  CLKBUFX3 U4250 ( .A(n9129), .Y(n9118) );
  CLKBUFX3 U4251 ( .A(n9132), .Y(n9087) );
  CLKBUFX3 U4252 ( .A(n9134), .Y(n9055) );
  CLKBUFX3 U4253 ( .A(n9144), .Y(n8929) );
  CLKBUFX3 U4254 ( .A(n9131), .Y(n9099) );
  CLKBUFX3 U4255 ( .A(n9134), .Y(n9060) );
  CLKBUFX3 U4256 ( .A(n9130), .Y(n9111) );
  CLKBUFX3 U4257 ( .A(n9133), .Y(n9065) );
  CLKBUFX3 U4258 ( .A(n9129), .Y(n9123) );
  CLKBUFX3 U4259 ( .A(n9131), .Y(n9092) );
  CLKBUFX3 U4260 ( .A(n9133), .Y(n9070) );
  CLKBUFX3 U4261 ( .A(n9130), .Y(n9104) );
  CLKBUFX3 U4262 ( .A(n9133), .Y(n9075) );
  CLKBUFX3 U4263 ( .A(n9144), .Y(n8927) );
  CLKBUFX3 U4264 ( .A(n9129), .Y(n9116) );
  CLKBUFX3 U4265 ( .A(n9132), .Y(n9080) );
  CLKBUFX3 U4266 ( .A(n9131), .Y(n9097) );
  CLKBUFX3 U4267 ( .A(n9132), .Y(n9085) );
  CLKBUFX3 U4268 ( .A(n9134), .Y(n9053) );
  CLKBUFX3 U4269 ( .A(n9130), .Y(n9109) );
  CLKBUFX3 U4270 ( .A(n9134), .Y(n9058) );
  CLKBUFX3 U4271 ( .A(n9129), .Y(n9121) );
  CLKBUFX3 U4272 ( .A(n9131), .Y(n9090) );
  CLKBUFX3 U4273 ( .A(n9134), .Y(n9063) );
  CLKBUFX3 U4274 ( .A(n9144), .Y(n8925) );
  CLKBUFX3 U4275 ( .A(n9131), .Y(n9102) );
  CLKBUFX3 U4276 ( .A(n9133), .Y(n9068) );
  CLKBUFX3 U4277 ( .A(n9144), .Y(n8932) );
  CLKBUFX3 U4278 ( .A(n9130), .Y(n9114) );
  CLKBUFX3 U4279 ( .A(n9133), .Y(n9073) );
  CLKBUFX3 U4280 ( .A(n9129), .Y(n9126) );
  CLKBUFX3 U4281 ( .A(n9131), .Y(n9095) );
  CLKBUFX3 U4282 ( .A(n9132), .Y(n9078) );
  CLKBUFX3 U4283 ( .A(n9129), .Y(n9124) );
  CLKBUFX3 U4284 ( .A(n9129), .Y(n9122) );
  CLKBUFX3 U4285 ( .A(n9129), .Y(n9119) );
  CLKBUFX3 U4286 ( .A(n9129), .Y(n9117) );
  CLKBUFX3 U4287 ( .A(n9130), .Y(n9115) );
  CLKBUFX3 U4288 ( .A(n9130), .Y(n9112) );
  CLKBUFX3 U4289 ( .A(n9130), .Y(n9110) );
  CLKBUFX3 U4290 ( .A(n9130), .Y(n9107) );
  CLKBUFX3 U4291 ( .A(n9130), .Y(n9105) );
  CLKBUFX3 U4292 ( .A(n9130), .Y(n9103) );
  CLKBUFX3 U4293 ( .A(n9131), .Y(n9100) );
  CLKBUFX3 U4294 ( .A(n9131), .Y(n9098) );
  CLKBUFX3 U4295 ( .A(n9131), .Y(n9096) );
  CLKBUFX3 U4296 ( .A(n9131), .Y(n9093) );
  CLKBUFX3 U4297 ( .A(n9131), .Y(n9091) );
  CLKBUFX3 U4298 ( .A(n9132), .Y(n9088) );
  CLKBUFX3 U4299 ( .A(n9132), .Y(n9086) );
  CLKBUFX3 U4300 ( .A(n9132), .Y(n9083) );
  CLKBUFX3 U4301 ( .A(n9132), .Y(n9081) );
  CLKBUFX3 U4302 ( .A(n9132), .Y(n9079) );
  CLKBUFX3 U4303 ( .A(n9133), .Y(n9076) );
  CLKBUFX3 U4304 ( .A(n9133), .Y(n9074) );
  CLKBUFX3 U4305 ( .A(n9133), .Y(n9071) );
  CLKBUFX3 U4306 ( .A(n9133), .Y(n9069) );
  CLKBUFX3 U4307 ( .A(n9133), .Y(n9066) );
  CLKBUFX3 U4308 ( .A(n9133), .Y(n9064) );
  CLKBUFX3 U4309 ( .A(n9134), .Y(n9061) );
  CLKBUFX3 U4310 ( .A(n9134), .Y(n9059) );
  CLKBUFX3 U4311 ( .A(n9134), .Y(n9056) );
  CLKBUFX3 U4312 ( .A(n9134), .Y(n9054) );
  CLKBUFX3 U4313 ( .A(n9134), .Y(n9051) );
  CLKBUFX3 U4314 ( .A(n9144), .Y(n8933) );
  CLKBUFX3 U4315 ( .A(n9144), .Y(n8930) );
  CLKBUFX3 U4316 ( .A(n9144), .Y(n8928) );
  CLKBUFX3 U4317 ( .A(n9144), .Y(n8926) );
  CLKBUFX3 U4318 ( .A(n9129), .Y(n9128) );
  CLKINVX1 U4319 ( .A(n8840), .Y(n8828) );
  CLKINVX1 U4320 ( .A(n8840), .Y(n8829) );
  CLKINVX1 U4321 ( .A(n8840), .Y(n8830) );
  CLKINVX1 U4322 ( .A(n8840), .Y(n8831) );
  CLKINVX1 U4323 ( .A(n8840), .Y(n8832) );
  CLKINVX1 U4324 ( .A(n8840), .Y(n8833) );
  CLKINVX1 U4325 ( .A(n8844), .Y(n8805) );
  CLKINVX1 U4326 ( .A(n8844), .Y(n8806) );
  CLKINVX1 U4327 ( .A(n8844), .Y(n8807) );
  CLKINVX1 U4328 ( .A(n8844), .Y(n8808) );
  CLKINVX1 U4329 ( .A(n8844), .Y(n8809) );
  CLKINVX1 U4330 ( .A(n8843), .Y(n8810) );
  CLKINVX1 U4331 ( .A(n8843), .Y(n8811) );
  CLKINVX1 U4332 ( .A(n8843), .Y(n8812) );
  CLKINVX1 U4333 ( .A(n8843), .Y(n8813) );
  CLKINVX1 U4334 ( .A(n8843), .Y(n8814) );
  CLKINVX1 U4335 ( .A(n8843), .Y(n8815) );
  CLKINVX1 U4336 ( .A(n8842), .Y(n8816) );
  CLKINVX1 U4337 ( .A(n8842), .Y(n8817) );
  CLKINVX1 U4338 ( .A(n8842), .Y(n8818) );
  CLKINVX1 U4339 ( .A(n8842), .Y(n8819) );
  CLKINVX1 U4340 ( .A(n8842), .Y(n8820) );
  CLKINVX1 U4341 ( .A(n8842), .Y(n8821) );
  CLKINVX1 U4342 ( .A(n8841), .Y(n8822) );
  CLKINVX1 U4343 ( .A(n8841), .Y(n8823) );
  CLKINVX1 U4344 ( .A(n8841), .Y(n8824) );
  CLKINVX1 U4345 ( .A(n8841), .Y(n8825) );
  CLKINVX1 U4346 ( .A(n8841), .Y(n8826) );
  CLKINVX1 U4347 ( .A(n8841), .Y(n8827) );
  CLKINVX1 U4348 ( .A(n8845), .Y(n8803) );
  CLKINVX1 U4349 ( .A(n8845), .Y(n8804) );
  CLKBUFX3 U4350 ( .A(n8701), .Y(n8658) );
  CLKBUFX3 U4351 ( .A(n8701), .Y(n8659) );
  CLKBUFX3 U4352 ( .A(n8701), .Y(n8660) );
  CLKBUFX3 U4353 ( .A(n8700), .Y(n8661) );
  CLKBUFX3 U4354 ( .A(n8700), .Y(n8662) );
  CLKBUFX3 U4355 ( .A(n8700), .Y(n8663) );
  CLKBUFX3 U4356 ( .A(n8699), .Y(n8664) );
  CLKBUFX3 U4357 ( .A(n8699), .Y(n8665) );
  CLKBUFX3 U4358 ( .A(n8699), .Y(n8666) );
  CLKBUFX3 U4359 ( .A(n8698), .Y(n8667) );
  CLKBUFX3 U4360 ( .A(n8705), .Y(n8647) );
  CLKBUFX3 U4361 ( .A(n8705), .Y(n8648) );
  CLKBUFX3 U4362 ( .A(n8704), .Y(n8649) );
  CLKBUFX3 U4363 ( .A(n8704), .Y(n8650) );
  CLKBUFX3 U4364 ( .A(n8704), .Y(n8651) );
  CLKBUFX3 U4365 ( .A(n8703), .Y(n8652) );
  CLKBUFX3 U4366 ( .A(n8703), .Y(n8653) );
  CLKBUFX3 U4367 ( .A(n8703), .Y(n8654) );
  CLKBUFX3 U4368 ( .A(n8702), .Y(n8655) );
  CLKBUFX3 U4369 ( .A(n8702), .Y(n8656) );
  CLKBUFX3 U4370 ( .A(n8702), .Y(n8657) );
  CLKBUFX3 U4371 ( .A(n8694), .Y(n8680) );
  CLKBUFX3 U4372 ( .A(n8694), .Y(n8681) );
  CLKBUFX3 U4373 ( .A(n8693), .Y(n8682) );
  CLKBUFX3 U4374 ( .A(n8693), .Y(n8683) );
  CLKBUFX3 U4375 ( .A(n8693), .Y(n8684) );
  CLKBUFX3 U4376 ( .A(n8692), .Y(n8685) );
  CLKBUFX3 U4377 ( .A(n8692), .Y(n8686) );
  CLKBUFX3 U4378 ( .A(n8692), .Y(n8687) );
  CLKBUFX3 U4379 ( .A(n8691), .Y(n8688) );
  CLKBUFX3 U4380 ( .A(n8698), .Y(n8668) );
  CLKBUFX3 U4381 ( .A(n8698), .Y(n8669) );
  CLKBUFX3 U4382 ( .A(n8697), .Y(n8670) );
  CLKBUFX3 U4383 ( .A(n8697), .Y(n8671) );
  CLKBUFX3 U4384 ( .A(n8697), .Y(n8672) );
  CLKBUFX3 U4385 ( .A(n8696), .Y(n8673) );
  CLKBUFX3 U4386 ( .A(n8696), .Y(n8674) );
  CLKBUFX3 U4387 ( .A(n8696), .Y(n8675) );
  CLKBUFX3 U4388 ( .A(n8695), .Y(n8676) );
  CLKBUFX3 U4389 ( .A(n8695), .Y(n8677) );
  CLKBUFX3 U4390 ( .A(n8695), .Y(n8678) );
  CLKBUFX3 U4391 ( .A(n8694), .Y(n8679) );
  CLKBUFX3 U4392 ( .A(n8716), .Y(n8615) );
  CLKBUFX3 U4393 ( .A(n8715), .Y(n8616) );
  CLKBUFX3 U4394 ( .A(n8715), .Y(n8617) );
  CLKBUFX3 U4395 ( .A(n8715), .Y(n8618) );
  CLKBUFX3 U4396 ( .A(n8714), .Y(n8619) );
  CLKBUFX3 U4397 ( .A(n8714), .Y(n8620) );
  CLKBUFX3 U4398 ( .A(n8714), .Y(n8621) );
  CLKBUFX3 U4399 ( .A(n8713), .Y(n8622) );
  CLKBUFX3 U4400 ( .A(n8713), .Y(n8623) );
  CLKBUFX3 U4401 ( .A(n8713), .Y(n8624) );
  CLKBUFX3 U4402 ( .A(n8719), .Y(n8605) );
  CLKBUFX3 U4403 ( .A(n8719), .Y(n8606) );
  CLKBUFX3 U4404 ( .A(n8718), .Y(n8607) );
  CLKBUFX3 U4405 ( .A(n8718), .Y(n8608) );
  CLKBUFX3 U4406 ( .A(n8718), .Y(n8609) );
  CLKBUFX3 U4407 ( .A(n8717), .Y(n8610) );
  CLKBUFX3 U4408 ( .A(n8717), .Y(n8611) );
  CLKBUFX3 U4409 ( .A(n8717), .Y(n8612) );
  CLKBUFX3 U4410 ( .A(n8716), .Y(n8613) );
  CLKBUFX3 U4411 ( .A(n8716), .Y(n8614) );
  CLKBUFX3 U4412 ( .A(n8708), .Y(n8637) );
  CLKBUFX3 U4413 ( .A(n8708), .Y(n8638) );
  CLKBUFX3 U4414 ( .A(n8708), .Y(n8639) );
  CLKBUFX3 U4415 ( .A(n8707), .Y(n8640) );
  CLKBUFX3 U4416 ( .A(n8707), .Y(n8641) );
  CLKBUFX3 U4417 ( .A(n8707), .Y(n8642) );
  CLKBUFX3 U4418 ( .A(n8706), .Y(n8643) );
  CLKBUFX3 U4419 ( .A(n8706), .Y(n8644) );
  CLKBUFX3 U4420 ( .A(n8706), .Y(n8645) );
  CLKBUFX3 U4421 ( .A(n8705), .Y(n8646) );
  CLKBUFX3 U4422 ( .A(n8712), .Y(n8625) );
  CLKBUFX3 U4423 ( .A(n8712), .Y(n8626) );
  CLKBUFX3 U4424 ( .A(n8712), .Y(n8627) );
  CLKBUFX3 U4425 ( .A(n8711), .Y(n8628) );
  CLKBUFX3 U4426 ( .A(n8711), .Y(n8629) );
  CLKBUFX3 U4427 ( .A(n8711), .Y(n8630) );
  CLKBUFX3 U4428 ( .A(n8710), .Y(n8631) );
  CLKBUFX3 U4429 ( .A(n8710), .Y(n8632) );
  CLKBUFX3 U4430 ( .A(n8710), .Y(n8633) );
  CLKBUFX3 U4431 ( .A(n8709), .Y(n8634) );
  CLKBUFX3 U4432 ( .A(n8709), .Y(n8635) );
  CLKBUFX3 U4433 ( .A(n8709), .Y(n8636) );
  CLKBUFX3 U4434 ( .A(n8719), .Y(n8604) );
  CLKBUFX3 U4435 ( .A(n8691), .Y(n8689) );
  CLKBUFX3 U4436 ( .A(n8763), .Y(n8751) );
  CLKBUFX3 U4437 ( .A(n8763), .Y(n8752) );
  CLKBUFX3 U4438 ( .A(n8762), .Y(n8753) );
  CLKBUFX3 U4439 ( .A(n8762), .Y(n8754) );
  CLKBUFX3 U4440 ( .A(n8767), .Y(n8744) );
  CLKBUFX3 U4441 ( .A(n8767), .Y(n8743) );
  CLKBUFX3 U4442 ( .A(n8768), .Y(n8742) );
  CLKBUFX3 U4443 ( .A(n8768), .Y(n8741) );
  CLKBUFX3 U4444 ( .A(n8769), .Y(n8740) );
  CLKBUFX3 U4445 ( .A(n8769), .Y(n8739) );
  CLKBUFX3 U4446 ( .A(n8764), .Y(n8749) );
  CLKBUFX3 U4447 ( .A(n8765), .Y(n8748) );
  CLKBUFX3 U4448 ( .A(n8765), .Y(n8747) );
  CLKBUFX3 U4449 ( .A(n8766), .Y(n8746) );
  CLKBUFX3 U4450 ( .A(n8766), .Y(n8745) );
  CLKBUFX3 U4451 ( .A(n8764), .Y(n8750) );
  CLKBUFX3 U4452 ( .A(n8919), .Y(n8891) );
  CLKBUFX3 U4453 ( .A(n8919), .Y(n8890) );
  CLKBUFX3 U4454 ( .A(n8918), .Y(n8892) );
  CLKBUFX3 U4455 ( .A(n8918), .Y(n8893) );
  CLKBUFX3 U4456 ( .A(n8917), .Y(n8894) );
  CLKBUFX3 U4457 ( .A(n8916), .Y(n8896) );
  CLKBUFX3 U4458 ( .A(n8917), .Y(n8895) );
  CLKBUFX3 U4459 ( .A(n8916), .Y(n8897) );
  CLKBUFX3 U4460 ( .A(n8915), .Y(n8898) );
  CLKBUFX3 U4461 ( .A(n8915), .Y(n8899) );
  CLKBUFX3 U4462 ( .A(n8914), .Y(n8900) );
  CLKBUFX3 U4463 ( .A(n8913), .Y(n8902) );
  CLKBUFX3 U4464 ( .A(n8914), .Y(n8901) );
  CLKBUFX3 U4465 ( .A(n8913), .Y(n8903) );
  CLKBUFX3 U4466 ( .A(n8912), .Y(n8904) );
  CLKBUFX3 U4467 ( .A(n8912), .Y(n8905) );
  CLKBUFX3 U4468 ( .A(n8911), .Y(n8907) );
  CLKBUFX3 U4469 ( .A(n8911), .Y(n8906) );
  CLKBUFX3 U4470 ( .A(n8761), .Y(n8755) );
  CLKBUFX3 U4471 ( .A(n8761), .Y(n8756) );
  CLKBUFX3 U4472 ( .A(n8760), .Y(n8758) );
  CLKBUFX3 U4473 ( .A(n8760), .Y(n8757) );
  CLKBUFX3 U4474 ( .A(n8909), .Y(n8850) );
  CLKBUFX3 U4475 ( .A(n8909), .Y(n8851) );
  CLKBUFX3 U4476 ( .A(n8908), .Y(n8852) );
  CLKBUFX3 U4477 ( .A(n8908), .Y(n8853) );
  CLKBUFX3 U4478 ( .A(n8691), .Y(n8690) );
  CLKINVX1 U4479 ( .A(n8839), .Y(n8834) );
  CLKINVX1 U4480 ( .A(n8839), .Y(n8835) );
  CLKINVX1 U4481 ( .A(n8839), .Y(n8836) );
  CLKINVX1 U4482 ( .A(n8839), .Y(n8837) );
  CLKINVX1 U4483 ( .A(n8839), .Y(n8838) );
  CLKBUFX3 U4484 ( .A(n8848), .Y(n8840) );
  CLKBUFX3 U4485 ( .A(n8846), .Y(n8844) );
  CLKBUFX3 U4486 ( .A(n8847), .Y(n8843) );
  CLKBUFX3 U4487 ( .A(n8847), .Y(n8842) );
  CLKBUFX3 U4488 ( .A(n8848), .Y(n8841) );
  CLKBUFX3 U4489 ( .A(n8920), .Y(n8919) );
  CLKBUFX3 U4490 ( .A(n8920), .Y(n8918) );
  CLKBUFX3 U4491 ( .A(n8920), .Y(n8917) );
  CLKBUFX3 U4492 ( .A(n8921), .Y(n8916) );
  CLKBUFX3 U4493 ( .A(n8921), .Y(n8915) );
  CLKBUFX3 U4494 ( .A(n8921), .Y(n8914) );
  CLKBUFX3 U4495 ( .A(n8922), .Y(n8913) );
  CLKBUFX3 U4496 ( .A(n8922), .Y(n8912) );
  CLKBUFX3 U4497 ( .A(n8922), .Y(n8911) );
  CLKBUFX3 U4498 ( .A(n8846), .Y(n8845) );
  CLKBUFX3 U4499 ( .A(n8770), .Y(n8738) );
  CLKBUFX3 U4500 ( .A(n8770), .Y(n8737) );
  CLKBUFX3 U4501 ( .A(n8771), .Y(n8736) );
  CLKBUFX3 U4502 ( .A(n8771), .Y(n8735) );
  CLKBUFX3 U4503 ( .A(n8777), .Y(n8761) );
  CLKBUFX3 U4504 ( .A(n8910), .Y(n8909) );
  CLKBUFX3 U4505 ( .A(n8910), .Y(n8908) );
  CLKBUFX3 U4506 ( .A(n8776), .Y(n8763) );
  CLKBUFX3 U4507 ( .A(n8776), .Y(n8762) );
  CLKBUFX3 U4508 ( .A(n8777), .Y(n8760) );
  CLKBUFX3 U4509 ( .A(n8774), .Y(n8767) );
  CLKBUFX3 U4510 ( .A(n8773), .Y(n8768) );
  CLKBUFX3 U4511 ( .A(n8773), .Y(n8769) );
  CLKBUFX3 U4512 ( .A(n8775), .Y(n8765) );
  CLKBUFX3 U4513 ( .A(n8774), .Y(n8766) );
  CLKBUFX3 U4514 ( .A(n8775), .Y(n8764) );
  CLKBUFX3 U4515 ( .A(n8780), .Y(n8759) );
  CLKBUFX3 U4516 ( .A(n9145), .Y(n9143) );
  CLKBUFX3 U4517 ( .A(n9146), .Y(n9142) );
  CLKBUFX3 U4518 ( .A(n9146), .Y(n9141) );
  CLKBUFX3 U4519 ( .A(n9147), .Y(n9140) );
  CLKBUFX3 U4520 ( .A(n9147), .Y(n9139) );
  CLKBUFX3 U4521 ( .A(n9148), .Y(n9138) );
  CLKBUFX3 U4522 ( .A(n9148), .Y(n9137) );
  CLKBUFX3 U4523 ( .A(n9149), .Y(n9136) );
  CLKBUFX3 U4524 ( .A(n9149), .Y(n9135) );
  CLKBUFX3 U4525 ( .A(n9152), .Y(n9129) );
  CLKBUFX3 U4526 ( .A(n9152), .Y(n9130) );
  CLKBUFX3 U4527 ( .A(n9151), .Y(n9131) );
  CLKBUFX3 U4528 ( .A(n9151), .Y(n9132) );
  CLKBUFX3 U4529 ( .A(n9150), .Y(n9133) );
  CLKBUFX3 U4530 ( .A(n9150), .Y(n9134) );
  CLKBUFX3 U4531 ( .A(n8729), .Y(n8691) );
  CLKBUFX3 U4532 ( .A(n8729), .Y(n8692) );
  CLKBUFX3 U4533 ( .A(n8726), .Y(n8701) );
  CLKBUFX3 U4534 ( .A(n8726), .Y(n8700) );
  CLKBUFX3 U4535 ( .A(n8726), .Y(n8699) );
  CLKBUFX3 U4536 ( .A(n8725), .Y(n8704) );
  CLKBUFX3 U4537 ( .A(n8725), .Y(n8703) );
  CLKBUFX3 U4538 ( .A(n8725), .Y(n8702) );
  CLKBUFX3 U4539 ( .A(n8728), .Y(n8693) );
  CLKBUFX3 U4540 ( .A(n8727), .Y(n8698) );
  CLKBUFX3 U4541 ( .A(n8727), .Y(n8697) );
  CLKBUFX3 U4542 ( .A(n8727), .Y(n8696) );
  CLKBUFX3 U4543 ( .A(n8728), .Y(n8695) );
  CLKBUFX3 U4544 ( .A(n8728), .Y(n8694) );
  CLKBUFX3 U4545 ( .A(n8721), .Y(n8715) );
  CLKBUFX3 U4546 ( .A(n8721), .Y(n8714) );
  CLKBUFX3 U4547 ( .A(n8722), .Y(n8713) );
  CLKBUFX3 U4548 ( .A(n8720), .Y(n8718) );
  CLKBUFX3 U4549 ( .A(n8720), .Y(n8717) );
  CLKBUFX3 U4550 ( .A(n8721), .Y(n8716) );
  CLKBUFX3 U4551 ( .A(n8723), .Y(n8708) );
  CLKBUFX3 U4552 ( .A(n8724), .Y(n8707) );
  CLKBUFX3 U4553 ( .A(n8724), .Y(n8706) );
  CLKBUFX3 U4554 ( .A(n8724), .Y(n8705) );
  CLKBUFX3 U4555 ( .A(n8722), .Y(n8712) );
  CLKBUFX3 U4556 ( .A(n8722), .Y(n8711) );
  CLKBUFX3 U4557 ( .A(n8723), .Y(n8710) );
  CLKBUFX3 U4558 ( .A(n8723), .Y(n8709) );
  CLKBUFX3 U4559 ( .A(n8720), .Y(n8719) );
  CLKBUFX3 U4560 ( .A(n8791), .Y(n8782) );
  CLKBUFX3 U4561 ( .A(n8790), .Y(n8784) );
  CLKBUFX3 U4562 ( .A(n8789), .Y(n8785) );
  CLKBUFX3 U4563 ( .A(n8790), .Y(n8783) );
  CLKBUFX3 U4564 ( .A(n8791), .Y(n8781) );
  CLKBUFX3 U4565 ( .A(n8801), .Y(n8793) );
  CLKBUFX3 U4566 ( .A(n8789), .Y(n8786) );
  CLKBUFX3 U4567 ( .A(n8788), .Y(n8787) );
  CLKBUFX3 U4568 ( .A(n8800), .Y(n8796) );
  CLKBUFX3 U4569 ( .A(n8801), .Y(n8794) );
  CLKBUFX3 U4570 ( .A(n8799), .Y(n8797) );
  CLKBUFX3 U4571 ( .A(n8800), .Y(n8795) );
  CLKBUFX3 U4572 ( .A(n9145), .Y(n9144) );
  CLKBUFX3 U4573 ( .A(n8799), .Y(n8798) );
  CLKBUFX3 U4574 ( .A(n8849), .Y(n8839) );
  CLKBUFX3 U4575 ( .A(n6195), .Y(n8849) );
  CLKBUFX3 U4576 ( .A(n9464), .Y(n8791) );
  CLKBUFX3 U4577 ( .A(n9464), .Y(n8788) );
  CLKBUFX3 U4578 ( .A(n9465), .Y(n8800) );
  CLKBUFX3 U4579 ( .A(n9464), .Y(n8790) );
  CLKBUFX3 U4580 ( .A(n9465), .Y(n8799) );
  CLKBUFX3 U4581 ( .A(n9464), .Y(n8789) );
  CLKBUFX3 U4582 ( .A(n9465), .Y(n8801) );
  CLKBUFX3 U4583 ( .A(n9580), .Y(n8920) );
  CLKBUFX3 U4584 ( .A(n9580), .Y(n8921) );
  CLKBUFX3 U4585 ( .A(n9580), .Y(n8922) );
  CLKBUFX3 U4586 ( .A(n6195), .Y(n8848) );
  CLKBUFX3 U4587 ( .A(n8923), .Y(n8910) );
  CLKBUFX3 U4588 ( .A(n9580), .Y(n8923) );
  CLKBUFX3 U4589 ( .A(n6195), .Y(n8846) );
  CLKBUFX3 U4590 ( .A(n6195), .Y(n8847) );
  CLKBUFX3 U4591 ( .A(n8778), .Y(n8777) );
  CLKBUFX3 U4592 ( .A(n8778), .Y(n8776) );
  CLKBUFX3 U4593 ( .A(n8779), .Y(n8773) );
  CLKBUFX3 U4594 ( .A(n8779), .Y(n8774) );
  CLKBUFX3 U4595 ( .A(n8779), .Y(n8775) );
  CLKBUFX3 U4596 ( .A(n8772), .Y(n8770) );
  CLKBUFX3 U4597 ( .A(n8772), .Y(n8771) );
  CLKBUFX3 U4598 ( .A(n9156), .Y(n9146) );
  CLKBUFX3 U4599 ( .A(n9155), .Y(n9147) );
  CLKBUFX3 U4600 ( .A(n9155), .Y(n9148) );
  CLKBUFX3 U4601 ( .A(n9154), .Y(n9149) );
  CLKBUFX3 U4602 ( .A(n9153), .Y(n9152) );
  CLKBUFX3 U4603 ( .A(n9153), .Y(n9151) );
  CLKBUFX3 U4604 ( .A(n9154), .Y(n9150) );
  CLKBUFX3 U4605 ( .A(n9156), .Y(n9145) );
  CLKBUFX3 U4606 ( .A(n8731), .Y(n8726) );
  CLKBUFX3 U4607 ( .A(n8732), .Y(n8725) );
  CLKBUFX3 U4608 ( .A(n8731), .Y(n8727) );
  CLKBUFX3 U4609 ( .A(n8730), .Y(n8728) );
  CLKBUFX3 U4610 ( .A(n8734), .Y(n8721) );
  CLKBUFX3 U4611 ( .A(n8732), .Y(n8724) );
  CLKBUFX3 U4612 ( .A(n8733), .Y(n8722) );
  CLKBUFX3 U4613 ( .A(n8733), .Y(n8723) );
  CLKBUFX3 U4614 ( .A(n8734), .Y(n8720) );
  CLKBUFX3 U4615 ( .A(n8802), .Y(n8792) );
  CLKBUFX3 U4616 ( .A(n9465), .Y(n8802) );
  CLKBUFX3 U4617 ( .A(n8730), .Y(n8729) );
  CLKBUFX3 U4618 ( .A(n9158), .Y(n8730) );
  CLKBUFX3 U4619 ( .A(n9158), .Y(n8731) );
  CLKBUFX3 U4620 ( .A(n9158), .Y(n8732) );
  CLKBUFX3 U4621 ( .A(n9158), .Y(n8733) );
  CLKBUFX3 U4622 ( .A(n9158), .Y(n8734) );
  CLKBUFX3 U4623 ( .A(n10477), .Y(n9155) );
  CLKBUFX3 U4624 ( .A(n10477), .Y(n9153) );
  CLKBUFX3 U4625 ( .A(n10477), .Y(n9154) );
  CLKBUFX3 U4626 ( .A(n10477), .Y(n9156) );
  CLKBUFX3 U4627 ( .A(fir_valid), .Y(n8778) );
  CLKBUFX3 U4628 ( .A(fir_valid), .Y(n8779) );
  CLKBUFX3 U4629 ( .A(n8780), .Y(n8772) );
  CLKBUFX3 U4630 ( .A(fir_valid), .Y(n8780) );
  CLKINVX1 U4632 ( .A(rst), .Y(n10477) );
  CLKINVX1 U4633 ( .A(n9157), .Y(n10479) );
  MXI2X1 U4634 ( .A(n8689), .B(n9159), .S0(counter[0]), .Y(n6187) );
  NAND2X1 U4635 ( .A(n10470), .B(n9160), .Y(n6186) );
  MXI2X1 U4636 ( .A(n10470), .B(n11215), .S0(n8689), .Y(n6185) );
  MXI2X1 U4637 ( .A(n9161), .B(n9162), .S0(counter[1]), .Y(n6184) );
  NAND2X1 U4638 ( .A(data_valid), .B(counter[0]), .Y(n9161) );
  OAI32X1 U4639 ( .A0(n9163), .A1(n6074), .A2(n8689), .B0(n6073), .B1(n9164), 
        .Y(n6183) );
  OA21XL U4640 ( .A0(counter[1]), .A1(n8690), .B0(n9162), .Y(n9164) );
  OA21XL U4641 ( .A0(counter[0]), .A1(n8690), .B0(n9159), .Y(n9162) );
  MXI2X1 U4642 ( .A(n9165), .B(n9166), .S0(n6072), .Y(n6182) );
  NAND2X1 U4643 ( .A(n9167), .B(data_valid), .Y(n9166) );
  OA21XL U4644 ( .A0(n8690), .A1(n9167), .B0(n9159), .Y(n9165) );
  MXI2X1 U4645 ( .A(n9168), .B(n9169), .S0(n6189), .Y(n6181) );
  NAND2X1 U4646 ( .A(n9170), .B(data_valid), .Y(n9168) );
  OAI2BB1X1 U4647 ( .A0N(n9171), .A1N(n6191), .B0(n9160), .Y(n6180) );
  NAND4X1 U4648 ( .A(n6067), .B(n9170), .C(data_valid), .D(n6189), .Y(n9160)
         );
  OAI21XL U4649 ( .A0(n8689), .A1(n6189), .B0(n9169), .Y(n9171) );
  OA21XL U4650 ( .A0(n9170), .A1(n8690), .B0(n9159), .Y(n9169) );
  NAND2X1 U4651 ( .A(n10470), .B(n8689), .Y(n9159) );
  OAI21XL U4652 ( .A0(n9172), .A1(n6194), .B0(n9173), .Y(n6179) );
  NAND4X1 U4653 ( .A(n6068), .B(n9170), .C(n6191), .D(n6190), .Y(n9173) );
  NOR2X1 U4654 ( .A(n10472), .B(n9174), .Y(n9172) );
  OAI21XL U4655 ( .A0(n9174), .A1(n6194), .B0(n6190), .Y(n6178) );
  OAI21XL U4656 ( .A0(n3079), .A1(data_valid), .B0(n9175), .Y(n6064) );
  OAI21XL U4657 ( .A0(n3078), .A1(data_valid), .B0(n9175), .Y(n6062) );
  OAI21XL U4658 ( .A0(n3077), .A1(data_valid), .B0(n9175), .Y(n6061) );
  OAI21XL U4659 ( .A0(n3076), .A1(data_valid), .B0(n9175), .Y(n6060) );
  OAI21XL U4660 ( .A0(n3075), .A1(data_valid), .B0(n9175), .Y(n6059) );
  OAI21XL U4661 ( .A0(n3074), .A1(data_valid), .B0(n9175), .Y(n6058) );
  OAI21XL U4662 ( .A0(n3073), .A1(data_valid), .B0(n9175), .Y(n6057) );
  OAI21XL U4663 ( .A0(n3072), .A1(data_valid), .B0(n9175), .Y(n6056) );
  OAI21XL U4664 ( .A0(n3071), .A1(data_valid), .B0(n9175), .Y(n6055) );
  OAI21XL U4665 ( .A0(n30701), .A1(data_valid), .B0(n9175), .Y(n6054) );
  OAI21XL U4666 ( .A0(n3069), .A1(data_valid), .B0(n9175), .Y(n6053) );
  OAI21XL U4667 ( .A0(n3068), .A1(data_valid), .B0(n9175), .Y(n6052) );
  OAI21XL U4668 ( .A0(n3067), .A1(data_valid), .B0(n9175), .Y(n6051) );
  NAND2X1 U4669 ( .A(hd01_35), .B(data_valid), .Y(n9175) );
  CLKMX2X2 U4670 ( .A(hd01[22]), .B(d01[22]), .S0(n8604), .Y(n6050) );
  CLKMX2X2 U4671 ( .A(hd01[21]), .B(d01[21]), .S0(n8636), .Y(n6049) );
  CLKMX2X2 U4672 ( .A(hd01[20]), .B(d01[20]), .S0(n8636), .Y(n6048) );
  CLKMX2X2 U4673 ( .A(hd01[19]), .B(d01[19]), .S0(n8635), .Y(n6047) );
  CLKMX2X2 U4674 ( .A(hd01[18]), .B(d01[18]), .S0(n8635), .Y(n6046) );
  CLKMX2X2 U4675 ( .A(hd01[17]), .B(d01[17]), .S0(n8635), .Y(n6045) );
  CLKMX2X2 U4676 ( .A(hd01[16]), .B(d01[16]), .S0(n8635), .Y(n6044) );
  CLKMX2X2 U4677 ( .A(hd01[15]), .B(d01[15]), .S0(n8635), .Y(n6043) );
  CLKMX2X2 U4678 ( .A(hd01[14]), .B(d01[14]), .S0(n8635), .Y(n6042) );
  CLKMX2X2 U4679 ( .A(hd01[13]), .B(d01[13]), .S0(n8635), .Y(n6041) );
  CLKMX2X2 U4680 ( .A(hd01[12]), .B(d01[12]), .S0(n8635), .Y(n6040) );
  CLKMX2X2 U4681 ( .A(hd01[11]), .B(d01[11]), .S0(n8635), .Y(n6039) );
  CLKMX2X2 U4682 ( .A(hd01[10]), .B(d01[10]), .S0(n8635), .Y(n6038) );
  CLKMX2X2 U4683 ( .A(hd01[9]), .B(d01[9]), .S0(n8635), .Y(n6037) );
  CLKMX2X2 U4684 ( .A(hd01[8]), .B(d01[8]), .S0(n8635), .Y(n6036) );
  CLKMX2X2 U4685 ( .A(hd01[7]), .B(d01[7]), .S0(n8635), .Y(n6035) );
  CLKMX2X2 U4686 ( .A(hd01[6]), .B(d01[6]), .S0(n8634), .Y(n6034) );
  CLKMX2X2 U4687 ( .A(hd01[5]), .B(d01[5]), .S0(n8634), .Y(n6033) );
  CLKMX2X2 U4688 ( .A(hd01[4]), .B(d01[4]), .S0(n8634), .Y(n6032) );
  CLKMX2X2 U4689 ( .A(hd01[3]), .B(d01[3]), .S0(n8634), .Y(n6031) );
  CLKMX2X2 U4690 ( .A(hd01[2]), .B(d01[2]), .S0(n8634), .Y(n6030) );
  CLKMX2X2 U4691 ( .A(hd01[1]), .B(d01[1]), .S0(n8634), .Y(n6029) );
  CLKMX2X2 U4692 ( .A(hd_a02[35]), .B(d02[35]), .S0(n8634), .Y(n6027) );
  CLKMX2X2 U4693 ( .A(hd_a02[34]), .B(d02[34]), .S0(n8634), .Y(n6026) );
  CLKMX2X2 U4694 ( .A(hd_a02[33]), .B(d02[33]), .S0(n8634), .Y(n6025) );
  CLKMX2X2 U4695 ( .A(hd_a02[32]), .B(d02[32]), .S0(n8634), .Y(n6024) );
  CLKMX2X2 U4696 ( .A(hd_a02[31]), .B(d02[31]), .S0(n8634), .Y(n6023) );
  CLKMX2X2 U4697 ( .A(hd_a02[30]), .B(d02[30]), .S0(n8634), .Y(n6022) );
  CLKMX2X2 U4698 ( .A(hd_a02[29]), .B(d02[29]), .S0(n8634), .Y(n6021) );
  CLKMX2X2 U4699 ( .A(hd_a02[28]), .B(d02[28]), .S0(n8633), .Y(n6020) );
  CLKMX2X2 U4700 ( .A(hd_a02[27]), .B(d02[27]), .S0(n8633), .Y(n6019) );
  CLKMX2X2 U4701 ( .A(hd_a02[26]), .B(d02[26]), .S0(n8633), .Y(n6018) );
  CLKMX2X2 U4702 ( .A(hd_a02[25]), .B(d02[25]), .S0(n8633), .Y(n6017) );
  CLKMX2X2 U4703 ( .A(hd_a02[24]), .B(d02[24]), .S0(n8633), .Y(n6016) );
  CLKMX2X2 U4704 ( .A(hd_a02[23]), .B(d02[23]), .S0(n8633), .Y(n6015) );
  CLKMX2X2 U4705 ( .A(hd_a02[22]), .B(d02[22]), .S0(n8633), .Y(n6014) );
  CLKMX2X2 U4706 ( .A(hd_a02[21]), .B(d02[21]), .S0(n8633), .Y(n6013) );
  CLKMX2X2 U4707 ( .A(hd_a02[20]), .B(d02[20]), .S0(n8633), .Y(n6012) );
  CLKMX2X2 U4708 ( .A(hd_a02[19]), .B(d02[19]), .S0(n8633), .Y(n6011) );
  CLKMX2X2 U4709 ( .A(hd_a02[18]), .B(d02[18]), .S0(n8633), .Y(n6010) );
  CLKMX2X2 U4710 ( .A(hd_a02[17]), .B(d02[17]), .S0(n8633), .Y(n6009) );
  CLKMX2X2 U4711 ( .A(hd_a02[16]), .B(d02[16]), .S0(n8633), .Y(n6008) );
  CLKMX2X2 U4712 ( .A(hd_a02[15]), .B(d02[15]), .S0(n8632), .Y(n6007) );
  CLKMX2X2 U4713 ( .A(hd_a02[14]), .B(d02[14]), .S0(n8632), .Y(n6006) );
  CLKMX2X2 U4714 ( .A(hd_a02[13]), .B(d02[13]), .S0(n8632), .Y(n6005) );
  CLKMX2X2 U4715 ( .A(hd_a02[12]), .B(d02[12]), .S0(n8632), .Y(n6004) );
  CLKMX2X2 U4716 ( .A(hd_a02[11]), .B(d02[11]), .S0(n8632), .Y(n6003) );
  CLKMX2X2 U4717 ( .A(hd_a02[10]), .B(d02[10]), .S0(n8632), .Y(n6002) );
  CLKMX2X2 U4718 ( .A(hd_a02[9]), .B(d02[9]), .S0(n8632), .Y(n6001) );
  CLKMX2X2 U4719 ( .A(hd_a02[8]), .B(d02[8]), .S0(n8632), .Y(n6000) );
  CLKMX2X2 U4720 ( .A(hd_a02[7]), .B(d02[7]), .S0(n8632), .Y(n5999) );
  CLKMX2X2 U4721 ( .A(hd_a02[6]), .B(d02[6]), .S0(n8632), .Y(n5998) );
  CLKMX2X2 U4722 ( .A(hd_a02[5]), .B(d02[5]), .S0(n8632), .Y(n5997) );
  CLKMX2X2 U4723 ( .A(hd_a02[4]), .B(d02[4]), .S0(n8632), .Y(n5996) );
  CLKMX2X2 U4724 ( .A(hd_a02[3]), .B(d02[3]), .S0(n8632), .Y(n5995) );
  CLKMX2X2 U4725 ( .A(hd_a02[2]), .B(d02[2]), .S0(n8631), .Y(n5994) );
  CLKMX2X2 U4726 ( .A(hd_a02[1]), .B(d02[1]), .S0(n8631), .Y(n5993) );
  CLKMX2X2 U4727 ( .A(hd_a03[35]), .B(d03[35]), .S0(n8631), .Y(n5991) );
  CLKMX2X2 U4728 ( .A(hd_a03[34]), .B(d03[34]), .S0(n8631), .Y(n5990) );
  CLKMX2X2 U4729 ( .A(hd_a03[33]), .B(d03[33]), .S0(n8631), .Y(n5989) );
  CLKMX2X2 U4730 ( .A(hd_a03[32]), .B(d03[32]), .S0(n8631), .Y(n5988) );
  CLKMX2X2 U4731 ( .A(hd_a03[31]), .B(d03[31]), .S0(n8631), .Y(n5987) );
  CLKMX2X2 U4732 ( .A(hd_a03[30]), .B(d03[30]), .S0(n8631), .Y(n5986) );
  CLKMX2X2 U4733 ( .A(hd_a03[29]), .B(d03[29]), .S0(n8631), .Y(n5985) );
  CLKMX2X2 U4734 ( .A(hd_a03[28]), .B(d03[28]), .S0(n8631), .Y(n5984) );
  CLKMX2X2 U4735 ( .A(hd_a03[27]), .B(d03[27]), .S0(n8631), .Y(n5983) );
  CLKMX2X2 U4736 ( .A(hd_a03[26]), .B(d03[26]), .S0(n8631), .Y(n5982) );
  CLKMX2X2 U4737 ( .A(hd_a03[25]), .B(d03[25]), .S0(n8630), .Y(n5981) );
  CLKMX2X2 U4738 ( .A(hd_a03[24]), .B(d03[24]), .S0(n8630), .Y(n5980) );
  CLKMX2X2 U4739 ( .A(hd_a03[23]), .B(d03[23]), .S0(n8630), .Y(n5979) );
  CLKMX2X2 U4740 ( .A(hd_a03[22]), .B(d03[22]), .S0(n8630), .Y(n5978) );
  CLKMX2X2 U4741 ( .A(hd_a03[21]), .B(d03[21]), .S0(n8630), .Y(n5977) );
  CLKMX2X2 U4742 ( .A(hd_a03[20]), .B(d03[20]), .S0(n8630), .Y(n5976) );
  CLKMX2X2 U4743 ( .A(hd_a03[19]), .B(d03[19]), .S0(n8630), .Y(n5975) );
  CLKMX2X2 U4744 ( .A(hd_a03[18]), .B(d03[18]), .S0(n8630), .Y(n5974) );
  CLKMX2X2 U4745 ( .A(hd_a03[17]), .B(d03[17]), .S0(n8630), .Y(n5973) );
  CLKMX2X2 U4746 ( .A(hd_a03[16]), .B(d03[16]), .S0(n8630), .Y(n5972) );
  CLKMX2X2 U4747 ( .A(hd_a03[15]), .B(d03[15]), .S0(n8630), .Y(n5971) );
  CLKMX2X2 U4748 ( .A(hd_a03[14]), .B(d03[14]), .S0(n8630), .Y(n5970) );
  CLKMX2X2 U4749 ( .A(hd_a03[13]), .B(d03[13]), .S0(n8629), .Y(n5969) );
  CLKMX2X2 U4750 ( .A(hd_a03[12]), .B(d03[12]), .S0(n8629), .Y(n5968) );
  CLKMX2X2 U4751 ( .A(hd_a03[11]), .B(d03[11]), .S0(n8629), .Y(n5967) );
  CLKMX2X2 U4752 ( .A(hd_a03[10]), .B(d03[10]), .S0(n8629), .Y(n5966) );
  CLKMX2X2 U4753 ( .A(hd_a03[9]), .B(d03[9]), .S0(n8629), .Y(n5965) );
  CLKMX2X2 U4754 ( .A(hd_a03[8]), .B(d03[8]), .S0(n8629), .Y(n5964) );
  CLKMX2X2 U4755 ( .A(hd_a03[7]), .B(d03[7]), .S0(n8629), .Y(n5963) );
  CLKMX2X2 U4756 ( .A(hd_a03[6]), .B(d03[6]), .S0(n8629), .Y(n5962) );
  CLKMX2X2 U4757 ( .A(hd_a03[5]), .B(d03[5]), .S0(n8629), .Y(n5961) );
  CLKMX2X2 U4758 ( .A(hd_a03[4]), .B(d03[4]), .S0(n8629), .Y(n5960) );
  CLKMX2X2 U4759 ( .A(hd_a03[3]), .B(d03[3]), .S0(n8629), .Y(n5959) );
  CLKMX2X2 U4760 ( .A(hd_a03[2]), .B(d03[2]), .S0(n8629), .Y(n5958) );
  CLKMX2X2 U4761 ( .A(hd_a03[1]), .B(d03[1]), .S0(n8629), .Y(n5957) );
  CLKMX2X2 U4762 ( .A(hd_a03[0]), .B(d03[0]), .S0(n8628), .Y(n5956) );
  CLKMX2X2 U4763 ( .A(hd_a04[35]), .B(d04[35]), .S0(n8628), .Y(n5955) );
  CLKMX2X2 U4764 ( .A(hd_a04[34]), .B(d04[34]), .S0(n8628), .Y(n5954) );
  CLKMX2X2 U4765 ( .A(hd_a04[33]), .B(d04[33]), .S0(n8628), .Y(n5953) );
  CLKMX2X2 U4766 ( .A(hd_a04[32]), .B(d04[32]), .S0(n8628), .Y(n5952) );
  CLKMX2X2 U4767 ( .A(hd_a04[31]), .B(d04[31]), .S0(n8628), .Y(n5951) );
  CLKMX2X2 U4768 ( .A(hd_a04[30]), .B(d04[30]), .S0(n8628), .Y(n5950) );
  CLKMX2X2 U4769 ( .A(hd_a04[29]), .B(d04[29]), .S0(n8628), .Y(n5949) );
  CLKMX2X2 U4770 ( .A(hd_a04[28]), .B(d04[28]), .S0(n8628), .Y(n5948) );
  CLKMX2X2 U4771 ( .A(hd_a04[27]), .B(d04[27]), .S0(n8628), .Y(n5947) );
  CLKMX2X2 U4772 ( .A(hd_a04[26]), .B(d04[26]), .S0(n8628), .Y(n5946) );
  CLKMX2X2 U4773 ( .A(hd_a04[25]), .B(d04[25]), .S0(n8628), .Y(n5945) );
  CLKMX2X2 U4774 ( .A(hd_a04[24]), .B(d04[24]), .S0(n8628), .Y(n5944) );
  CLKMX2X2 U4775 ( .A(hd_a04[23]), .B(d04[23]), .S0(n8627), .Y(n5943) );
  CLKMX2X2 U4776 ( .A(hd_a04[22]), .B(d04[22]), .S0(n8627), .Y(n5942) );
  CLKMX2X2 U4777 ( .A(hd_a04[21]), .B(d04[21]), .S0(n8627), .Y(n5941) );
  CLKMX2X2 U4778 ( .A(hd_a04[20]), .B(d04[20]), .S0(n8627), .Y(n5940) );
  CLKMX2X2 U4779 ( .A(hd_a04[19]), .B(d04[19]), .S0(n8627), .Y(n5939) );
  CLKMX2X2 U4780 ( .A(hd_a04[18]), .B(d04[18]), .S0(n8627), .Y(n5938) );
  CLKMX2X2 U4781 ( .A(hd_a04[17]), .B(d04[17]), .S0(n8627), .Y(n5937) );
  CLKMX2X2 U4782 ( .A(hd_a04[16]), .B(d04[16]), .S0(n8627), .Y(n5936) );
  CLKMX2X2 U4783 ( .A(hd_a04[15]), .B(d04[15]), .S0(n8627), .Y(n5935) );
  CLKMX2X2 U4784 ( .A(hd_a04[14]), .B(d04[14]), .S0(n8627), .Y(n5934) );
  CLKMX2X2 U4785 ( .A(hd_a04[13]), .B(d04[13]), .S0(n8627), .Y(n5933) );
  CLKMX2X2 U4786 ( .A(hd_a04[12]), .B(d04[12]), .S0(n8627), .Y(n5932) );
  CLKMX2X2 U4787 ( .A(hd_a04[11]), .B(d04[11]), .S0(n8627), .Y(n5931) );
  CLKMX2X2 U4788 ( .A(hd_a04[10]), .B(d04[10]), .S0(n8626), .Y(n5930) );
  CLKMX2X2 U4789 ( .A(hd_a04[9]), .B(d04[9]), .S0(n8626), .Y(n5929) );
  CLKMX2X2 U4790 ( .A(hd_a04[8]), .B(d04[8]), .S0(n8626), .Y(n5928) );
  CLKMX2X2 U4791 ( .A(hd_a04[7]), .B(d04[7]), .S0(n8626), .Y(n5927) );
  CLKMX2X2 U4792 ( .A(hd_a04[6]), .B(d04[6]), .S0(n8626), .Y(n5926) );
  CLKMX2X2 U4793 ( .A(hd_a04[5]), .B(d04[5]), .S0(n8626), .Y(n5925) );
  CLKMX2X2 U4794 ( .A(hd_a04[4]), .B(d04[4]), .S0(n8626), .Y(n5924) );
  CLKMX2X2 U4795 ( .A(hd_a04[3]), .B(d04[3]), .S0(n8626), .Y(n5923) );
  CLKMX2X2 U4796 ( .A(hd_a04[2]), .B(d04[2]), .S0(n8626), .Y(n5922) );
  CLKMX2X2 U4797 ( .A(hd_a04[1]), .B(d04[1]), .S0(n8626), .Y(n5921) );
  CLKMX2X2 U4798 ( .A(hd_a04[0]), .B(d04[0]), .S0(n8626), .Y(n5920) );
  CLKMX2X2 U4799 ( .A(hd_a05[35]), .B(d05[35]), .S0(n8626), .Y(n5919) );
  CLKMX2X2 U4800 ( .A(hd_a05[34]), .B(d05[34]), .S0(n8626), .Y(n5918) );
  CLKMX2X2 U4801 ( .A(hd_a05[33]), .B(d05[33]), .S0(n8625), .Y(n5917) );
  CLKMX2X2 U4802 ( .A(hd_a05[32]), .B(d05[32]), .S0(n8625), .Y(n5916) );
  CLKMX2X2 U4803 ( .A(hd_a05[31]), .B(d05[31]), .S0(n8625), .Y(n5915) );
  CLKMX2X2 U4804 ( .A(hd_a05[30]), .B(d05[30]), .S0(n8625), .Y(n5914) );
  CLKMX2X2 U4805 ( .A(hd_a05[29]), .B(d05[29]), .S0(n8625), .Y(n5913) );
  CLKMX2X2 U4806 ( .A(hd_a05[28]), .B(d05[28]), .S0(n8625), .Y(n5912) );
  CLKMX2X2 U4807 ( .A(hd_a05[27]), .B(d05[27]), .S0(n8625), .Y(n5911) );
  CLKMX2X2 U4808 ( .A(hd_a05[26]), .B(d05[26]), .S0(n8630), .Y(n5910) );
  CLKMX2X2 U4809 ( .A(hd_a05[25]), .B(d05[25]), .S0(n8646), .Y(n5909) );
  CLKMX2X2 U4810 ( .A(hd_a05[24]), .B(d05[24]), .S0(n8646), .Y(n5908) );
  CLKMX2X2 U4811 ( .A(hd_a05[23]), .B(d05[23]), .S0(n8646), .Y(n5907) );
  CLKMX2X2 U4812 ( .A(hd_a05[22]), .B(d05[22]), .S0(n8646), .Y(n5906) );
  CLKMX2X2 U4813 ( .A(hd_a05[21]), .B(d05[21]), .S0(n8646), .Y(n5905) );
  CLKMX2X2 U4814 ( .A(hd_a05[20]), .B(d05[20]), .S0(n8646), .Y(n5904) );
  CLKMX2X2 U4815 ( .A(hd_a05[19]), .B(d05[19]), .S0(n8646), .Y(n5903) );
  CLKMX2X2 U4816 ( .A(hd_a05[18]), .B(d05[18]), .S0(n8646), .Y(n5902) );
  CLKMX2X2 U4817 ( .A(hd_a05[17]), .B(d05[17]), .S0(n8646), .Y(n5901) );
  CLKMX2X2 U4818 ( .A(hd_a05[16]), .B(d05[16]), .S0(n8646), .Y(n5900) );
  CLKMX2X2 U4819 ( .A(hd_a05[15]), .B(d05[15]), .S0(n8646), .Y(n5899) );
  CLKMX2X2 U4820 ( .A(hd_a05[14]), .B(d05[14]), .S0(n8645), .Y(n5898) );
  CLKMX2X2 U4821 ( .A(hd_a05[13]), .B(d05[13]), .S0(n8645), .Y(n5897) );
  CLKMX2X2 U4822 ( .A(hd_a05[12]), .B(d05[12]), .S0(n8645), .Y(n5896) );
  CLKMX2X2 U4823 ( .A(hd_a05[11]), .B(d05[11]), .S0(n8645), .Y(n5895) );
  CLKMX2X2 U4824 ( .A(hd_a05[10]), .B(d05[10]), .S0(n8645), .Y(n5894) );
  CLKMX2X2 U4825 ( .A(hd_a05[9]), .B(d05[9]), .S0(n8645), .Y(n5893) );
  CLKMX2X2 U4826 ( .A(hd_a05[8]), .B(d05[8]), .S0(n8645), .Y(n5892) );
  CLKMX2X2 U4827 ( .A(hd_a05[7]), .B(d05[7]), .S0(n8645), .Y(n5891) );
  CLKMX2X2 U4828 ( .A(hd_a05[6]), .B(d05[6]), .S0(n8645), .Y(n5890) );
  CLKMX2X2 U4829 ( .A(hd_a05[5]), .B(d05[5]), .S0(n8645), .Y(n5889) );
  CLKMX2X2 U4830 ( .A(hd_a05[4]), .B(d05[4]), .S0(n8645), .Y(n5888) );
  CLKMX2X2 U4831 ( .A(hd_a05[3]), .B(d05[3]), .S0(n8645), .Y(n5887) );
  CLKMX2X2 U4832 ( .A(hd_a05[2]), .B(d05[2]), .S0(n8645), .Y(n5886) );
  CLKMX2X2 U4833 ( .A(hd_a05[1]), .B(d05[1]), .S0(n8644), .Y(n5885) );
  CLKMX2X2 U4834 ( .A(hd_a05[0]), .B(d05[0]), .S0(n8644), .Y(n5884) );
  CLKMX2X2 U4835 ( .A(hd_a06[35]), .B(d06[35]), .S0(n8644), .Y(n5883) );
  CLKMX2X2 U4836 ( .A(hd_a06[34]), .B(d06[34]), .S0(n8644), .Y(n5882) );
  CLKMX2X2 U4837 ( .A(hd_a06[33]), .B(d06[33]), .S0(n8644), .Y(n5881) );
  CLKMX2X2 U4838 ( .A(hd_a06[32]), .B(d06[32]), .S0(n8644), .Y(n5880) );
  CLKMX2X2 U4839 ( .A(hd_a06[31]), .B(d06[31]), .S0(n8644), .Y(n5879) );
  CLKMX2X2 U4840 ( .A(hd_a06[30]), .B(d06[30]), .S0(n8644), .Y(n5878) );
  CLKMX2X2 U4841 ( .A(hd_a06[29]), .B(d06[29]), .S0(n8644), .Y(n5877) );
  CLKMX2X2 U4842 ( .A(hd_a06[28]), .B(d06[28]), .S0(n8644), .Y(n5876) );
  CLKMX2X2 U4843 ( .A(hd_a06[27]), .B(d06[27]), .S0(n8644), .Y(n5875) );
  CLKMX2X2 U4844 ( .A(hd_a06[26]), .B(d06[26]), .S0(n8644), .Y(n5874) );
  CLKMX2X2 U4845 ( .A(hd_a06[25]), .B(d06[25]), .S0(n8644), .Y(n5873) );
  CLKMX2X2 U4846 ( .A(hd_a06[24]), .B(d06[24]), .S0(n8643), .Y(n5872) );
  CLKMX2X2 U4847 ( .A(hd_a06[23]), .B(d06[23]), .S0(n8643), .Y(n5871) );
  CLKMX2X2 U4848 ( .A(hd_a06[22]), .B(d06[22]), .S0(n8643), .Y(n5870) );
  CLKMX2X2 U4849 ( .A(hd_a06[21]), .B(d06[21]), .S0(n8643), .Y(n5869) );
  CLKMX2X2 U4850 ( .A(hd_a06[20]), .B(d06[20]), .S0(n8643), .Y(n5868) );
  CLKMX2X2 U4851 ( .A(hd_a06[19]), .B(d06[19]), .S0(n8643), .Y(n5867) );
  CLKMX2X2 U4852 ( .A(hd_a06[18]), .B(d06[18]), .S0(n8643), .Y(n5866) );
  CLKMX2X2 U4853 ( .A(hd_a06[17]), .B(d06[17]), .S0(n8643), .Y(n5865) );
  CLKMX2X2 U4854 ( .A(hd_a06[16]), .B(d06[16]), .S0(n8643), .Y(n5864) );
  CLKMX2X2 U4855 ( .A(hd_a06[15]), .B(d06[15]), .S0(n8643), .Y(n5863) );
  CLKMX2X2 U4856 ( .A(hd_a06[14]), .B(d06[14]), .S0(n8643), .Y(n5862) );
  CLKMX2X2 U4857 ( .A(hd_a06[13]), .B(d06[13]), .S0(n8643), .Y(n5861) );
  CLKMX2X2 U4858 ( .A(hd_a06[12]), .B(d06[12]), .S0(n8643), .Y(n5860) );
  CLKMX2X2 U4859 ( .A(hd_a06[11]), .B(d06[11]), .S0(n8642), .Y(n5859) );
  CLKMX2X2 U4860 ( .A(hd_a06[10]), .B(d06[10]), .S0(n8642), .Y(n5858) );
  CLKMX2X2 U4861 ( .A(hd_a06[9]), .B(d06[9]), .S0(n8642), .Y(n5857) );
  CLKMX2X2 U4862 ( .A(hd_a06[8]), .B(d06[8]), .S0(n8642), .Y(n5856) );
  CLKMX2X2 U4863 ( .A(hd_a06[7]), .B(d06[7]), .S0(n8642), .Y(n5855) );
  CLKMX2X2 U4864 ( .A(hd_a06[6]), .B(d06[6]), .S0(n8642), .Y(n5854) );
  CLKMX2X2 U4865 ( .A(hd_a06[5]), .B(d06[5]), .S0(n8642), .Y(n5853) );
  CLKMX2X2 U4866 ( .A(hd_a06[4]), .B(d06[4]), .S0(n8642), .Y(n5852) );
  CLKMX2X2 U4867 ( .A(hd_a06[3]), .B(d06[3]), .S0(n8642), .Y(n5851) );
  CLKMX2X2 U4868 ( .A(hd_a06[2]), .B(d06[2]), .S0(n8642), .Y(n5850) );
  CLKMX2X2 U4869 ( .A(hd_a06[1]), .B(d06[1]), .S0(n8642), .Y(n5849) );
  CLKMX2X2 U4870 ( .A(hd_a06[0]), .B(d06[0]), .S0(n8642), .Y(n5848) );
  CLKMX2X2 U4871 ( .A(hd_a07[35]), .B(d07[35]), .S0(n8642), .Y(n5847) );
  CLKMX2X2 U4872 ( .A(hd_a07[34]), .B(d07[34]), .S0(n8641), .Y(n5846) );
  CLKMX2X2 U4873 ( .A(hd_a07[33]), .B(d07[33]), .S0(n8641), .Y(n5845) );
  CLKMX2X2 U4874 ( .A(hd_a07[32]), .B(d07[32]), .S0(n8641), .Y(n5844) );
  CLKMX2X2 U4875 ( .A(hd_a07[31]), .B(d07[31]), .S0(n8641), .Y(n5843) );
  CLKMX2X2 U4876 ( .A(hd_a07[30]), .B(d07[30]), .S0(n8641), .Y(n5842) );
  CLKMX2X2 U4877 ( .A(hd_a07[29]), .B(d07[29]), .S0(n8641), .Y(n5841) );
  CLKMX2X2 U4878 ( .A(hd_a07[28]), .B(d07[28]), .S0(n8641), .Y(n5840) );
  CLKMX2X2 U4879 ( .A(hd_a07[27]), .B(d07[27]), .S0(n8641), .Y(n5839) );
  CLKMX2X2 U4880 ( .A(hd_a07[26]), .B(d07[26]), .S0(n8641), .Y(n5838) );
  CLKMX2X2 U4881 ( .A(hd_a07[25]), .B(d07[25]), .S0(n8641), .Y(n5837) );
  CLKMX2X2 U4882 ( .A(hd_a07[24]), .B(d07[24]), .S0(n8641), .Y(n5836) );
  CLKMX2X2 U4883 ( .A(hd_a07[23]), .B(d07[23]), .S0(n8641), .Y(n5835) );
  CLKMX2X2 U4884 ( .A(hd_a07[22]), .B(d07[22]), .S0(n8640), .Y(n5834) );
  CLKMX2X2 U4885 ( .A(hd_a07[21]), .B(d07[21]), .S0(n8640), .Y(n5833) );
  CLKMX2X2 U4886 ( .A(hd_a07[20]), .B(d07[20]), .S0(n8640), .Y(n5832) );
  CLKMX2X2 U4887 ( .A(hd_a07[19]), .B(d07[19]), .S0(n8640), .Y(n5831) );
  CLKMX2X2 U4888 ( .A(hd_a07[18]), .B(d07[18]), .S0(n8640), .Y(n5830) );
  CLKMX2X2 U4889 ( .A(hd_a07[17]), .B(d07[17]), .S0(n8640), .Y(n5829) );
  CLKMX2X2 U4890 ( .A(hd_a07[16]), .B(d07[16]), .S0(n8640), .Y(n5828) );
  CLKMX2X2 U4891 ( .A(hd_a07[15]), .B(d07[15]), .S0(n8640), .Y(n5827) );
  CLKMX2X2 U4892 ( .A(hd_a07[14]), .B(d07[14]), .S0(n8640), .Y(n5826) );
  CLKMX2X2 U4893 ( .A(hd_a07[13]), .B(d07[13]), .S0(n8640), .Y(n5825) );
  CLKMX2X2 U4894 ( .A(hd_a07[12]), .B(d07[12]), .S0(n8640), .Y(n5824) );
  CLKMX2X2 U4895 ( .A(hd_a07[11]), .B(d07[11]), .S0(n8640), .Y(n5823) );
  CLKMX2X2 U4896 ( .A(hd_a07[10]), .B(d07[10]), .S0(n8640), .Y(n5822) );
  CLKMX2X2 U4897 ( .A(hd_a07[9]), .B(d07[9]), .S0(n8639), .Y(n5821) );
  CLKMX2X2 U4898 ( .A(hd_a07[8]), .B(d07[8]), .S0(n8639), .Y(n5820) );
  CLKMX2X2 U4899 ( .A(hd_a07[7]), .B(d07[7]), .S0(n8639), .Y(n5819) );
  CLKMX2X2 U4900 ( .A(hd_a07[6]), .B(d07[6]), .S0(n8639), .Y(n5818) );
  CLKMX2X2 U4901 ( .A(hd_a07[5]), .B(d07[5]), .S0(n8639), .Y(n5817) );
  CLKMX2X2 U4902 ( .A(hd_a07[4]), .B(d07[4]), .S0(n8639), .Y(n5816) );
  CLKMX2X2 U4903 ( .A(hd_a07[3]), .B(d07[3]), .S0(n8639), .Y(n5815) );
  CLKMX2X2 U4904 ( .A(hd_a07[2]), .B(d07[2]), .S0(n8639), .Y(n5814) );
  CLKMX2X2 U4905 ( .A(hd_a07[1]), .B(d07[1]), .S0(n8639), .Y(n5813) );
  CLKMX2X2 U4906 ( .A(hd_a07[0]), .B(d07[0]), .S0(n8639), .Y(n5812) );
  CLKMX2X2 U4907 ( .A(hd_a08[35]), .B(d08[35]), .S0(n8639), .Y(n5811) );
  CLKMX2X2 U4908 ( .A(hd_a08[34]), .B(d08[34]), .S0(n8639), .Y(n5810) );
  CLKMX2X2 U4909 ( .A(hd_a08[33]), .B(d08[33]), .S0(n8639), .Y(n5809) );
  CLKMX2X2 U4910 ( .A(hd_a08[32]), .B(d08[32]), .S0(n8638), .Y(n5808) );
  CLKMX2X2 U4911 ( .A(hd_a08[31]), .B(d08[31]), .S0(n8638), .Y(n5807) );
  CLKMX2X2 U4912 ( .A(hd_a08[30]), .B(d08[30]), .S0(n8638), .Y(n5806) );
  CLKMX2X2 U4913 ( .A(hd_a08[29]), .B(d08[29]), .S0(n8638), .Y(n5805) );
  CLKMX2X2 U4914 ( .A(hd_a08[28]), .B(d08[28]), .S0(n8638), .Y(n5804) );
  CLKMX2X2 U4915 ( .A(hd_a08[27]), .B(d08[27]), .S0(n8638), .Y(n5803) );
  CLKMX2X2 U4916 ( .A(hd_a08[26]), .B(d08[26]), .S0(n8638), .Y(n5802) );
  CLKMX2X2 U4917 ( .A(hd_a08[25]), .B(d08[25]), .S0(n8638), .Y(n5801) );
  CLKMX2X2 U4918 ( .A(hd_a08[24]), .B(d08[24]), .S0(n8638), .Y(n5800) );
  CLKMX2X2 U4919 ( .A(hd_a08[23]), .B(d08[23]), .S0(n8638), .Y(n5799) );
  CLKMX2X2 U4920 ( .A(hd_a08[22]), .B(d08[22]), .S0(n8638), .Y(n5798) );
  CLKMX2X2 U4921 ( .A(hd_a08[21]), .B(d08[21]), .S0(n8638), .Y(n5797) );
  CLKMX2X2 U4922 ( .A(hd_a08[20]), .B(d08[20]), .S0(n8638), .Y(n5796) );
  CLKMX2X2 U4923 ( .A(hd_a08[19]), .B(d08[19]), .S0(n8637), .Y(n5795) );
  CLKMX2X2 U4924 ( .A(hd_a08[18]), .B(d08[18]), .S0(n8637), .Y(n5794) );
  CLKMX2X2 U4925 ( .A(hd_a08[17]), .B(d08[17]), .S0(n8637), .Y(n5793) );
  CLKMX2X2 U4926 ( .A(hd_a08[16]), .B(d08[16]), .S0(n8637), .Y(n5792) );
  CLKMX2X2 U4927 ( .A(hd_a08[15]), .B(d08[15]), .S0(n8637), .Y(n5791) );
  CLKMX2X2 U4928 ( .A(hd_a08[14]), .B(d08[14]), .S0(n8637), .Y(n5790) );
  CLKMX2X2 U4929 ( .A(hd_a08[13]), .B(d08[13]), .S0(n8637), .Y(n5789) );
  CLKMX2X2 U4930 ( .A(hd_a08[12]), .B(d08[12]), .S0(n8637), .Y(n5788) );
  CLKMX2X2 U4931 ( .A(hd_a08[11]), .B(d08[11]), .S0(n8637), .Y(n5787) );
  CLKMX2X2 U4932 ( .A(hd_a08[10]), .B(d08[10]), .S0(n8637), .Y(n5786) );
  CLKMX2X2 U4933 ( .A(hd_a08[9]), .B(d08[9]), .S0(n8637), .Y(n5785) );
  CLKMX2X2 U4934 ( .A(hd_a08[8]), .B(d08[8]), .S0(n8637), .Y(n5784) );
  CLKMX2X2 U4935 ( .A(hd_a08[7]), .B(d08[7]), .S0(n8637), .Y(n5783) );
  CLKMX2X2 U4936 ( .A(hd_a08[6]), .B(d08[6]), .S0(n8636), .Y(n5782) );
  CLKMX2X2 U4937 ( .A(hd_a08[5]), .B(d08[5]), .S0(n8636), .Y(n5781) );
  CLKMX2X2 U4938 ( .A(hd_a08[4]), .B(d08[4]), .S0(n8636), .Y(n5780) );
  CLKMX2X2 U4939 ( .A(hd_a08[3]), .B(d08[3]), .S0(n8636), .Y(n5779) );
  CLKMX2X2 U4940 ( .A(hd_a08[2]), .B(d08[2]), .S0(n8646), .Y(n5778) );
  CLKMX2X2 U4941 ( .A(hd_a08[1]), .B(d08[1]), .S0(n8636), .Y(n5777) );
  CLKMX2X2 U4942 ( .A(hd_a08[0]), .B(d08[0]), .S0(n8636), .Y(n5776) );
  CLKMX2X2 U4943 ( .A(hd_a09[35]), .B(d09[35]), .S0(n8636), .Y(n5775) );
  CLKMX2X2 U4944 ( .A(hd_a09[34]), .B(d09[34]), .S0(n8636), .Y(n5774) );
  CLKMX2X2 U4945 ( .A(hd_a09[33]), .B(d09[33]), .S0(n8636), .Y(n5773) );
  CLKMX2X2 U4946 ( .A(hd_a09[32]), .B(d09[32]), .S0(n8636), .Y(n5772) );
  CLKMX2X2 U4947 ( .A(hd_a09[31]), .B(d09[31]), .S0(n8636), .Y(n5771) );
  CLKMX2X2 U4948 ( .A(hd_a09[30]), .B(d09[30]), .S0(n8641), .Y(n5770) );
  CLKMX2X2 U4949 ( .A(hd_a09[29]), .B(d09[29]), .S0(n8614), .Y(n5769) );
  CLKMX2X2 U4950 ( .A(hd_a09[28]), .B(d09[28]), .S0(n8614), .Y(n5768) );
  CLKMX2X2 U4951 ( .A(hd_a09[27]), .B(d09[27]), .S0(n8614), .Y(n5767) );
  CLKMX2X2 U4952 ( .A(hd_a09[26]), .B(d09[26]), .S0(n8614), .Y(n5766) );
  CLKMX2X2 U4953 ( .A(hd_a09[25]), .B(d09[25]), .S0(n8614), .Y(n5765) );
  CLKMX2X2 U4954 ( .A(hd_a09[24]), .B(d09[24]), .S0(n8614), .Y(n5764) );
  CLKMX2X2 U4955 ( .A(hd_a09[23]), .B(d09[23]), .S0(n8614), .Y(n5763) );
  CLKMX2X2 U4956 ( .A(hd_a09[22]), .B(d09[22]), .S0(n8614), .Y(n5762) );
  CLKMX2X2 U4957 ( .A(hd_a09[21]), .B(d09[21]), .S0(n8614), .Y(n5761) );
  CLKMX2X2 U4958 ( .A(hd_a09[20]), .B(d09[20]), .S0(n8614), .Y(n5760) );
  CLKMX2X2 U4959 ( .A(hd_a09[19]), .B(d09[19]), .S0(n8613), .Y(n5759) );
  CLKMX2X2 U4960 ( .A(hd_a09[18]), .B(d09[18]), .S0(n8613), .Y(n5758) );
  CLKMX2X2 U4961 ( .A(hd_a09[17]), .B(d09[17]), .S0(n8613), .Y(n5757) );
  CLKMX2X2 U4962 ( .A(hd_a09[16]), .B(d09[16]), .S0(n8613), .Y(n5756) );
  CLKMX2X2 U4963 ( .A(hd_a09[15]), .B(d09[15]), .S0(n8613), .Y(n5755) );
  CLKMX2X2 U4964 ( .A(hd_a09[14]), .B(d09[14]), .S0(n8613), .Y(n5754) );
  CLKMX2X2 U4965 ( .A(hd_a09[13]), .B(d09[13]), .S0(n8613), .Y(n5753) );
  CLKMX2X2 U4966 ( .A(hd_a09[12]), .B(d09[12]), .S0(n8613), .Y(n5752) );
  CLKMX2X2 U4967 ( .A(hd_a09[11]), .B(d09[11]), .S0(n8613), .Y(n5751) );
  CLKMX2X2 U4968 ( .A(hd_a09[10]), .B(d09[10]), .S0(n8613), .Y(n5750) );
  CLKMX2X2 U4969 ( .A(hd_a09[9]), .B(d09[9]), .S0(n8613), .Y(n5749) );
  CLKMX2X2 U4970 ( .A(hd_a09[8]), .B(d09[8]), .S0(n8613), .Y(n5748) );
  CLKMX2X2 U4971 ( .A(hd_a09[7]), .B(d09[7]), .S0(n8613), .Y(n5747) );
  CLKMX2X2 U4972 ( .A(hd_a09[6]), .B(d09[6]), .S0(n8612), .Y(n5746) );
  CLKMX2X2 U4973 ( .A(hd_a09[5]), .B(d09[5]), .S0(n8612), .Y(n5745) );
  CLKMX2X2 U4974 ( .A(hd_a09[4]), .B(d09[4]), .S0(n8612), .Y(n5744) );
  CLKMX2X2 U4975 ( .A(hd_a09[3]), .B(d09[3]), .S0(n8612), .Y(n5743) );
  CLKMX2X2 U4976 ( .A(hd_a09[2]), .B(d09[2]), .S0(n8612), .Y(n5742) );
  CLKMX2X2 U4977 ( .A(hd_a09[1]), .B(d09[1]), .S0(n8612), .Y(n5741) );
  CLKMX2X2 U4978 ( .A(hd_a09[0]), .B(d09[0]), .S0(n8612), .Y(n5740) );
  CLKMX2X2 U4979 ( .A(hd_a10[35]), .B(d10[35]), .S0(n8612), .Y(n5739) );
  CLKMX2X2 U4980 ( .A(hd_a10[34]), .B(d10[34]), .S0(n8612), .Y(n5738) );
  CLKMX2X2 U4981 ( .A(hd_a10[33]), .B(d10[33]), .S0(n8612), .Y(n5737) );
  CLKMX2X2 U4982 ( .A(hd_a10[32]), .B(d10[32]), .S0(n8612), .Y(n5736) );
  CLKMX2X2 U4983 ( .A(hd_a10[31]), .B(d10[31]), .S0(n8612), .Y(n5735) );
  CLKMX2X2 U4984 ( .A(hd_a10[30]), .B(d10[30]), .S0(n8612), .Y(n5734) );
  CLKMX2X2 U4985 ( .A(hd_a10[29]), .B(d10[29]), .S0(n8611), .Y(n5733) );
  CLKMX2X2 U4986 ( .A(hd_a10[28]), .B(d10[28]), .S0(n8611), .Y(n5732) );
  CLKMX2X2 U4987 ( .A(hd_a10[27]), .B(d10[27]), .S0(n8611), .Y(n5731) );
  CLKMX2X2 U4988 ( .A(hd_a10[26]), .B(d10[26]), .S0(n8611), .Y(n5730) );
  CLKMX2X2 U4989 ( .A(hd_a10[25]), .B(d10[25]), .S0(n8611), .Y(n5729) );
  CLKMX2X2 U4990 ( .A(hd_a10[24]), .B(d10[24]), .S0(n8611), .Y(n5728) );
  CLKMX2X2 U4991 ( .A(hd_a10[23]), .B(d10[23]), .S0(n8611), .Y(n5727) );
  CLKMX2X2 U4992 ( .A(hd_a10[22]), .B(d10[22]), .S0(n8611), .Y(n5726) );
  CLKMX2X2 U4993 ( .A(hd_a10[21]), .B(d10[21]), .S0(n8611), .Y(n5725) );
  CLKMX2X2 U4994 ( .A(hd_a10[20]), .B(d10[20]), .S0(n8611), .Y(n5724) );
  CLKMX2X2 U4995 ( .A(hd_a10[19]), .B(d10[19]), .S0(n8611), .Y(n5723) );
  CLKMX2X2 U4996 ( .A(hd_a10[18]), .B(d10[18]), .S0(n8611), .Y(n5722) );
  CLKMX2X2 U4997 ( .A(hd_a10[17]), .B(d10[17]), .S0(n8611), .Y(n5721) );
  CLKMX2X2 U4998 ( .A(hd_a10[16]), .B(d10[16]), .S0(n8610), .Y(n5720) );
  CLKMX2X2 U4999 ( .A(hd_a10[15]), .B(d10[15]), .S0(n8610), .Y(n5719) );
  CLKMX2X2 U5000 ( .A(hd_a10[14]), .B(d10[14]), .S0(n8610), .Y(n5718) );
  CLKMX2X2 U5001 ( .A(hd_a10[13]), .B(d10[13]), .S0(n8610), .Y(n5717) );
  CLKMX2X2 U5002 ( .A(hd_a10[12]), .B(d10[12]), .S0(n8610), .Y(n5716) );
  CLKMX2X2 U5003 ( .A(hd_a10[11]), .B(d10[11]), .S0(n8610), .Y(n5715) );
  CLKMX2X2 U5004 ( .A(hd_a10[10]), .B(d10[10]), .S0(n8610), .Y(n5714) );
  CLKMX2X2 U5005 ( .A(hd_a10[9]), .B(d10[9]), .S0(n8610), .Y(n5713) );
  CLKMX2X2 U5006 ( .A(hd_a10[8]), .B(d10[8]), .S0(n8610), .Y(n5712) );
  CLKMX2X2 U5007 ( .A(hd_a10[7]), .B(d10[7]), .S0(n8610), .Y(n5711) );
  CLKMX2X2 U5008 ( .A(hd_a10[6]), .B(d10[6]), .S0(n8610), .Y(n5710) );
  CLKMX2X2 U5009 ( .A(hd_a10[5]), .B(d10[5]), .S0(n8610), .Y(n5709) );
  CLKMX2X2 U5010 ( .A(hd_a10[4]), .B(d10[4]), .S0(n8610), .Y(n5708) );
  CLKMX2X2 U5011 ( .A(hd_a10[3]), .B(d10[3]), .S0(n8609), .Y(n5707) );
  CLKMX2X2 U5012 ( .A(hd_a10[2]), .B(d10[2]), .S0(n8609), .Y(n5706) );
  CLKMX2X2 U5013 ( .A(hd_a10[1]), .B(d10[1]), .S0(n8609), .Y(n5705) );
  CLKMX2X2 U5014 ( .A(hd_a10[0]), .B(d10[0]), .S0(n8609), .Y(n5704) );
  CLKMX2X2 U5015 ( .A(hd_a11[35]), .B(d11[35]), .S0(n8609), .Y(n5703) );
  CLKMX2X2 U5016 ( .A(hd_a11[34]), .B(d11[34]), .S0(n8609), .Y(n5702) );
  CLKMX2X2 U5017 ( .A(hd_a11[33]), .B(d11[33]), .S0(n8609), .Y(n5701) );
  CLKMX2X2 U5018 ( .A(hd_a11[32]), .B(d11[32]), .S0(n8609), .Y(n5700) );
  CLKMX2X2 U5019 ( .A(hd_a11[31]), .B(d11[31]), .S0(n8609), .Y(n5699) );
  CLKMX2X2 U5020 ( .A(hd_a11[30]), .B(d11[30]), .S0(n8609), .Y(n5698) );
  CLKMX2X2 U5021 ( .A(hd_a11[29]), .B(d11[29]), .S0(n8609), .Y(n5697) );
  CLKMX2X2 U5022 ( .A(hd_a11[28]), .B(d11[28]), .S0(n8609), .Y(n5696) );
  CLKMX2X2 U5023 ( .A(hd_a11[27]), .B(d11[27]), .S0(n8608), .Y(n5695) );
  CLKMX2X2 U5024 ( .A(hd_a11[26]), .B(d11[26]), .S0(n8608), .Y(n5694) );
  CLKMX2X2 U5025 ( .A(hd_a11[25]), .B(d11[25]), .S0(n8608), .Y(n5693) );
  CLKMX2X2 U5026 ( .A(hd_a11[24]), .B(d11[24]), .S0(n8608), .Y(n5692) );
  CLKMX2X2 U5027 ( .A(hd_a11[23]), .B(d11[23]), .S0(n8608), .Y(n5691) );
  CLKMX2X2 U5028 ( .A(hd_a11[22]), .B(d11[22]), .S0(n8608), .Y(n5690) );
  CLKMX2X2 U5029 ( .A(hd_a11[21]), .B(d11[21]), .S0(n8608), .Y(n5689) );
  CLKMX2X2 U5030 ( .A(hd_a11[20]), .B(d11[20]), .S0(n8608), .Y(n5688) );
  CLKMX2X2 U5031 ( .A(hd_a11[19]), .B(d11[19]), .S0(n8608), .Y(n5687) );
  CLKMX2X2 U5032 ( .A(hd_a11[18]), .B(d11[18]), .S0(n8608), .Y(n5686) );
  CLKMX2X2 U5033 ( .A(hd_a11[17]), .B(d11[17]), .S0(n8608), .Y(n5685) );
  CLKMX2X2 U5034 ( .A(hd_a11[16]), .B(d11[16]), .S0(n8608), .Y(n5684) );
  CLKMX2X2 U5035 ( .A(hd_a11[15]), .B(d11[15]), .S0(n8608), .Y(n5683) );
  CLKMX2X2 U5036 ( .A(hd_a11[14]), .B(d11[14]), .S0(n8607), .Y(n5682) );
  CLKMX2X2 U5037 ( .A(hd_a11[13]), .B(d11[13]), .S0(n8607), .Y(n5681) );
  CLKMX2X2 U5038 ( .A(hd_a11[12]), .B(d11[12]), .S0(n8607), .Y(n5680) );
  CLKMX2X2 U5039 ( .A(hd_a11[11]), .B(d11[11]), .S0(n8607), .Y(n5679) );
  CLKMX2X2 U5040 ( .A(hd_a11[10]), .B(d11[10]), .S0(n8607), .Y(n5678) );
  CLKMX2X2 U5041 ( .A(hd_a11[9]), .B(d11[9]), .S0(n8607), .Y(n5677) );
  CLKMX2X2 U5042 ( .A(hd_a11[8]), .B(d11[8]), .S0(n8607), .Y(n5676) );
  CLKMX2X2 U5043 ( .A(hd_a11[7]), .B(d11[7]), .S0(n8607), .Y(n5675) );
  CLKMX2X2 U5044 ( .A(hd_a11[6]), .B(d11[6]), .S0(n8607), .Y(n5674) );
  CLKMX2X2 U5045 ( .A(hd_a11[5]), .B(d11[5]), .S0(n8607), .Y(n5673) );
  CLKMX2X2 U5046 ( .A(hd_a11[4]), .B(d11[4]), .S0(n8607), .Y(n5672) );
  CLKMX2X2 U5047 ( .A(hd_a11[3]), .B(d11[3]), .S0(n8607), .Y(n5671) );
  CLKMX2X2 U5048 ( .A(hd_a11[2]), .B(d11[2]), .S0(n8607), .Y(n5670) );
  CLKMX2X2 U5049 ( .A(hd_a11[1]), .B(d11[1]), .S0(n8606), .Y(n5669) );
  CLKMX2X2 U5050 ( .A(hd_a11[0]), .B(d11[0]), .S0(n8606), .Y(n5668) );
  CLKMX2X2 U5051 ( .A(hd_a12[35]), .B(d12[35]), .S0(n8606), .Y(n5667) );
  CLKMX2X2 U5052 ( .A(hd_a12[34]), .B(d12[34]), .S0(n8606), .Y(n5666) );
  CLKMX2X2 U5053 ( .A(hd_a12[33]), .B(d12[33]), .S0(n8606), .Y(n5665) );
  CLKMX2X2 U5054 ( .A(hd_a12[32]), .B(d12[32]), .S0(n8606), .Y(n5664) );
  CLKMX2X2 U5055 ( .A(hd_a12[31]), .B(d12[31]), .S0(n8606), .Y(n5663) );
  CLKMX2X2 U5056 ( .A(hd_a12[30]), .B(d12[30]), .S0(n8606), .Y(n5662) );
  CLKMX2X2 U5057 ( .A(hd_a12[29]), .B(d12[29]), .S0(n8606), .Y(n5661) );
  CLKMX2X2 U5058 ( .A(hd_a12[28]), .B(d12[28]), .S0(n8606), .Y(n5660) );
  CLKMX2X2 U5059 ( .A(hd_a12[27]), .B(d12[27]), .S0(n8606), .Y(n5659) );
  CLKMX2X2 U5060 ( .A(hd_a12[26]), .B(d12[26]), .S0(n8606), .Y(n5658) );
  CLKMX2X2 U5061 ( .A(hd_a12[25]), .B(d12[25]), .S0(n8606), .Y(n5657) );
  CLKMX2X2 U5062 ( .A(hd_a12[24]), .B(d12[24]), .S0(n8605), .Y(n5656) );
  CLKMX2X2 U5063 ( .A(hd_a12[23]), .B(d12[23]), .S0(n8605), .Y(n5655) );
  CLKMX2X2 U5064 ( .A(hd_a12[22]), .B(d12[22]), .S0(n8605), .Y(n5654) );
  CLKMX2X2 U5065 ( .A(hd_a12[21]), .B(d12[21]), .S0(n8605), .Y(n5653) );
  CLKMX2X2 U5066 ( .A(hd_a12[20]), .B(d12[20]), .S0(n8605), .Y(n5652) );
  CLKMX2X2 U5067 ( .A(hd_a12[19]), .B(d12[19]), .S0(n8605), .Y(n5651) );
  CLKMX2X2 U5068 ( .A(hd_a12[18]), .B(d12[18]), .S0(n8605), .Y(n5650) );
  CLKMX2X2 U5069 ( .A(hd_a12[17]), .B(d12[17]), .S0(n8605), .Y(n5649) );
  CLKMX2X2 U5070 ( .A(hd_a12[16]), .B(d12[16]), .S0(n8605), .Y(n5648) );
  CLKMX2X2 U5071 ( .A(hd_a12[15]), .B(d12[15]), .S0(n8605), .Y(n5647) );
  CLKMX2X2 U5072 ( .A(hd_a12[14]), .B(d12[14]), .S0(n8605), .Y(n5646) );
  CLKMX2X2 U5073 ( .A(hd_a12[13]), .B(d12[13]), .S0(n8605), .Y(n5645) );
  CLKMX2X2 U5074 ( .A(hd_a12[12]), .B(d12[12]), .S0(n8605), .Y(n5644) );
  CLKMX2X2 U5075 ( .A(hd_a12[11]), .B(d12[11]), .S0(n8604), .Y(n5643) );
  CLKMX2X2 U5076 ( .A(hd_a12[10]), .B(d12[10]), .S0(n8604), .Y(n5642) );
  CLKMX2X2 U5077 ( .A(hd_a12[9]), .B(d12[9]), .S0(n8604), .Y(n5641) );
  CLKMX2X2 U5078 ( .A(hd_a12[8]), .B(d12[8]), .S0(n8604), .Y(n5640) );
  CLKMX2X2 U5079 ( .A(hd_a12[7]), .B(d12[7]), .S0(n8604), .Y(n5639) );
  CLKMX2X2 U5080 ( .A(hd_a12[6]), .B(d12[6]), .S0(n8604), .Y(n5638) );
  CLKMX2X2 U5081 ( .A(hd_a12[5]), .B(d12[5]), .S0(n8604), .Y(n5637) );
  CLKMX2X2 U5082 ( .A(hd_a12[4]), .B(d12[4]), .S0(n8604), .Y(n5636) );
  CLKMX2X2 U5083 ( .A(hd_a12[3]), .B(d12[3]), .S0(n8604), .Y(n5635) );
  CLKMX2X2 U5084 ( .A(hd_a12[2]), .B(d12[2]), .S0(n8604), .Y(n5634) );
  CLKMX2X2 U5085 ( .A(hd_a12[1]), .B(d12[1]), .S0(n8604), .Y(n5633) );
  CLKMX2X2 U5086 ( .A(hd_a12[0]), .B(d12[0]), .S0(n8604), .Y(n5632) );
  CLKMX2X2 U5087 ( .A(hd_a13[35]), .B(d13[35]), .S0(n8609), .Y(n5631) );
  CLKMX2X2 U5088 ( .A(hd_a13[34]), .B(d13[34]), .S0(n8625), .Y(n5630) );
  CLKMX2X2 U5089 ( .A(hd_a13[33]), .B(d13[33]), .S0(n8625), .Y(n5629) );
  CLKMX2X2 U5090 ( .A(hd_a13[32]), .B(d13[32]), .S0(n8625), .Y(n5628) );
  CLKMX2X2 U5091 ( .A(hd_a13[31]), .B(d13[31]), .S0(n8625), .Y(n5627) );
  CLKMX2X2 U5092 ( .A(hd_a13[30]), .B(d13[30]), .S0(n8625), .Y(n5626) );
  CLKMX2X2 U5093 ( .A(hd_a13[29]), .B(d13[29]), .S0(n8624), .Y(n5625) );
  CLKMX2X2 U5094 ( .A(hd_a13[28]), .B(d13[28]), .S0(n8624), .Y(n5624) );
  CLKMX2X2 U5095 ( .A(hd_a13[27]), .B(d13[27]), .S0(n8624), .Y(n5623) );
  CLKMX2X2 U5096 ( .A(hd_a13[26]), .B(d13[26]), .S0(n8624), .Y(n5622) );
  CLKMX2X2 U5097 ( .A(hd_a13[25]), .B(d13[25]), .S0(n8624), .Y(n5621) );
  CLKMX2X2 U5098 ( .A(hd_a13[24]), .B(d13[24]), .S0(n8624), .Y(n5620) );
  CLKMX2X2 U5099 ( .A(hd_a13[23]), .B(d13[23]), .S0(n8624), .Y(n5619) );
  CLKMX2X2 U5100 ( .A(hd_a13[22]), .B(d13[22]), .S0(n8624), .Y(n5618) );
  CLKMX2X2 U5101 ( .A(hd_a13[21]), .B(d13[21]), .S0(n8624), .Y(n5617) );
  CLKMX2X2 U5102 ( .A(hd_a13[20]), .B(d13[20]), .S0(n8624), .Y(n5616) );
  CLKMX2X2 U5103 ( .A(hd_a13[19]), .B(d13[19]), .S0(n8624), .Y(n5615) );
  CLKMX2X2 U5104 ( .A(hd_a13[18]), .B(d13[18]), .S0(n8624), .Y(n5614) );
  CLKMX2X2 U5105 ( .A(hd_a13[17]), .B(d13[17]), .S0(n8624), .Y(n5613) );
  CLKMX2X2 U5106 ( .A(hd_a13[16]), .B(d13[16]), .S0(n8623), .Y(n5612) );
  CLKMX2X2 U5107 ( .A(hd_a13[15]), .B(d13[15]), .S0(n8623), .Y(n5611) );
  CLKMX2X2 U5108 ( .A(hd_a13[14]), .B(d13[14]), .S0(n8623), .Y(n5610) );
  CLKMX2X2 U5109 ( .A(hd_a13[13]), .B(d13[13]), .S0(n8623), .Y(n5609) );
  CLKMX2X2 U5110 ( .A(hd_a13[12]), .B(d13[12]), .S0(n8623), .Y(n5608) );
  CLKMX2X2 U5111 ( .A(hd_a13[11]), .B(d13[11]), .S0(n8623), .Y(n5607) );
  CLKMX2X2 U5112 ( .A(hd_a13[10]), .B(d13[10]), .S0(n8623), .Y(n5606) );
  CLKMX2X2 U5113 ( .A(hd_a13[9]), .B(d13[9]), .S0(n8623), .Y(n5605) );
  CLKMX2X2 U5114 ( .A(hd_a13[8]), .B(d13[8]), .S0(n8623), .Y(n5604) );
  CLKMX2X2 U5115 ( .A(hd_a13[7]), .B(d13[7]), .S0(n8623), .Y(n5603) );
  CLKMX2X2 U5116 ( .A(hd_a13[6]), .B(d13[6]), .S0(n8623), .Y(n5602) );
  CLKMX2X2 U5117 ( .A(hd_a13[5]), .B(d13[5]), .S0(n8623), .Y(n5601) );
  CLKMX2X2 U5118 ( .A(hd_a13[4]), .B(d13[4]), .S0(n8623), .Y(n5600) );
  CLKMX2X2 U5119 ( .A(hd_a13[3]), .B(d13[3]), .S0(n8622), .Y(n5599) );
  CLKMX2X2 U5120 ( .A(hd_a13[2]), .B(d13[2]), .S0(n8622), .Y(n5598) );
  CLKMX2X2 U5121 ( .A(hd_a13[1]), .B(d13[1]), .S0(n8622), .Y(n5597) );
  CLKMX2X2 U5122 ( .A(hd_a13[0]), .B(d13[0]), .S0(n8622), .Y(n5596) );
  CLKMX2X2 U5123 ( .A(hd_a14[35]), .B(d14[35]), .S0(n8622), .Y(n5595) );
  CLKMX2X2 U5124 ( .A(hd_a14[34]), .B(d14[34]), .S0(n8622), .Y(n5594) );
  CLKMX2X2 U5125 ( .A(hd_a14[33]), .B(d14[33]), .S0(n8622), .Y(n5593) );
  CLKMX2X2 U5126 ( .A(hd_a14[32]), .B(d14[32]), .S0(n8622), .Y(n5592) );
  CLKMX2X2 U5127 ( .A(hd_a14[31]), .B(d14[31]), .S0(n8622), .Y(n5591) );
  CLKMX2X2 U5128 ( .A(hd_a14[30]), .B(d14[30]), .S0(n8622), .Y(n5590) );
  CLKMX2X2 U5129 ( .A(hd_a14[29]), .B(d14[29]), .S0(n8622), .Y(n5589) );
  CLKMX2X2 U5130 ( .A(hd_a14[28]), .B(d14[28]), .S0(n8622), .Y(n5588) );
  CLKMX2X2 U5131 ( .A(hd_a14[27]), .B(d14[27]), .S0(n8622), .Y(n5587) );
  CLKMX2X2 U5132 ( .A(hd_a14[26]), .B(d14[26]), .S0(n8621), .Y(n5586) );
  CLKMX2X2 U5133 ( .A(hd_a14[25]), .B(d14[25]), .S0(n8621), .Y(n5585) );
  CLKMX2X2 U5134 ( .A(hd_a14[24]), .B(d14[24]), .S0(n8621), .Y(n5584) );
  CLKMX2X2 U5135 ( .A(hd_a14[23]), .B(d14[23]), .S0(n8621), .Y(n5583) );
  CLKMX2X2 U5136 ( .A(hd_a14[22]), .B(d14[22]), .S0(n8621), .Y(n5582) );
  CLKMX2X2 U5137 ( .A(hd_a14[21]), .B(d14[21]), .S0(n8621), .Y(n5581) );
  CLKMX2X2 U5138 ( .A(hd_a14[20]), .B(d14[20]), .S0(n8621), .Y(n5580) );
  CLKMX2X2 U5139 ( .A(hd_a14[19]), .B(d14[19]), .S0(n8621), .Y(n5579) );
  CLKMX2X2 U5140 ( .A(hd_a14[18]), .B(d14[18]), .S0(n8621), .Y(n5578) );
  CLKMX2X2 U5141 ( .A(hd_a14[17]), .B(d14[17]), .S0(n8621), .Y(n5577) );
  CLKMX2X2 U5142 ( .A(hd_a14[16]), .B(d14[16]), .S0(n8621), .Y(n5576) );
  CLKMX2X2 U5143 ( .A(hd_a14[15]), .B(d14[15]), .S0(n8621), .Y(n5575) );
  CLKMX2X2 U5144 ( .A(hd_a14[14]), .B(d14[14]), .S0(n8621), .Y(n5574) );
  CLKMX2X2 U5145 ( .A(hd_a14[13]), .B(d14[13]), .S0(n8620), .Y(n5573) );
  CLKMX2X2 U5146 ( .A(hd_a14[12]), .B(d14[12]), .S0(n8620), .Y(n5572) );
  CLKMX2X2 U5147 ( .A(hd_a14[11]), .B(d14[11]), .S0(n8620), .Y(n5571) );
  CLKMX2X2 U5148 ( .A(hd_a14[10]), .B(d14[10]), .S0(n8620), .Y(n5570) );
  CLKMX2X2 U5149 ( .A(hd_a14[9]), .B(d14[9]), .S0(n8620), .Y(n5569) );
  CLKMX2X2 U5150 ( .A(hd_a14[8]), .B(d14[8]), .S0(n8620), .Y(n5568) );
  CLKMX2X2 U5151 ( .A(hd_a14[7]), .B(d14[7]), .S0(n8620), .Y(n5567) );
  CLKMX2X2 U5152 ( .A(hd_a14[6]), .B(d14[6]), .S0(n8620), .Y(n5566) );
  CLKMX2X2 U5153 ( .A(hd_a14[5]), .B(d14[5]), .S0(n8620), .Y(n5565) );
  CLKMX2X2 U5154 ( .A(hd_a14[4]), .B(d14[4]), .S0(n8620), .Y(n5564) );
  CLKMX2X2 U5155 ( .A(hd_a14[3]), .B(d14[3]), .S0(n8620), .Y(n5563) );
  CLKMX2X2 U5156 ( .A(hd_a14[2]), .B(d14[2]), .S0(n8620), .Y(n5562) );
  CLKMX2X2 U5157 ( .A(hd_a14[1]), .B(d14[1]), .S0(n8619), .Y(n5561) );
  CLKMX2X2 U5158 ( .A(hd_a14[0]), .B(d14[0]), .S0(n8619), .Y(n5560) );
  CLKMX2X2 U5159 ( .A(hd_a15[35]), .B(d15[35]), .S0(n8619), .Y(n5559) );
  CLKMX2X2 U5160 ( .A(hd_a15[34]), .B(d15[34]), .S0(n8619), .Y(n5558) );
  CLKMX2X2 U5161 ( .A(hd_a15[33]), .B(d15[33]), .S0(n8619), .Y(n5557) );
  CLKMX2X2 U5162 ( .A(hd_a15[32]), .B(d15[32]), .S0(n8619), .Y(n5556) );
  CLKMX2X2 U5163 ( .A(hd_a15[31]), .B(d15[31]), .S0(n8619), .Y(n5555) );
  CLKMX2X2 U5164 ( .A(hd_a15[30]), .B(d15[30]), .S0(n8619), .Y(n5554) );
  CLKMX2X2 U5165 ( .A(hd_a15[29]), .B(d15[29]), .S0(n8619), .Y(n5553) );
  CLKMX2X2 U5166 ( .A(hd_a15[28]), .B(d15[28]), .S0(n8619), .Y(n5552) );
  CLKMX2X2 U5167 ( .A(hd_a15[27]), .B(d15[27]), .S0(n8619), .Y(n5551) );
  CLKMX2X2 U5168 ( .A(hd_a15[26]), .B(d15[26]), .S0(n8619), .Y(n5550) );
  CLKMX2X2 U5169 ( .A(hd_a15[25]), .B(d15[25]), .S0(n8619), .Y(n5549) );
  CLKMX2X2 U5170 ( .A(hd_a15[24]), .B(d15[24]), .S0(n8618), .Y(n5548) );
  CLKMX2X2 U5171 ( .A(hd_a15[23]), .B(d15[23]), .S0(n8618), .Y(n5547) );
  CLKMX2X2 U5172 ( .A(hd_a15[22]), .B(d15[22]), .S0(n8618), .Y(n5546) );
  CLKMX2X2 U5173 ( .A(hd_a15[21]), .B(d15[21]), .S0(n8618), .Y(n5545) );
  CLKMX2X2 U5174 ( .A(hd_a15[20]), .B(d15[20]), .S0(n8618), .Y(n5544) );
  CLKMX2X2 U5175 ( .A(hd_a15[19]), .B(d15[19]), .S0(n8618), .Y(n5543) );
  CLKMX2X2 U5176 ( .A(hd_a15[18]), .B(d15[18]), .S0(n8618), .Y(n5542) );
  CLKMX2X2 U5177 ( .A(hd_a15[17]), .B(d15[17]), .S0(n8618), .Y(n5541) );
  CLKMX2X2 U5178 ( .A(hd_a15[16]), .B(d15[16]), .S0(n8618), .Y(n5540) );
  CLKMX2X2 U5179 ( .A(hd_a15[15]), .B(d15[15]), .S0(n8618), .Y(n5539) );
  CLKMX2X2 U5180 ( .A(hd_a15[14]), .B(d15[14]), .S0(n8618), .Y(n5538) );
  CLKMX2X2 U5181 ( .A(hd_a15[13]), .B(d15[13]), .S0(n8618), .Y(n5537) );
  CLKMX2X2 U5182 ( .A(hd_a15[12]), .B(d15[12]), .S0(n8618), .Y(n5536) );
  CLKMX2X2 U5183 ( .A(hd_a15[11]), .B(d15[11]), .S0(n8617), .Y(n5535) );
  CLKMX2X2 U5184 ( .A(hd_a15[10]), .B(d15[10]), .S0(n8617), .Y(n5534) );
  CLKMX2X2 U5185 ( .A(hd_a15[9]), .B(d15[9]), .S0(n8617), .Y(n5533) );
  CLKMX2X2 U5186 ( .A(hd_a15[8]), .B(d15[8]), .S0(n8617), .Y(n5532) );
  CLKMX2X2 U5187 ( .A(hd_a15[7]), .B(d15[7]), .S0(n8617), .Y(n5531) );
  CLKMX2X2 U5188 ( .A(hd_a15[6]), .B(d15[6]), .S0(n8617), .Y(n5530) );
  CLKMX2X2 U5189 ( .A(hd_a15[5]), .B(d15[5]), .S0(n8617), .Y(n5529) );
  CLKMX2X2 U5190 ( .A(hd_a15[4]), .B(d15[4]), .S0(n8617), .Y(n5528) );
  CLKMX2X2 U5191 ( .A(hd_a15[3]), .B(d15[3]), .S0(n8617), .Y(n5527) );
  CLKMX2X2 U5192 ( .A(hd_a15[2]), .B(d15[2]), .S0(n8617), .Y(n5526) );
  CLKMX2X2 U5193 ( .A(hd_a15[1]), .B(d15[1]), .S0(n8617), .Y(n5525) );
  CLKMX2X2 U5194 ( .A(hd_a15[0]), .B(d15[0]), .S0(n8617), .Y(n5524) );
  CLKMX2X2 U5195 ( .A(hd_a16[35]), .B(d16[35]), .S0(n8617), .Y(n5523) );
  CLKMX2X2 U5196 ( .A(hd_a16[34]), .B(d16[34]), .S0(n8616), .Y(n5522) );
  CLKMX2X2 U5197 ( .A(hd_a16[33]), .B(d16[33]), .S0(n8616), .Y(n5521) );
  CLKMX2X2 U5198 ( .A(hd_a16[32]), .B(d16[32]), .S0(n8616), .Y(n5520) );
  CLKMX2X2 U5199 ( .A(hd_a16[31]), .B(d16[31]), .S0(n8616), .Y(n5519) );
  CLKMX2X2 U5200 ( .A(hd_a16[30]), .B(d16[30]), .S0(n8616), .Y(n5518) );
  CLKMX2X2 U5201 ( .A(hd_a16[29]), .B(d16[29]), .S0(n8616), .Y(n5517) );
  CLKMX2X2 U5202 ( .A(hd_a16[28]), .B(d16[28]), .S0(n8616), .Y(n5516) );
  CLKMX2X2 U5203 ( .A(hd_a16[27]), .B(d16[27]), .S0(n8616), .Y(n5515) );
  CLKMX2X2 U5204 ( .A(hd_a16[26]), .B(d16[26]), .S0(n8616), .Y(n5514) );
  CLKMX2X2 U5205 ( .A(hd_a16[25]), .B(d16[25]), .S0(n8616), .Y(n5513) );
  CLKMX2X2 U5206 ( .A(hd_a16[24]), .B(d16[24]), .S0(n8616), .Y(n5512) );
  CLKMX2X2 U5207 ( .A(hd_a16[23]), .B(d16[23]), .S0(n8616), .Y(n5511) );
  CLKMX2X2 U5208 ( .A(hd_a16[22]), .B(d16[22]), .S0(n8616), .Y(n5510) );
  CLKMX2X2 U5209 ( .A(hd_a16[21]), .B(d16[21]), .S0(n8615), .Y(n5509) );
  CLKMX2X2 U5210 ( .A(hd_a16[20]), .B(d16[20]), .S0(n8615), .Y(n5508) );
  CLKMX2X2 U5211 ( .A(hd_a16[19]), .B(d16[19]), .S0(n8615), .Y(n5507) );
  CLKMX2X2 U5212 ( .A(hd_a16[18]), .B(d16[18]), .S0(n8615), .Y(n5506) );
  CLKMX2X2 U5213 ( .A(hd_a16[17]), .B(d16[17]), .S0(n8615), .Y(n5505) );
  CLKMX2X2 U5214 ( .A(hd_a16[16]), .B(d16[16]), .S0(n8615), .Y(n5504) );
  CLKMX2X2 U5215 ( .A(hd_a16[15]), .B(d16[15]), .S0(n8615), .Y(n5503) );
  CLKMX2X2 U5216 ( .A(hd_a16[14]), .B(d16[14]), .S0(n8615), .Y(n5502) );
  CLKMX2X2 U5217 ( .A(hd_a16[13]), .B(d16[13]), .S0(n8615), .Y(n5501) );
  CLKMX2X2 U5218 ( .A(hd_a16[12]), .B(d16[12]), .S0(n8615), .Y(n5500) );
  CLKMX2X2 U5219 ( .A(hd_a16[11]), .B(d16[11]), .S0(n8615), .Y(n5499) );
  CLKMX2X2 U5220 ( .A(hd_a16[10]), .B(d16[10]), .S0(n8615), .Y(n5498) );
  CLKMX2X2 U5221 ( .A(hd_a16[9]), .B(d16[9]), .S0(n8615), .Y(n5497) );
  CLKMX2X2 U5222 ( .A(hd_a16[8]), .B(d16[8]), .S0(n8614), .Y(n5496) );
  CLKMX2X2 U5223 ( .A(hd_a16[7]), .B(d16[7]), .S0(n8614), .Y(n5495) );
  CLKMX2X2 U5224 ( .A(hd_a16[6]), .B(d16[6]), .S0(n8614), .Y(n5494) );
  CLKMX2X2 U5225 ( .A(hd_a16[5]), .B(d16[5]), .S0(n8620), .Y(n5493) );
  CLKMX2X2 U5226 ( .A(hd_a16[4]), .B(d16[4]), .S0(n8625), .Y(n5492) );
  CLKMX2X2 U5227 ( .A(hd_a16[3]), .B(d16[3]), .S0(n8679), .Y(n5491) );
  CLKMX2X2 U5228 ( .A(hd_a16[2]), .B(d16[2]), .S0(n8678), .Y(n5490) );
  CLKMX2X2 U5229 ( .A(hd_a16[1]), .B(d16[1]), .S0(n8678), .Y(n5489) );
  CLKMX2X2 U5230 ( .A(hd_a16[0]), .B(d16[0]), .S0(n8678), .Y(n5488) );
  CLKMX2X2 U5231 ( .A(hd_a17[35]), .B(d17[35]), .S0(n8678), .Y(n5487) );
  CLKMX2X2 U5232 ( .A(hd_a17[34]), .B(d17[34]), .S0(n8678), .Y(n5486) );
  CLKMX2X2 U5233 ( .A(hd_a17[33]), .B(d17[33]), .S0(n8678), .Y(n5485) );
  CLKMX2X2 U5234 ( .A(hd_a17[32]), .B(d17[32]), .S0(n8678), .Y(n5484) );
  CLKMX2X2 U5235 ( .A(hd_a17[31]), .B(d17[31]), .S0(n8678), .Y(n5483) );
  CLKMX2X2 U5236 ( .A(hd_a17[30]), .B(d17[30]), .S0(n8678), .Y(n5482) );
  CLKMX2X2 U5237 ( .A(hd_a17[29]), .B(d17[29]), .S0(n8678), .Y(n5481) );
  CLKMX2X2 U5238 ( .A(hd_a17[28]), .B(d17[28]), .S0(n8678), .Y(n5480) );
  CLKMX2X2 U5239 ( .A(hd_a17[27]), .B(d17[27]), .S0(n8678), .Y(n5479) );
  CLKMX2X2 U5240 ( .A(hd_a17[26]), .B(d17[26]), .S0(n8678), .Y(n5478) );
  CLKMX2X2 U5241 ( .A(hd_a17[25]), .B(d17[25]), .S0(n8677), .Y(n5477) );
  CLKMX2X2 U5242 ( .A(hd_a17[24]), .B(d17[24]), .S0(n8677), .Y(n5476) );
  CLKMX2X2 U5243 ( .A(hd_a17[23]), .B(d17[23]), .S0(n8677), .Y(n5475) );
  CLKMX2X2 U5244 ( .A(hd_a17[22]), .B(d17[22]), .S0(n8677), .Y(n5474) );
  CLKMX2X2 U5245 ( .A(hd_a17[21]), .B(d17[21]), .S0(n8677), .Y(n5473) );
  CLKMX2X2 U5246 ( .A(hd_a17[20]), .B(d17[20]), .S0(n8677), .Y(n5472) );
  CLKMX2X2 U5247 ( .A(hd_a17[19]), .B(d17[19]), .S0(n8677), .Y(n5471) );
  CLKMX2X2 U5248 ( .A(hd_a17[18]), .B(d17[18]), .S0(n8677), .Y(n5470) );
  CLKMX2X2 U5249 ( .A(hd_a17[17]), .B(d17[17]), .S0(n8677), .Y(n5469) );
  CLKMX2X2 U5250 ( .A(hd_a17[16]), .B(d17[16]), .S0(n8677), .Y(n5468) );
  CLKMX2X2 U5251 ( .A(hd_a17[15]), .B(d17[15]), .S0(n8677), .Y(n5467) );
  CLKMX2X2 U5252 ( .A(hd_a17[14]), .B(d17[14]), .S0(n8677), .Y(n5466) );
  CLKMX2X2 U5253 ( .A(hd_a17[13]), .B(d17[13]), .S0(n8677), .Y(n5465) );
  CLKMX2X2 U5254 ( .A(hd_a17[12]), .B(d17[12]), .S0(n8676), .Y(n5464) );
  CLKMX2X2 U5255 ( .A(hd_a17[11]), .B(d17[11]), .S0(n8676), .Y(n5463) );
  CLKMX2X2 U5256 ( .A(hd_a17[10]), .B(d17[10]), .S0(n8676), .Y(n5462) );
  CLKMX2X2 U5257 ( .A(hd_a17[9]), .B(d17[9]), .S0(n8676), .Y(n5461) );
  CLKMX2X2 U5258 ( .A(hd_a17[8]), .B(d17[8]), .S0(n8676), .Y(n5460) );
  CLKMX2X2 U5259 ( .A(hd_a17[7]), .B(d17[7]), .S0(n8676), .Y(n5459) );
  CLKMX2X2 U5260 ( .A(hd_a17[6]), .B(d17[6]), .S0(n8676), .Y(n5458) );
  CLKMX2X2 U5261 ( .A(hd_a17[5]), .B(d17[5]), .S0(n8676), .Y(n5457) );
  CLKMX2X2 U5262 ( .A(hd_a17[4]), .B(d17[4]), .S0(n8676), .Y(n5456) );
  CLKMX2X2 U5263 ( .A(hd_a17[3]), .B(d17[3]), .S0(n8676), .Y(n5455) );
  CLKMX2X2 U5264 ( .A(hd_a17[2]), .B(d17[2]), .S0(n8676), .Y(n5454) );
  CLKMX2X2 U5265 ( .A(hd_a17[1]), .B(d17[1]), .S0(n8676), .Y(n5453) );
  CLKMX2X2 U5266 ( .A(hd_a17[0]), .B(d17[0]), .S0(n8676), .Y(n5452) );
  CLKMX2X2 U5267 ( .A(hd_a18[35]), .B(d18[35]), .S0(n8675), .Y(n5451) );
  CLKMX2X2 U5268 ( .A(hd_a18[34]), .B(d18[34]), .S0(n8675), .Y(n5450) );
  CLKMX2X2 U5269 ( .A(hd_a18[33]), .B(d18[33]), .S0(n8675), .Y(n5449) );
  CLKMX2X2 U5270 ( .A(hd_a18[32]), .B(d18[32]), .S0(n8675), .Y(n5448) );
  CLKMX2X2 U5271 ( .A(hd_a18[31]), .B(d18[31]), .S0(n8675), .Y(n5447) );
  CLKMX2X2 U5272 ( .A(hd_a18[30]), .B(d18[30]), .S0(n8675), .Y(n5446) );
  CLKMX2X2 U5273 ( .A(hd_a18[29]), .B(d18[29]), .S0(n8675), .Y(n5445) );
  CLKMX2X2 U5274 ( .A(hd_a18[28]), .B(d18[28]), .S0(n8675), .Y(n5444) );
  CLKMX2X2 U5275 ( .A(hd_a18[27]), .B(d18[27]), .S0(n8675), .Y(n5443) );
  CLKMX2X2 U5276 ( .A(hd_a18[26]), .B(d18[26]), .S0(n8675), .Y(n5442) );
  CLKMX2X2 U5277 ( .A(hd_a18[25]), .B(d18[25]), .S0(n8675), .Y(n5441) );
  CLKMX2X2 U5278 ( .A(hd_a18[24]), .B(d18[24]), .S0(n8675), .Y(n5440) );
  CLKMX2X2 U5279 ( .A(hd_a18[23]), .B(d18[23]), .S0(n8675), .Y(n5439) );
  CLKMX2X2 U5280 ( .A(hd_a18[22]), .B(d18[22]), .S0(n8674), .Y(n5438) );
  CLKMX2X2 U5281 ( .A(hd_a18[21]), .B(d18[21]), .S0(n8674), .Y(n5437) );
  CLKMX2X2 U5282 ( .A(hd_a18[20]), .B(d18[20]), .S0(n8674), .Y(n5436) );
  CLKMX2X2 U5283 ( .A(hd_a18[19]), .B(d18[19]), .S0(n8674), .Y(n5435) );
  CLKMX2X2 U5284 ( .A(hd_a18[18]), .B(d18[18]), .S0(n8674), .Y(n5434) );
  CLKMX2X2 U5285 ( .A(hd_a18[17]), .B(d18[17]), .S0(n8674), .Y(n5433) );
  CLKMX2X2 U5286 ( .A(hd_a18[16]), .B(d18[16]), .S0(n8674), .Y(n5432) );
  CLKMX2X2 U5287 ( .A(hd_a18[15]), .B(d18[15]), .S0(n8674), .Y(n5431) );
  CLKMX2X2 U5288 ( .A(hd_a18[14]), .B(d18[14]), .S0(n8674), .Y(n5430) );
  CLKMX2X2 U5289 ( .A(hd_a18[13]), .B(d18[13]), .S0(n8674), .Y(n5429) );
  CLKMX2X2 U5290 ( .A(hd_a18[12]), .B(d18[12]), .S0(n8674), .Y(n5428) );
  CLKMX2X2 U5291 ( .A(hd_a18[11]), .B(d18[11]), .S0(n8674), .Y(n5427) );
  CLKMX2X2 U5292 ( .A(hd_a18[10]), .B(d18[10]), .S0(n8674), .Y(n5426) );
  CLKMX2X2 U5293 ( .A(hd_a18[9]), .B(d18[9]), .S0(n8673), .Y(n5425) );
  CLKMX2X2 U5294 ( .A(hd_a18[8]), .B(d18[8]), .S0(n8673), .Y(n5424) );
  CLKMX2X2 U5295 ( .A(hd_a18[7]), .B(d18[7]), .S0(n8673), .Y(n5423) );
  CLKMX2X2 U5296 ( .A(hd_a18[6]), .B(d18[6]), .S0(n8673), .Y(n5422) );
  CLKMX2X2 U5297 ( .A(hd_a18[5]), .B(d18[5]), .S0(n8673), .Y(n5421) );
  CLKMX2X2 U5298 ( .A(hd_a18[4]), .B(d18[4]), .S0(n8673), .Y(n5420) );
  CLKMX2X2 U5299 ( .A(hd_a18[3]), .B(d18[3]), .S0(n8673), .Y(n5419) );
  CLKMX2X2 U5300 ( .A(hd_a18[2]), .B(d18[2]), .S0(n8673), .Y(n5418) );
  CLKMX2X2 U5301 ( .A(hd_a18[1]), .B(d18[1]), .S0(n8673), .Y(n5417) );
  CLKMX2X2 U5302 ( .A(hd_a18[0]), .B(d18[0]), .S0(n8673), .Y(n5416) );
  CLKMX2X2 U5303 ( .A(hd_a19[35]), .B(d19[35]), .S0(n8673), .Y(n5415) );
  CLKMX2X2 U5304 ( .A(hd_a19[34]), .B(d19[34]), .S0(n8673), .Y(n5414) );
  CLKMX2X2 U5305 ( .A(hd_a19[33]), .B(d19[33]), .S0(n8672), .Y(n5413) );
  CLKMX2X2 U5306 ( .A(hd_a19[32]), .B(d19[32]), .S0(n8672), .Y(n5412) );
  CLKMX2X2 U5307 ( .A(hd_a19[31]), .B(d19[31]), .S0(n8672), .Y(n5411) );
  CLKMX2X2 U5308 ( .A(hd_a19[30]), .B(d19[30]), .S0(n8672), .Y(n5410) );
  CLKMX2X2 U5309 ( .A(hd_a19[29]), .B(d19[29]), .S0(n8672), .Y(n5409) );
  CLKMX2X2 U5310 ( .A(hd_a19[28]), .B(d19[28]), .S0(n8672), .Y(n5408) );
  CLKMX2X2 U5311 ( .A(hd_a19[27]), .B(d19[27]), .S0(n8672), .Y(n5407) );
  CLKMX2X2 U5312 ( .A(hd_a19[26]), .B(d19[26]), .S0(n8672), .Y(n5406) );
  CLKMX2X2 U5313 ( .A(hd_a19[25]), .B(d19[25]), .S0(n8672), .Y(n5405) );
  CLKMX2X2 U5314 ( .A(hd_a19[24]), .B(d19[24]), .S0(n8672), .Y(n5404) );
  CLKMX2X2 U5315 ( .A(hd_a19[23]), .B(d19[23]), .S0(n8672), .Y(n5403) );
  CLKMX2X2 U5316 ( .A(hd_a19[22]), .B(d19[22]), .S0(n8672), .Y(n5402) );
  CLKMX2X2 U5317 ( .A(hd_a19[21]), .B(d19[21]), .S0(n8672), .Y(n5401) );
  CLKMX2X2 U5318 ( .A(hd_a19[20]), .B(d19[20]), .S0(n8671), .Y(n5400) );
  CLKMX2X2 U5319 ( .A(hd_a19[19]), .B(d19[19]), .S0(n8671), .Y(n5399) );
  CLKMX2X2 U5320 ( .A(hd_a19[18]), .B(d19[18]), .S0(n8671), .Y(n5398) );
  CLKMX2X2 U5321 ( .A(hd_a19[17]), .B(d19[17]), .S0(n8671), .Y(n5397) );
  CLKMX2X2 U5322 ( .A(hd_a19[16]), .B(d19[16]), .S0(n8671), .Y(n5396) );
  CLKMX2X2 U5323 ( .A(hd_a19[15]), .B(d19[15]), .S0(n8671), .Y(n5395) );
  CLKMX2X2 U5324 ( .A(hd_a19[14]), .B(d19[14]), .S0(n8671), .Y(n5394) );
  CLKMX2X2 U5325 ( .A(hd_a19[13]), .B(d19[13]), .S0(n8671), .Y(n5393) );
  CLKMX2X2 U5326 ( .A(hd_a19[12]), .B(d19[12]), .S0(n8671), .Y(n5392) );
  CLKMX2X2 U5327 ( .A(hd_a19[11]), .B(d19[11]), .S0(n8671), .Y(n5391) );
  CLKMX2X2 U5328 ( .A(hd_a19[10]), .B(d19[10]), .S0(n8671), .Y(n5390) );
  CLKMX2X2 U5329 ( .A(hd_a19[9]), .B(d19[9]), .S0(n8671), .Y(n5389) );
  CLKMX2X2 U5330 ( .A(hd_a19[8]), .B(d19[8]), .S0(n8671), .Y(n5388) );
  CLKMX2X2 U5331 ( .A(hd_a19[7]), .B(d19[7]), .S0(n8670), .Y(n5387) );
  CLKMX2X2 U5332 ( .A(hd_a19[6]), .B(d19[6]), .S0(n8670), .Y(n5386) );
  CLKMX2X2 U5333 ( .A(hd_a19[5]), .B(d19[5]), .S0(n8670), .Y(n5385) );
  CLKMX2X2 U5334 ( .A(hd_a19[4]), .B(d19[4]), .S0(n8670), .Y(n5384) );
  CLKMX2X2 U5335 ( .A(hd_a19[3]), .B(d19[3]), .S0(n8670), .Y(n5383) );
  CLKMX2X2 U5336 ( .A(hd_a19[2]), .B(d19[2]), .S0(n8670), .Y(n5382) );
  CLKMX2X2 U5337 ( .A(hd_a19[1]), .B(d19[1]), .S0(n8670), .Y(n5381) );
  CLKMX2X2 U5338 ( .A(hd_a19[0]), .B(d19[0]), .S0(n8670), .Y(n5380) );
  CLKMX2X2 U5339 ( .A(hd_a20[35]), .B(d20[35]), .S0(n8670), .Y(n5379) );
  CLKMX2X2 U5340 ( .A(hd_a20[34]), .B(d20[34]), .S0(n8670), .Y(n5378) );
  CLKMX2X2 U5341 ( .A(hd_a20[33]), .B(d20[33]), .S0(n8670), .Y(n5377) );
  CLKMX2X2 U5342 ( .A(hd_a20[32]), .B(d20[32]), .S0(n8670), .Y(n5376) );
  CLKMX2X2 U5343 ( .A(hd_a20[31]), .B(d20[31]), .S0(n8670), .Y(n5375) );
  CLKMX2X2 U5344 ( .A(hd_a20[30]), .B(d20[30]), .S0(n8669), .Y(n5374) );
  CLKMX2X2 U5345 ( .A(hd_a20[29]), .B(d20[29]), .S0(n8669), .Y(n5373) );
  CLKMX2X2 U5346 ( .A(hd_a20[28]), .B(d20[28]), .S0(n8669), .Y(n5372) );
  CLKMX2X2 U5347 ( .A(hd_a20[27]), .B(d20[27]), .S0(n8669), .Y(n5371) );
  CLKMX2X2 U5348 ( .A(hd_a20[26]), .B(d20[26]), .S0(n8669), .Y(n5370) );
  CLKMX2X2 U5349 ( .A(hd_a20[25]), .B(d20[25]), .S0(n8669), .Y(n5369) );
  CLKMX2X2 U5350 ( .A(hd_a20[24]), .B(d20[24]), .S0(n8669), .Y(n5368) );
  CLKMX2X2 U5351 ( .A(hd_a20[23]), .B(d20[23]), .S0(n8669), .Y(n5367) );
  CLKMX2X2 U5352 ( .A(hd_a20[22]), .B(d20[22]), .S0(n8669), .Y(n5366) );
  CLKMX2X2 U5353 ( .A(hd_a20[21]), .B(d20[21]), .S0(n8669), .Y(n5365) );
  CLKMX2X2 U5354 ( .A(hd_a20[20]), .B(d20[20]), .S0(n8669), .Y(n5364) );
  CLKMX2X2 U5355 ( .A(hd_a20[19]), .B(d20[19]), .S0(n8669), .Y(n5363) );
  CLKMX2X2 U5356 ( .A(hd_a20[18]), .B(d20[18]), .S0(n8669), .Y(n5362) );
  CLKMX2X2 U5357 ( .A(hd_a20[17]), .B(d20[17]), .S0(n8668), .Y(n5361) );
  CLKMX2X2 U5358 ( .A(hd_a20[16]), .B(d20[16]), .S0(n8668), .Y(n5360) );
  CLKMX2X2 U5359 ( .A(hd_a20[15]), .B(d20[15]), .S0(n8668), .Y(n5359) );
  CLKMX2X2 U5360 ( .A(hd_a20[14]), .B(d20[14]), .S0(n8668), .Y(n5358) );
  CLKMX2X2 U5361 ( .A(hd_a20[13]), .B(d20[13]), .S0(n8668), .Y(n5357) );
  CLKMX2X2 U5362 ( .A(hd_a20[12]), .B(d20[12]), .S0(n8668), .Y(n5356) );
  CLKMX2X2 U5363 ( .A(hd_a20[11]), .B(d20[11]), .S0(n8668), .Y(n5355) );
  CLKMX2X2 U5364 ( .A(hd_a20[10]), .B(d20[10]), .S0(n8668), .Y(n5354) );
  CLKMX2X2 U5365 ( .A(hd_a20[9]), .B(d20[9]), .S0(n8668), .Y(n5353) );
  CLKMX2X2 U5366 ( .A(hd_a20[8]), .B(d20[8]), .S0(n8673), .Y(n5352) );
  CLKMX2X2 U5367 ( .A(hd_a20[7]), .B(d20[7]), .S0(n8689), .Y(n5351) );
  CLKMX2X2 U5368 ( .A(hd_a20[6]), .B(d20[6]), .S0(n8689), .Y(n5350) );
  CLKMX2X2 U5369 ( .A(hd_a20[5]), .B(d20[5]), .S0(n8689), .Y(n5349) );
  CLKMX2X2 U5370 ( .A(hd_a20[4]), .B(d20[4]), .S0(n8689), .Y(n5348) );
  CLKMX2X2 U5371 ( .A(hd_a20[3]), .B(d20[3]), .S0(n8689), .Y(n5347) );
  CLKMX2X2 U5372 ( .A(hd_a20[2]), .B(d20[2]), .S0(n8689), .Y(n5346) );
  CLKMX2X2 U5373 ( .A(hd_a20[1]), .B(d20[1]), .S0(n8689), .Y(n5345) );
  CLKMX2X2 U5374 ( .A(hd_a20[0]), .B(d20[0]), .S0(n8689), .Y(n5344) );
  CLKMX2X2 U5375 ( .A(hd_a21[35]), .B(d21[35]), .S0(n8689), .Y(n5343) );
  CLKMX2X2 U5376 ( .A(hd_a21[34]), .B(d21[34]), .S0(n8688), .Y(n5342) );
  CLKMX2X2 U5377 ( .A(hd_a21[33]), .B(d21[33]), .S0(n8688), .Y(n5341) );
  CLKMX2X2 U5378 ( .A(hd_a21[32]), .B(d21[32]), .S0(n8688), .Y(n5340) );
  CLKMX2X2 U5379 ( .A(hd_a21[31]), .B(d21[31]), .S0(n8688), .Y(n5339) );
  CLKMX2X2 U5380 ( .A(hd_a21[30]), .B(d21[30]), .S0(n8688), .Y(n5338) );
  CLKMX2X2 U5381 ( .A(hd_a21[29]), .B(d21[29]), .S0(n8688), .Y(n5337) );
  CLKMX2X2 U5382 ( .A(hd_a21[28]), .B(d21[28]), .S0(n8688), .Y(n5336) );
  CLKMX2X2 U5383 ( .A(hd_a21[27]), .B(d21[27]), .S0(n8688), .Y(n5335) );
  CLKMX2X2 U5384 ( .A(hd_a21[26]), .B(d21[26]), .S0(n8688), .Y(n5334) );
  CLKMX2X2 U5385 ( .A(hd_a21[25]), .B(d21[25]), .S0(n8688), .Y(n5333) );
  CLKMX2X2 U5386 ( .A(hd_a21[24]), .B(d21[24]), .S0(n8688), .Y(n5332) );
  CLKMX2X2 U5387 ( .A(hd_a21[23]), .B(d21[23]), .S0(n8688), .Y(n5331) );
  CLKMX2X2 U5388 ( .A(hd_a21[22]), .B(d21[22]), .S0(n8688), .Y(n5330) );
  CLKMX2X2 U5389 ( .A(hd_a21[21]), .B(d21[21]), .S0(n8687), .Y(n5329) );
  CLKMX2X2 U5390 ( .A(hd_a21[20]), .B(d21[20]), .S0(n8687), .Y(n5328) );
  CLKMX2X2 U5391 ( .A(hd_a21[19]), .B(d21[19]), .S0(n8687), .Y(n5327) );
  CLKMX2X2 U5392 ( .A(hd_a21[18]), .B(d21[18]), .S0(n8687), .Y(n5326) );
  CLKMX2X2 U5393 ( .A(hd_a21[17]), .B(d21[17]), .S0(n8687), .Y(n5325) );
  CLKMX2X2 U5394 ( .A(hd_a21[16]), .B(d21[16]), .S0(n8687), .Y(n5324) );
  CLKMX2X2 U5395 ( .A(hd_a21[15]), .B(d21[15]), .S0(n8687), .Y(n5323) );
  CLKMX2X2 U5396 ( .A(hd_a21[14]), .B(d21[14]), .S0(n8687), .Y(n5322) );
  CLKMX2X2 U5397 ( .A(hd_a21[13]), .B(d21[13]), .S0(n8687), .Y(n5321) );
  CLKMX2X2 U5398 ( .A(hd_a21[12]), .B(d21[12]), .S0(n8687), .Y(n5320) );
  CLKMX2X2 U5399 ( .A(hd_a21[11]), .B(d21[11]), .S0(n8687), .Y(n5319) );
  CLKMX2X2 U5400 ( .A(hd_a21[10]), .B(d21[10]), .S0(n8687), .Y(n5318) );
  CLKMX2X2 U5401 ( .A(hd_a21[9]), .B(d21[9]), .S0(n8687), .Y(n5317) );
  CLKMX2X2 U5402 ( .A(hd_a21[8]), .B(d21[8]), .S0(n8686), .Y(n5316) );
  CLKMX2X2 U5403 ( .A(hd_a21[7]), .B(d21[7]), .S0(n8686), .Y(n5315) );
  CLKMX2X2 U5404 ( .A(hd_a21[6]), .B(d21[6]), .S0(n8686), .Y(n5314) );
  CLKMX2X2 U5405 ( .A(hd_a21[5]), .B(d21[5]), .S0(n8686), .Y(n5313) );
  CLKMX2X2 U5406 ( .A(hd_a21[4]), .B(d21[4]), .S0(n8686), .Y(n5312) );
  CLKMX2X2 U5407 ( .A(hd_a21[3]), .B(d21[3]), .S0(n8686), .Y(n5311) );
  CLKMX2X2 U5408 ( .A(hd_a21[2]), .B(d21[2]), .S0(n8686), .Y(n5310) );
  CLKMX2X2 U5409 ( .A(hd_a21[1]), .B(d21[1]), .S0(n8686), .Y(n5309) );
  CLKMX2X2 U5410 ( .A(hd_a21[0]), .B(d21[0]), .S0(n8686), .Y(n5308) );
  CLKMX2X2 U5411 ( .A(hd_a22[35]), .B(d22[35]), .S0(n8686), .Y(n5307) );
  CLKMX2X2 U5412 ( .A(hd_a22[34]), .B(d22[34]), .S0(n8686), .Y(n5306) );
  CLKMX2X2 U5413 ( .A(hd_a22[33]), .B(d22[33]), .S0(n8686), .Y(n5305) );
  CLKMX2X2 U5414 ( .A(hd_a22[32]), .B(d22[32]), .S0(n8686), .Y(n5304) );
  CLKMX2X2 U5415 ( .A(hd_a22[31]), .B(d22[31]), .S0(n8685), .Y(n5303) );
  CLKMX2X2 U5416 ( .A(hd_a22[30]), .B(d22[30]), .S0(n8685), .Y(n5302) );
  CLKMX2X2 U5417 ( .A(hd_a22[29]), .B(d22[29]), .S0(n8685), .Y(n5301) );
  CLKMX2X2 U5418 ( .A(hd_a22[28]), .B(d22[28]), .S0(n8685), .Y(n5300) );
  CLKMX2X2 U5419 ( .A(hd_a22[27]), .B(d22[27]), .S0(n8685), .Y(n5299) );
  CLKMX2X2 U5420 ( .A(hd_a22[26]), .B(d22[26]), .S0(n8685), .Y(n5298) );
  CLKMX2X2 U5421 ( .A(hd_a22[25]), .B(d22[25]), .S0(n8685), .Y(n5297) );
  CLKMX2X2 U5422 ( .A(hd_a22[24]), .B(d22[24]), .S0(n8685), .Y(n5296) );
  CLKMX2X2 U5423 ( .A(hd_a22[23]), .B(d22[23]), .S0(n8685), .Y(n5295) );
  CLKMX2X2 U5424 ( .A(hd_a22[22]), .B(d22[22]), .S0(n8685), .Y(n5294) );
  CLKMX2X2 U5425 ( .A(hd_a22[21]), .B(d22[21]), .S0(n8685), .Y(n5293) );
  CLKMX2X2 U5426 ( .A(hd_a22[20]), .B(d22[20]), .S0(n8685), .Y(n5292) );
  CLKMX2X2 U5427 ( .A(hd_a22[19]), .B(d22[19]), .S0(n8685), .Y(n5291) );
  CLKMX2X2 U5428 ( .A(hd_a22[18]), .B(d22[18]), .S0(n8684), .Y(n5290) );
  CLKMX2X2 U5429 ( .A(hd_a22[17]), .B(d22[17]), .S0(n8684), .Y(n5289) );
  CLKMX2X2 U5430 ( .A(hd_a22[16]), .B(d22[16]), .S0(n8684), .Y(n5288) );
  CLKMX2X2 U5431 ( .A(hd_a22[15]), .B(d22[15]), .S0(n8684), .Y(n5287) );
  CLKMX2X2 U5432 ( .A(hd_a22[14]), .B(d22[14]), .S0(n8684), .Y(n5286) );
  CLKMX2X2 U5433 ( .A(hd_a22[13]), .B(d22[13]), .S0(n8684), .Y(n5285) );
  CLKMX2X2 U5434 ( .A(hd_a22[12]), .B(d22[12]), .S0(n8684), .Y(n5284) );
  CLKMX2X2 U5435 ( .A(hd_a22[11]), .B(d22[11]), .S0(n8684), .Y(n5283) );
  CLKMX2X2 U5436 ( .A(hd_a22[10]), .B(d22[10]), .S0(n8684), .Y(n5282) );
  CLKMX2X2 U5437 ( .A(hd_a22[9]), .B(d22[9]), .S0(n8684), .Y(n5281) );
  CLKMX2X2 U5438 ( .A(hd_a22[8]), .B(d22[8]), .S0(n8684), .Y(n5280) );
  CLKMX2X2 U5439 ( .A(hd_a22[7]), .B(d22[7]), .S0(n8684), .Y(n5279) );
  CLKMX2X2 U5440 ( .A(hd_a22[6]), .B(d22[6]), .S0(n8683), .Y(n5278) );
  CLKMX2X2 U5441 ( .A(hd_a22[5]), .B(d22[5]), .S0(n8683), .Y(n5277) );
  CLKMX2X2 U5442 ( .A(hd_a22[4]), .B(d22[4]), .S0(n8683), .Y(n5276) );
  CLKMX2X2 U5443 ( .A(hd_a22[3]), .B(d22[3]), .S0(n8683), .Y(n5275) );
  CLKMX2X2 U5444 ( .A(hd_a22[2]), .B(d22[2]), .S0(n8683), .Y(n5274) );
  CLKMX2X2 U5445 ( .A(hd_a22[1]), .B(d22[1]), .S0(n8683), .Y(n5273) );
  CLKMX2X2 U5446 ( .A(hd_a22[0]), .B(d22[0]), .S0(n8683), .Y(n5272) );
  CLKMX2X2 U5447 ( .A(hd_a23[35]), .B(d23[35]), .S0(n8683), .Y(n5271) );
  CLKMX2X2 U5448 ( .A(hd_a23[34]), .B(d23[34]), .S0(n8683), .Y(n5270) );
  CLKMX2X2 U5449 ( .A(hd_a23[33]), .B(d23[33]), .S0(n8683), .Y(n5269) );
  CLKMX2X2 U5450 ( .A(hd_a23[32]), .B(d23[32]), .S0(n8683), .Y(n5268) );
  CLKMX2X2 U5451 ( .A(hd_a23[31]), .B(d23[31]), .S0(n8683), .Y(n5267) );
  CLKMX2X2 U5452 ( .A(hd_a23[30]), .B(d23[30]), .S0(n8683), .Y(n5266) );
  CLKMX2X2 U5453 ( .A(hd_a23[29]), .B(d23[29]), .S0(n8682), .Y(n5265) );
  CLKMX2X2 U5454 ( .A(hd_a23[28]), .B(d23[28]), .S0(n8682), .Y(n5264) );
  CLKMX2X2 U5455 ( .A(hd_a23[27]), .B(d23[27]), .S0(n8682), .Y(n5263) );
  CLKMX2X2 U5456 ( .A(hd_a23[26]), .B(d23[26]), .S0(n8682), .Y(n5262) );
  CLKMX2X2 U5457 ( .A(hd_a23[25]), .B(d23[25]), .S0(n8682), .Y(n5261) );
  CLKMX2X2 U5458 ( .A(hd_a23[24]), .B(d23[24]), .S0(n8682), .Y(n5260) );
  CLKMX2X2 U5459 ( .A(hd_a23[23]), .B(d23[23]), .S0(n8682), .Y(n5259) );
  CLKMX2X2 U5460 ( .A(hd_a23[22]), .B(d23[22]), .S0(n8682), .Y(n5258) );
  CLKMX2X2 U5461 ( .A(hd_a23[21]), .B(d23[21]), .S0(n8682), .Y(n5257) );
  CLKMX2X2 U5462 ( .A(hd_a23[20]), .B(d23[20]), .S0(n8682), .Y(n5256) );
  CLKMX2X2 U5463 ( .A(hd_a23[19]), .B(d23[19]), .S0(n8682), .Y(n5255) );
  CLKMX2X2 U5464 ( .A(hd_a23[18]), .B(d23[18]), .S0(n8682), .Y(n5254) );
  CLKMX2X2 U5465 ( .A(hd_a23[17]), .B(d23[17]), .S0(n8682), .Y(n5253) );
  CLKMX2X2 U5466 ( .A(hd_a23[16]), .B(d23[16]), .S0(n8681), .Y(n5252) );
  CLKMX2X2 U5467 ( .A(hd_a23[15]), .B(d23[15]), .S0(n8681), .Y(n5251) );
  CLKMX2X2 U5468 ( .A(hd_a23[14]), .B(d23[14]), .S0(n8681), .Y(n5250) );
  CLKMX2X2 U5469 ( .A(hd_a23[13]), .B(d23[13]), .S0(n8681), .Y(n5249) );
  CLKMX2X2 U5470 ( .A(hd_a23[12]), .B(d23[12]), .S0(n8681), .Y(n5248) );
  CLKMX2X2 U5471 ( .A(hd_a23[11]), .B(d23[11]), .S0(n8681), .Y(n5247) );
  CLKMX2X2 U5472 ( .A(hd_a23[10]), .B(d23[10]), .S0(n8681), .Y(n5246) );
  CLKMX2X2 U5473 ( .A(hd_a23[9]), .B(d23[9]), .S0(n8681), .Y(n5245) );
  CLKMX2X2 U5474 ( .A(hd_a23[8]), .B(d23[8]), .S0(n8681), .Y(n5244) );
  CLKMX2X2 U5475 ( .A(hd_a23[7]), .B(d23[7]), .S0(n8681), .Y(n5243) );
  CLKMX2X2 U5476 ( .A(hd_a23[6]), .B(d23[6]), .S0(n8681), .Y(n5242) );
  CLKMX2X2 U5477 ( .A(hd_a23[5]), .B(d23[5]), .S0(n8681), .Y(n5241) );
  CLKMX2X2 U5478 ( .A(hd_a23[4]), .B(d23[4]), .S0(n8681), .Y(n5240) );
  CLKMX2X2 U5479 ( .A(hd_a23[3]), .B(d23[3]), .S0(n8680), .Y(n5239) );
  CLKMX2X2 U5480 ( .A(hd_a23[2]), .B(d23[2]), .S0(n8680), .Y(n5238) );
  CLKMX2X2 U5481 ( .A(hd_a23[1]), .B(d23[1]), .S0(n8680), .Y(n5237) );
  CLKMX2X2 U5482 ( .A(hd_a23[0]), .B(d23[0]), .S0(n8680), .Y(n5236) );
  CLKMX2X2 U5483 ( .A(hd_a24[35]), .B(d24[35]), .S0(n8680), .Y(n5235) );
  CLKMX2X2 U5484 ( .A(hd_a24[34]), .B(d24[34]), .S0(n8680), .Y(n5234) );
  CLKMX2X2 U5485 ( .A(hd_a24[33]), .B(d24[33]), .S0(n8680), .Y(n5233) );
  CLKMX2X2 U5486 ( .A(hd_a24[32]), .B(d24[32]), .S0(n8680), .Y(n5232) );
  CLKMX2X2 U5487 ( .A(hd_a24[31]), .B(d24[31]), .S0(n8680), .Y(n5231) );
  CLKMX2X2 U5488 ( .A(hd_a24[30]), .B(d24[30]), .S0(n8680), .Y(n5230) );
  CLKMX2X2 U5489 ( .A(hd_a24[29]), .B(d24[29]), .S0(n8680), .Y(n5229) );
  CLKMX2X2 U5490 ( .A(hd_a24[28]), .B(d24[28]), .S0(n8680), .Y(n5228) );
  CLKMX2X2 U5491 ( .A(hd_a24[27]), .B(d24[27]), .S0(n8680), .Y(n5227) );
  CLKMX2X2 U5492 ( .A(hd_a24[26]), .B(d24[26]), .S0(n8679), .Y(n5226) );
  CLKMX2X2 U5493 ( .A(hd_a24[25]), .B(d24[25]), .S0(n8679), .Y(n5225) );
  CLKMX2X2 U5494 ( .A(hd_a24[24]), .B(d24[24]), .S0(n8679), .Y(n5224) );
  CLKMX2X2 U5495 ( .A(hd_a24[23]), .B(d24[23]), .S0(n8679), .Y(n5223) );
  CLKMX2X2 U5496 ( .A(hd_a24[22]), .B(d24[22]), .S0(n8679), .Y(n5222) );
  CLKMX2X2 U5497 ( .A(hd_a24[21]), .B(d24[21]), .S0(n8679), .Y(n5221) );
  CLKMX2X2 U5498 ( .A(hd_a24[20]), .B(d24[20]), .S0(n8679), .Y(n5220) );
  CLKMX2X2 U5499 ( .A(hd_a24[19]), .B(d24[19]), .S0(n8679), .Y(n5219) );
  CLKMX2X2 U5500 ( .A(hd_a24[18]), .B(d24[18]), .S0(n8679), .Y(n5218) );
  CLKMX2X2 U5501 ( .A(hd_a24[17]), .B(d24[17]), .S0(n8679), .Y(n5217) );
  CLKMX2X2 U5502 ( .A(hd_a24[16]), .B(d24[16]), .S0(n8679), .Y(n5216) );
  CLKMX2X2 U5503 ( .A(hd_a24[15]), .B(d24[15]), .S0(n8679), .Y(n5215) );
  CLKMX2X2 U5504 ( .A(hd_a24[14]), .B(d24[14]), .S0(n8684), .Y(n5214) );
  CLKMX2X2 U5505 ( .A(hd_a24[13]), .B(d24[13]), .S0(n8657), .Y(n5213) );
  CLKMX2X2 U5506 ( .A(hd_a24[12]), .B(d24[12]), .S0(n8657), .Y(n5212) );
  CLKMX2X2 U5507 ( .A(hd_a24[11]), .B(d24[11]), .S0(n8657), .Y(n5211) );
  CLKMX2X2 U5508 ( .A(hd_a24[10]), .B(d24[10]), .S0(n8657), .Y(n5210) );
  CLKMX2X2 U5509 ( .A(hd_a24[9]), .B(d24[9]), .S0(n8657), .Y(n5209) );
  CLKMX2X2 U5510 ( .A(hd_a24[8]), .B(d24[8]), .S0(n8657), .Y(n5208) );
  CLKMX2X2 U5511 ( .A(hd_a24[7]), .B(d24[7]), .S0(n8657), .Y(n5207) );
  CLKMX2X2 U5512 ( .A(hd_a24[6]), .B(d24[6]), .S0(n8657), .Y(n5206) );
  CLKMX2X2 U5513 ( .A(hd_a24[5]), .B(d24[5]), .S0(n8656), .Y(n5205) );
  CLKMX2X2 U5514 ( .A(hd_a24[4]), .B(d24[4]), .S0(n8656), .Y(n5204) );
  CLKMX2X2 U5515 ( .A(hd_a24[3]), .B(d24[3]), .S0(n8656), .Y(n5203) );
  CLKMX2X2 U5516 ( .A(hd_a24[2]), .B(d24[2]), .S0(n8656), .Y(n5202) );
  CLKMX2X2 U5517 ( .A(hd_a24[1]), .B(d24[1]), .S0(n8656), .Y(n5201) );
  CLKMX2X2 U5518 ( .A(hd_a24[0]), .B(d24[0]), .S0(n8656), .Y(n5200) );
  CLKMX2X2 U5519 ( .A(hd_a25[35]), .B(d25[35]), .S0(n8656), .Y(n5199) );
  CLKMX2X2 U5520 ( .A(hd_a25[34]), .B(d25[34]), .S0(n8656), .Y(n5198) );
  CLKMX2X2 U5521 ( .A(hd_a25[33]), .B(d25[33]), .S0(n8656), .Y(n5197) );
  CLKMX2X2 U5522 ( .A(hd_a25[32]), .B(d25[32]), .S0(n8656), .Y(n5196) );
  CLKMX2X2 U5523 ( .A(hd_a25[31]), .B(d25[31]), .S0(n8656), .Y(n5195) );
  CLKMX2X2 U5524 ( .A(hd_a25[30]), .B(d25[30]), .S0(n8656), .Y(n5194) );
  CLKMX2X2 U5525 ( .A(hd_a25[29]), .B(d25[29]), .S0(n8656), .Y(n5193) );
  CLKMX2X2 U5526 ( .A(hd_a25[28]), .B(d25[28]), .S0(n8655), .Y(n5192) );
  CLKMX2X2 U5527 ( .A(hd_a25[27]), .B(d25[27]), .S0(n8655), .Y(n5191) );
  CLKMX2X2 U5528 ( .A(hd_a25[26]), .B(d25[26]), .S0(n8655), .Y(n5190) );
  CLKMX2X2 U5529 ( .A(hd_a25[25]), .B(d25[25]), .S0(n8655), .Y(n5189) );
  CLKMX2X2 U5530 ( .A(hd_a25[24]), .B(d25[24]), .S0(n8655), .Y(n5188) );
  CLKMX2X2 U5531 ( .A(hd_a25[23]), .B(d25[23]), .S0(n8655), .Y(n5187) );
  CLKMX2X2 U5532 ( .A(hd_a25[22]), .B(d25[22]), .S0(n8655), .Y(n5186) );
  CLKMX2X2 U5533 ( .A(hd_a25[21]), .B(d25[21]), .S0(n8655), .Y(n5185) );
  CLKMX2X2 U5534 ( .A(hd_a25[20]), .B(d25[20]), .S0(n8655), .Y(n5184) );
  CLKMX2X2 U5535 ( .A(hd_a25[19]), .B(d25[19]), .S0(n8655), .Y(n5183) );
  CLKMX2X2 U5536 ( .A(hd_a25[18]), .B(d25[18]), .S0(n8655), .Y(n5182) );
  CLKMX2X2 U5537 ( .A(hd_a25[17]), .B(d25[17]), .S0(n8655), .Y(n5181) );
  CLKMX2X2 U5538 ( .A(hd_a25[16]), .B(d25[16]), .S0(n8655), .Y(n5180) );
  CLKMX2X2 U5539 ( .A(hd_a25[15]), .B(d25[15]), .S0(n8654), .Y(n5179) );
  CLKMX2X2 U5540 ( .A(hd_a25[14]), .B(d25[14]), .S0(n8654), .Y(n5178) );
  CLKMX2X2 U5541 ( .A(hd_a25[13]), .B(d25[13]), .S0(n8654), .Y(n5177) );
  CLKMX2X2 U5542 ( .A(hd_a25[12]), .B(d25[12]), .S0(n8654), .Y(n5176) );
  CLKMX2X2 U5543 ( .A(hd_a25[11]), .B(d25[11]), .S0(n8654), .Y(n5175) );
  CLKMX2X2 U5544 ( .A(hd_a25[10]), .B(d25[10]), .S0(n8654), .Y(n5174) );
  CLKMX2X2 U5545 ( .A(hd_a25[9]), .B(d25[9]), .S0(n8654), .Y(n5173) );
  CLKMX2X2 U5546 ( .A(hd_a25[8]), .B(d25[8]), .S0(n8654), .Y(n5172) );
  CLKMX2X2 U5547 ( .A(hd_a25[7]), .B(d25[7]), .S0(n8654), .Y(n5171) );
  CLKMX2X2 U5548 ( .A(hd_a25[6]), .B(d25[6]), .S0(n8654), .Y(n5170) );
  CLKMX2X2 U5549 ( .A(hd_a25[5]), .B(d25[5]), .S0(n8654), .Y(n5169) );
  CLKMX2X2 U5550 ( .A(hd_a25[4]), .B(d25[4]), .S0(n8654), .Y(n5168) );
  CLKMX2X2 U5551 ( .A(hd_a25[3]), .B(d25[3]), .S0(n8654), .Y(n5167) );
  CLKMX2X2 U5552 ( .A(hd_a25[2]), .B(d25[2]), .S0(n8653), .Y(n5166) );
  CLKMX2X2 U5553 ( .A(hd_a25[1]), .B(d25[1]), .S0(n8653), .Y(n5165) );
  CLKMX2X2 U5554 ( .A(hd_a25[0]), .B(d25[0]), .S0(n8653), .Y(n5164) );
  CLKMX2X2 U5555 ( .A(hd_a26[35]), .B(d26[35]), .S0(n8653), .Y(n5163) );
  CLKMX2X2 U5556 ( .A(hd_a26[34]), .B(d26[34]), .S0(n8653), .Y(n5162) );
  CLKMX2X2 U5557 ( .A(hd_a26[33]), .B(d26[33]), .S0(n8653), .Y(n5161) );
  CLKMX2X2 U5558 ( .A(hd_a26[32]), .B(d26[32]), .S0(n8653), .Y(n5160) );
  CLKMX2X2 U5559 ( .A(hd_a26[31]), .B(d26[31]), .S0(n8653), .Y(n5159) );
  CLKMX2X2 U5560 ( .A(hd_a26[30]), .B(d26[30]), .S0(n8653), .Y(n5158) );
  CLKMX2X2 U5561 ( .A(hd_a26[29]), .B(d26[29]), .S0(n8653), .Y(n5157) );
  CLKMX2X2 U5562 ( .A(hd_a26[28]), .B(d26[28]), .S0(n8653), .Y(n5156) );
  CLKMX2X2 U5563 ( .A(hd_a26[27]), .B(d26[27]), .S0(n8653), .Y(n5155) );
  CLKMX2X2 U5564 ( .A(hd_a26[26]), .B(d26[26]), .S0(n8653), .Y(n5154) );
  CLKMX2X2 U5565 ( .A(hd_a26[25]), .B(d26[25]), .S0(n8652), .Y(n5153) );
  CLKMX2X2 U5566 ( .A(hd_a26[24]), .B(d26[24]), .S0(n8652), .Y(n5152) );
  CLKMX2X2 U5567 ( .A(hd_a26[23]), .B(d26[23]), .S0(n8652), .Y(n5151) );
  CLKMX2X2 U5568 ( .A(hd_a26[22]), .B(d26[22]), .S0(n8652), .Y(n5150) );
  CLKMX2X2 U5569 ( .A(hd_a26[21]), .B(d26[21]), .S0(n8652), .Y(n5149) );
  CLKMX2X2 U5570 ( .A(hd_a26[20]), .B(d26[20]), .S0(n8652), .Y(n5148) );
  CLKMX2X2 U5571 ( .A(hd_a26[19]), .B(d26[19]), .S0(n8652), .Y(n5147) );
  CLKMX2X2 U5572 ( .A(hd_a26[18]), .B(d26[18]), .S0(n8652), .Y(n5146) );
  CLKMX2X2 U5573 ( .A(hd_a26[17]), .B(d26[17]), .S0(n8652), .Y(n5145) );
  CLKMX2X2 U5574 ( .A(hd_a26[16]), .B(d26[16]), .S0(n8652), .Y(n5144) );
  CLKMX2X2 U5575 ( .A(hd_a26[15]), .B(d26[15]), .S0(n8652), .Y(n5143) );
  CLKMX2X2 U5576 ( .A(hd_a26[14]), .B(d26[14]), .S0(n8652), .Y(n5142) );
  CLKMX2X2 U5577 ( .A(hd_a26[13]), .B(d26[13]), .S0(n8651), .Y(n5141) );
  CLKMX2X2 U5578 ( .A(hd_a26[12]), .B(d26[12]), .S0(n8651), .Y(n5140) );
  CLKMX2X2 U5579 ( .A(hd_a26[11]), .B(d26[11]), .S0(n8651), .Y(n5139) );
  CLKMX2X2 U5580 ( .A(hd_a26[10]), .B(d26[10]), .S0(n8651), .Y(n5138) );
  CLKMX2X2 U5581 ( .A(hd_a26[9]), .B(d26[9]), .S0(n8651), .Y(n5137) );
  CLKMX2X2 U5582 ( .A(hd_a26[8]), .B(d26[8]), .S0(n8651), .Y(n5136) );
  CLKMX2X2 U5583 ( .A(hd_a26[7]), .B(d26[7]), .S0(n8651), .Y(n5135) );
  CLKMX2X2 U5584 ( .A(hd_a26[6]), .B(d26[6]), .S0(n8651), .Y(n5134) );
  CLKMX2X2 U5585 ( .A(hd_a26[5]), .B(d26[5]), .S0(n8651), .Y(n5133) );
  CLKMX2X2 U5586 ( .A(hd_a26[4]), .B(d26[4]), .S0(n8651), .Y(n5132) );
  CLKMX2X2 U5587 ( .A(hd_a26[3]), .B(d26[3]), .S0(n8651), .Y(n5131) );
  CLKMX2X2 U5588 ( .A(hd_a26[2]), .B(d26[2]), .S0(n8651), .Y(n5130) );
  CLKMX2X2 U5589 ( .A(hd_a26[1]), .B(d26[1]), .S0(n8651), .Y(n5129) );
  CLKMX2X2 U5590 ( .A(hd_a26[0]), .B(d26[0]), .S0(n8650), .Y(n5128) );
  CLKMX2X2 U5591 ( .A(hd_a27[35]), .B(d27[35]), .S0(n8650), .Y(n5127) );
  CLKMX2X2 U5592 ( .A(hd_a27[34]), .B(d27[34]), .S0(n8650), .Y(n5126) );
  CLKMX2X2 U5593 ( .A(hd_a27[33]), .B(d27[33]), .S0(n8650), .Y(n5125) );
  CLKMX2X2 U5594 ( .A(hd_a27[32]), .B(d27[32]), .S0(n8650), .Y(n5124) );
  CLKMX2X2 U5595 ( .A(hd_a27[31]), .B(d27[31]), .S0(n8650), .Y(n5123) );
  CLKMX2X2 U5596 ( .A(hd_a27[30]), .B(d27[30]), .S0(n8650), .Y(n5122) );
  CLKMX2X2 U5597 ( .A(hd_a27[29]), .B(d27[29]), .S0(n8650), .Y(n5121) );
  CLKMX2X2 U5598 ( .A(hd_a27[28]), .B(d27[28]), .S0(n8650), .Y(n5120) );
  CLKMX2X2 U5599 ( .A(hd_a27[27]), .B(d27[27]), .S0(n8650), .Y(n5119) );
  CLKMX2X2 U5600 ( .A(hd_a27[26]), .B(d27[26]), .S0(n8650), .Y(n5118) );
  CLKMX2X2 U5601 ( .A(hd_a27[25]), .B(d27[25]), .S0(n8650), .Y(n5117) );
  CLKMX2X2 U5602 ( .A(hd_a27[24]), .B(d27[24]), .S0(n8650), .Y(n5116) );
  CLKMX2X2 U5603 ( .A(hd_a27[23]), .B(d27[23]), .S0(n8649), .Y(n5115) );
  CLKMX2X2 U5604 ( .A(hd_a27[22]), .B(d27[22]), .S0(n8649), .Y(n5114) );
  CLKMX2X2 U5605 ( .A(hd_a27[21]), .B(d27[21]), .S0(n8649), .Y(n5113) );
  CLKMX2X2 U5606 ( .A(hd_a27[20]), .B(d27[20]), .S0(n8649), .Y(n5112) );
  CLKMX2X2 U5607 ( .A(hd_a27[19]), .B(d27[19]), .S0(n8649), .Y(n5111) );
  CLKMX2X2 U5608 ( .A(hd_a27[18]), .B(d27[18]), .S0(n8649), .Y(n5110) );
  CLKMX2X2 U5609 ( .A(hd_a27[17]), .B(d27[17]), .S0(n8649), .Y(n5109) );
  CLKMX2X2 U5610 ( .A(hd_a27[16]), .B(d27[16]), .S0(n8649), .Y(n5108) );
  CLKMX2X2 U5611 ( .A(hd_a27[15]), .B(d27[15]), .S0(n8649), .Y(n5107) );
  CLKMX2X2 U5612 ( .A(hd_a27[14]), .B(d27[14]), .S0(n8649), .Y(n5106) );
  CLKMX2X2 U5613 ( .A(hd_a27[13]), .B(d27[13]), .S0(n8649), .Y(n5105) );
  CLKMX2X2 U5614 ( .A(hd_a27[12]), .B(d27[12]), .S0(n8649), .Y(n5104) );
  CLKMX2X2 U5615 ( .A(hd_a27[11]), .B(d27[11]), .S0(n8649), .Y(n5103) );
  CLKMX2X2 U5616 ( .A(hd_a27[10]), .B(d27[10]), .S0(n8648), .Y(n5102) );
  CLKMX2X2 U5617 ( .A(hd_a27[9]), .B(d27[9]), .S0(n8648), .Y(n5101) );
  CLKMX2X2 U5618 ( .A(hd_a27[8]), .B(d27[8]), .S0(n8648), .Y(n5100) );
  CLKMX2X2 U5619 ( .A(hd_a27[7]), .B(d27[7]), .S0(n8648), .Y(n5099) );
  CLKMX2X2 U5620 ( .A(hd_a27[6]), .B(d27[6]), .S0(n8648), .Y(n5098) );
  CLKMX2X2 U5621 ( .A(hd_a27[5]), .B(d27[5]), .S0(n8648), .Y(n5097) );
  CLKMX2X2 U5622 ( .A(hd_a27[4]), .B(d27[4]), .S0(n8648), .Y(n5096) );
  CLKMX2X2 U5623 ( .A(hd_a27[3]), .B(d27[3]), .S0(n8648), .Y(n5095) );
  CLKMX2X2 U5624 ( .A(hd_a27[2]), .B(d27[2]), .S0(n8648), .Y(n5094) );
  CLKMX2X2 U5625 ( .A(hd_a27[1]), .B(d27[1]), .S0(n8648), .Y(n5093) );
  CLKMX2X2 U5626 ( .A(hd_a27[0]), .B(d27[0]), .S0(n8648), .Y(n5092) );
  CLKMX2X2 U5627 ( .A(hd_a28[35]), .B(d28[35]), .S0(n8648), .Y(n5091) );
  CLKMX2X2 U5628 ( .A(hd_a28[34]), .B(d28[34]), .S0(n8648), .Y(n5090) );
  CLKMX2X2 U5629 ( .A(hd_a28[33]), .B(d28[33]), .S0(n8647), .Y(n5089) );
  CLKMX2X2 U5630 ( .A(hd_a28[32]), .B(d28[32]), .S0(n8647), .Y(n5088) );
  CLKMX2X2 U5631 ( .A(hd_a28[31]), .B(d28[31]), .S0(n8647), .Y(n5087) );
  CLKMX2X2 U5632 ( .A(hd_a28[30]), .B(d28[30]), .S0(n8647), .Y(n5086) );
  CLKMX2X2 U5633 ( .A(hd_a28[29]), .B(d28[29]), .S0(n8647), .Y(n5085) );
  CLKMX2X2 U5634 ( .A(hd_a28[28]), .B(d28[28]), .S0(n8647), .Y(n5084) );
  CLKMX2X2 U5635 ( .A(hd_a28[27]), .B(d28[27]), .S0(n8647), .Y(n5083) );
  CLKMX2X2 U5636 ( .A(hd_a28[26]), .B(d28[26]), .S0(n8647), .Y(n5082) );
  CLKMX2X2 U5637 ( .A(hd_a28[25]), .B(d28[25]), .S0(n8647), .Y(n5081) );
  CLKMX2X2 U5638 ( .A(hd_a28[24]), .B(d28[24]), .S0(n8647), .Y(n5080) );
  CLKMX2X2 U5639 ( .A(hd_a28[23]), .B(d28[23]), .S0(n8647), .Y(n5079) );
  CLKMX2X2 U5640 ( .A(hd_a28[22]), .B(d28[22]), .S0(n8647), .Y(n5078) );
  CLKMX2X2 U5641 ( .A(hd_a28[21]), .B(d28[21]), .S0(n8647), .Y(n5077) );
  CLKMX2X2 U5642 ( .A(hd_a28[20]), .B(d28[20]), .S0(n8646), .Y(n5076) );
  CLKMX2X2 U5643 ( .A(hd_a28[19]), .B(d28[19]), .S0(n8652), .Y(n5075) );
  CLKMX2X2 U5644 ( .A(hd_a28[18]), .B(d28[18]), .S0(n8668), .Y(n5074) );
  CLKMX2X2 U5645 ( .A(hd_a28[17]), .B(d28[17]), .S0(n8668), .Y(n5073) );
  CLKMX2X2 U5646 ( .A(hd_a28[16]), .B(d28[16]), .S0(n8668), .Y(n5072) );
  CLKMX2X2 U5647 ( .A(hd_a28[15]), .B(d28[15]), .S0(n8667), .Y(n5071) );
  CLKMX2X2 U5648 ( .A(hd_a28[14]), .B(d28[14]), .S0(n8667), .Y(n5070) );
  CLKMX2X2 U5649 ( .A(hd_a28[13]), .B(d28[13]), .S0(n8667), .Y(n5069) );
  CLKMX2X2 U5650 ( .A(hd_a28[12]), .B(d28[12]), .S0(n8667), .Y(n5068) );
  CLKMX2X2 U5651 ( .A(hd_a28[11]), .B(d28[11]), .S0(n8668), .Y(n5067) );
  CLKMX2X2 U5652 ( .A(hd_a28[10]), .B(d28[10]), .S0(n8667), .Y(n5066) );
  CLKMX2X2 U5653 ( .A(hd_a28[9]), .B(d28[9]), .S0(n8667), .Y(n5065) );
  CLKMX2X2 U5654 ( .A(hd_a28[8]), .B(d28[8]), .S0(n8667), .Y(n5064) );
  CLKMX2X2 U5655 ( .A(hd_a28[7]), .B(d28[7]), .S0(n8667), .Y(n5063) );
  CLKMX2X2 U5656 ( .A(hd_a28[6]), .B(d28[6]), .S0(n8667), .Y(n5062) );
  CLKMX2X2 U5657 ( .A(hd_a28[5]), .B(d28[5]), .S0(n8667), .Y(n5061) );
  CLKMX2X2 U5658 ( .A(hd_a28[4]), .B(d28[4]), .S0(n8667), .Y(n5060) );
  CLKMX2X2 U5659 ( .A(hd_a28[3]), .B(d28[3]), .S0(n8667), .Y(n5059) );
  CLKMX2X2 U5660 ( .A(hd_a28[2]), .B(d28[2]), .S0(n8667), .Y(n5058) );
  CLKMX2X2 U5661 ( .A(hd_a28[1]), .B(d28[1]), .S0(n8666), .Y(n5057) );
  CLKMX2X2 U5662 ( .A(hd_a28[0]), .B(d28[0]), .S0(n8666), .Y(n5056) );
  CLKMX2X2 U5663 ( .A(hd_a29[35]), .B(d29[35]), .S0(n8666), .Y(n5055) );
  CLKMX2X2 U5664 ( .A(hd_a29[34]), .B(d29[34]), .S0(n8666), .Y(n5054) );
  CLKMX2X2 U5665 ( .A(hd_a29[33]), .B(d29[33]), .S0(n8666), .Y(n5053) );
  CLKMX2X2 U5666 ( .A(hd_a29[32]), .B(d29[32]), .S0(n8666), .Y(n5052) );
  CLKMX2X2 U5667 ( .A(hd_a29[31]), .B(d29[31]), .S0(n8666), .Y(n5051) );
  CLKMX2X2 U5668 ( .A(hd_a29[30]), .B(d29[30]), .S0(n8666), .Y(n5050) );
  CLKMX2X2 U5669 ( .A(hd_a29[29]), .B(d29[29]), .S0(n8666), .Y(n5049) );
  CLKMX2X2 U5670 ( .A(hd_a29[28]), .B(d29[28]), .S0(n8666), .Y(n5048) );
  CLKMX2X2 U5671 ( .A(hd_a29[27]), .B(d29[27]), .S0(n8666), .Y(n5047) );
  CLKMX2X2 U5672 ( .A(hd_a29[26]), .B(d29[26]), .S0(n8666), .Y(n5046) );
  CLKMX2X2 U5673 ( .A(hd_a29[25]), .B(d29[25]), .S0(n8666), .Y(n5045) );
  CLKMX2X2 U5674 ( .A(hd_a29[24]), .B(d29[24]), .S0(n8665), .Y(n5044) );
  CLKMX2X2 U5675 ( .A(hd_a29[23]), .B(d29[23]), .S0(n8665), .Y(n5043) );
  CLKMX2X2 U5676 ( .A(hd_a29[22]), .B(d29[22]), .S0(n8665), .Y(n5042) );
  CLKMX2X2 U5677 ( .A(hd_a29[21]), .B(d29[21]), .S0(n8665), .Y(n5041) );
  CLKMX2X2 U5678 ( .A(hd_a29[20]), .B(d29[20]), .S0(n8665), .Y(n5040) );
  CLKMX2X2 U5679 ( .A(hd_a29[19]), .B(d29[19]), .S0(n8665), .Y(n5039) );
  CLKMX2X2 U5680 ( .A(hd_a29[18]), .B(d29[18]), .S0(n8665), .Y(n5038) );
  CLKMX2X2 U5681 ( .A(hd_a29[17]), .B(d29[17]), .S0(n8665), .Y(n5037) );
  CLKMX2X2 U5682 ( .A(hd_a29[16]), .B(d29[16]), .S0(n8665), .Y(n5036) );
  CLKMX2X2 U5683 ( .A(hd_a29[15]), .B(d29[15]), .S0(n8665), .Y(n5035) );
  CLKMX2X2 U5684 ( .A(hd_a29[14]), .B(d29[14]), .S0(n8665), .Y(n5034) );
  CLKMX2X2 U5685 ( .A(hd_a29[13]), .B(d29[13]), .S0(n8665), .Y(n5033) );
  CLKMX2X2 U5686 ( .A(hd_a29[12]), .B(d29[12]), .S0(n8665), .Y(n5032) );
  CLKMX2X2 U5687 ( .A(hd_a29[11]), .B(d29[11]), .S0(n8664), .Y(n5031) );
  CLKMX2X2 U5688 ( .A(hd_a29[10]), .B(d29[10]), .S0(n8664), .Y(n5030) );
  CLKMX2X2 U5689 ( .A(hd_a29[9]), .B(d29[9]), .S0(n8664), .Y(n5029) );
  CLKMX2X2 U5690 ( .A(hd_a29[8]), .B(d29[8]), .S0(n8664), .Y(n5028) );
  CLKMX2X2 U5691 ( .A(hd_a29[7]), .B(d29[7]), .S0(n8664), .Y(n5027) );
  CLKMX2X2 U5692 ( .A(hd_a29[6]), .B(d29[6]), .S0(n8664), .Y(n5026) );
  CLKMX2X2 U5693 ( .A(hd_a29[5]), .B(d29[5]), .S0(n8664), .Y(n5025) );
  CLKMX2X2 U5694 ( .A(hd_a29[4]), .B(d29[4]), .S0(n8664), .Y(n5024) );
  CLKMX2X2 U5695 ( .A(hd_a29[3]), .B(d29[3]), .S0(n8664), .Y(n5023) );
  CLKMX2X2 U5696 ( .A(hd_a29[2]), .B(d29[2]), .S0(n8664), .Y(n5022) );
  CLKMX2X2 U5697 ( .A(hd_a29[1]), .B(d29[1]), .S0(n8664), .Y(n5021) );
  CLKMX2X2 U5698 ( .A(hd_a29[0]), .B(d29[0]), .S0(n8664), .Y(n5020) );
  CLKMX2X2 U5699 ( .A(hd_a30[0]), .B(d30[0]), .S0(n8664), .Y(n5019) );
  CLKMX2X2 U5700 ( .A(hd_a30[1]), .B(d30[1]), .S0(n8663), .Y(n5018) );
  CLKMX2X2 U5701 ( .A(hd_a30[2]), .B(d30[2]), .S0(n8663), .Y(n5017) );
  CLKMX2X2 U5702 ( .A(hd_a30[3]), .B(d30[3]), .S0(n8663), .Y(n5016) );
  CLKMX2X2 U5703 ( .A(hd_a30[4]), .B(d30[4]), .S0(n8663), .Y(n5015) );
  CLKMX2X2 U5704 ( .A(hd_a30[5]), .B(d30[5]), .S0(n8663), .Y(n5014) );
  CLKMX2X2 U5705 ( .A(hd_a30[6]), .B(d30[6]), .S0(n8663), .Y(n5013) );
  CLKMX2X2 U5706 ( .A(hd_a30[7]), .B(d30[7]), .S0(n8663), .Y(n5012) );
  CLKMX2X2 U5707 ( .A(hd_a30[8]), .B(d30[8]), .S0(n8663), .Y(n5011) );
  CLKMX2X2 U5708 ( .A(hd_a30[9]), .B(d30[9]), .S0(n8663), .Y(n5010) );
  CLKMX2X2 U5709 ( .A(hd_a30[10]), .B(d30[10]), .S0(n8663), .Y(n5009) );
  CLKMX2X2 U5710 ( .A(hd_a30[11]), .B(d30[11]), .S0(n8663), .Y(n5008) );
  CLKMX2X2 U5711 ( .A(hd_a30[12]), .B(d30[12]), .S0(n8663), .Y(n5007) );
  CLKMX2X2 U5712 ( .A(hd_a30[13]), .B(d30[13]), .S0(n8663), .Y(n5006) );
  CLKMX2X2 U5713 ( .A(hd_a30[14]), .B(d30[14]), .S0(n8662), .Y(n5005) );
  CLKMX2X2 U5714 ( .A(hd_a30[15]), .B(d30[15]), .S0(n8662), .Y(n5004) );
  CLKMX2X2 U5715 ( .A(hd_a30[16]), .B(d30[16]), .S0(n8662), .Y(n5003) );
  CLKMX2X2 U5716 ( .A(hd_a30[17]), .B(d30[17]), .S0(n8662), .Y(n5002) );
  CLKMX2X2 U5717 ( .A(hd_a30[18]), .B(d30[18]), .S0(n8662), .Y(n5001) );
  CLKMX2X2 U5718 ( .A(hd_a30[19]), .B(d30[19]), .S0(n8662), .Y(n5000) );
  CLKMX2X2 U5719 ( .A(hd_a30[20]), .B(d30[20]), .S0(n8662), .Y(n4999) );
  CLKMX2X2 U5720 ( .A(hd_a30[21]), .B(d30[21]), .S0(n8662), .Y(n4998) );
  CLKMX2X2 U5721 ( .A(hd_a30[22]), .B(d30[22]), .S0(n8662), .Y(n4997) );
  CLKMX2X2 U5722 ( .A(hd_a30[23]), .B(d30[23]), .S0(n8662), .Y(n4996) );
  CLKMX2X2 U5723 ( .A(hd_a30[24]), .B(d30[24]), .S0(n8662), .Y(n4995) );
  CLKMX2X2 U5724 ( .A(hd_a30[25]), .B(d30[25]), .S0(n8662), .Y(n4994) );
  CLKMX2X2 U5725 ( .A(hd_a30[26]), .B(d30[26]), .S0(n8661), .Y(n4993) );
  CLKMX2X2 U5726 ( .A(hd_a30[27]), .B(d30[27]), .S0(n8661), .Y(n4992) );
  CLKMX2X2 U5727 ( .A(hd_a30[28]), .B(d30[28]), .S0(n8661), .Y(n4991) );
  CLKMX2X2 U5728 ( .A(hd_a30[29]), .B(d30[29]), .S0(n8661), .Y(n4990) );
  CLKMX2X2 U5729 ( .A(hd_a30[30]), .B(d30[30]), .S0(n8661), .Y(n4989) );
  CLKMX2X2 U5730 ( .A(hd_a30[31]), .B(d30[31]), .S0(n8661), .Y(n4988) );
  CLKMX2X2 U5731 ( .A(hd_a30[32]), .B(d30[32]), .S0(n8661), .Y(n4987) );
  CLKMX2X2 U5732 ( .A(hd_a30[33]), .B(d30[33]), .S0(n8661), .Y(n4986) );
  CLKMX2X2 U5733 ( .A(hd_a30[34]), .B(d30[34]), .S0(n8661), .Y(n4985) );
  CLKMX2X2 U5734 ( .A(hd_a30[35]), .B(d30[35]), .S0(n8661), .Y(n4984) );
  CLKMX2X2 U5735 ( .A(hd_a31[0]), .B(d31[0]), .S0(n8661), .Y(n4983) );
  CLKMX2X2 U5736 ( .A(hd_a31[1]), .B(d31[1]), .S0(n8661), .Y(n4982) );
  CLKMX2X2 U5737 ( .A(hd_a31[2]), .B(d31[2]), .S0(n8661), .Y(n4981) );
  CLKMX2X2 U5738 ( .A(hd_a31[3]), .B(d31[3]), .S0(n8660), .Y(n4980) );
  CLKMX2X2 U5739 ( .A(hd_a31[4]), .B(d31[4]), .S0(n8660), .Y(n4979) );
  CLKMX2X2 U5740 ( .A(hd_a31[5]), .B(d31[5]), .S0(n8660), .Y(n4978) );
  CLKMX2X2 U5741 ( .A(hd_a31[6]), .B(d31[6]), .S0(n8660), .Y(n4977) );
  CLKMX2X2 U5742 ( .A(hd_a31[7]), .B(d31[7]), .S0(n8660), .Y(n4976) );
  CLKMX2X2 U5743 ( .A(hd_a31[8]), .B(d31[8]), .S0(n8660), .Y(n4975) );
  CLKMX2X2 U5744 ( .A(hd_a31[9]), .B(d31[9]), .S0(n8660), .Y(n4974) );
  CLKMX2X2 U5745 ( .A(hd_a31[10]), .B(d31[10]), .S0(n8660), .Y(n4973) );
  CLKMX2X2 U5746 ( .A(hd_a31[11]), .B(d31[11]), .S0(n8660), .Y(n4972) );
  CLKMX2X2 U5747 ( .A(hd_a31[12]), .B(d31[12]), .S0(n8660), .Y(n4971) );
  CLKMX2X2 U5748 ( .A(hd_a31[13]), .B(d31[13]), .S0(n8660), .Y(n4970) );
  CLKMX2X2 U5749 ( .A(hd_a31[14]), .B(d31[14]), .S0(n8660), .Y(n4969) );
  CLKMX2X2 U5750 ( .A(hd_a31[15]), .B(d31[15]), .S0(n8660), .Y(n4968) );
  CLKMX2X2 U5751 ( .A(hd_a31[16]), .B(d31[16]), .S0(n8659), .Y(n4967) );
  CLKMX2X2 U5752 ( .A(hd_a31[17]), .B(d31[17]), .S0(n8659), .Y(n4966) );
  CLKMX2X2 U5753 ( .A(hd_a31[18]), .B(d31[18]), .S0(n8659), .Y(n4965) );
  CLKMX2X2 U5754 ( .A(hd_a31[19]), .B(d31[19]), .S0(n8659), .Y(n4964) );
  CLKMX2X2 U5755 ( .A(hd_a31[20]), .B(d31[20]), .S0(n8659), .Y(n4963) );
  CLKMX2X2 U5756 ( .A(hd_a31[21]), .B(d31[21]), .S0(n8659), .Y(n4962) );
  CLKMX2X2 U5757 ( .A(hd_a31[22]), .B(d31[22]), .S0(n8659), .Y(n4961) );
  CLKMX2X2 U5758 ( .A(hd_a31[23]), .B(d31[23]), .S0(n8659), .Y(n4960) );
  CLKMX2X2 U5759 ( .A(hd_a31[24]), .B(d31[24]), .S0(n8659), .Y(n4959) );
  CLKMX2X2 U5760 ( .A(hd_a31[25]), .B(d31[25]), .S0(n8659), .Y(n4958) );
  CLKMX2X2 U5761 ( .A(hd_a31[26]), .B(d31[26]), .S0(n8659), .Y(n4957) );
  CLKMX2X2 U5762 ( .A(hd_a31[27]), .B(d31[27]), .S0(n8659), .Y(n4956) );
  CLKMX2X2 U5763 ( .A(hd_a31[28]), .B(d31[28]), .S0(n8659), .Y(n4955) );
  CLKMX2X2 U5764 ( .A(hd_a31[29]), .B(d31[29]), .S0(n8658), .Y(n4954) );
  CLKMX2X2 U5765 ( .A(hd_a31[30]), .B(d31[30]), .S0(n8658), .Y(n4953) );
  CLKMX2X2 U5766 ( .A(hd_a31[31]), .B(d31[31]), .S0(n8658), .Y(n4952) );
  CLKMX2X2 U5767 ( .A(hd_a32[16]), .B(d32[16]), .S0(n8658), .Y(n4951) );
  CLKMX2X2 U5768 ( .A(hd_a32[17]), .B(d32[17]), .S0(n8658), .Y(n4950) );
  CLKMX2X2 U5769 ( .A(hd_a32[18]), .B(d32[18]), .S0(n8658), .Y(n4949) );
  CLKMX2X2 U5770 ( .A(hd_a32[19]), .B(d32[19]), .S0(n8658), .Y(n4948) );
  CLKMX2X2 U5771 ( .A(hd_a32[20]), .B(d32[20]), .S0(n8658), .Y(n4947) );
  CLKMX2X2 U5772 ( .A(hd_a32[21]), .B(d32[21]), .S0(n8658), .Y(n4946) );
  CLKMX2X2 U5773 ( .A(hd_a32[22]), .B(d32[22]), .S0(n8658), .Y(n4945) );
  CLKMX2X2 U5774 ( .A(hd_a32[23]), .B(d32[23]), .S0(n8658), .Y(n4944) );
  CLKMX2X2 U5775 ( .A(hd_a32[24]), .B(d32[24]), .S0(n8658), .Y(n4943) );
  CLKMX2X2 U5776 ( .A(hd_a32[25]), .B(d32[25]), .S0(n8658), .Y(n4942) );
  CLKMX2X2 U5777 ( .A(hd_a32[26]), .B(d32[26]), .S0(n8657), .Y(n4941) );
  CLKMX2X2 U5778 ( .A(hd_a32[27]), .B(d32[27]), .S0(n8657), .Y(n4940) );
  CLKMX2X2 U5779 ( .A(hd_a32[28]), .B(d32[28]), .S0(n8657), .Y(n4939) );
  CLKMX2X2 U5780 ( .A(hd_a32[29]), .B(d32[29]), .S0(n8657), .Y(n4938) );
  CLKMX2X2 U5781 ( .A(hd_a32[30]), .B(d32[30]), .S0(n8657), .Y(n4937) );
  CLKMX2X2 U5782 ( .A(hd_a32[31]), .B(n11219), .S0(n8662), .Y(n4936) );
  CLKINVX1 U5783 ( .A(n9176), .Y(n4935) );
  AOI222XL U5784 ( .A0(n11221), .A1(n6200), .B0(n9177), .B1(fir_d[0]), .C0(N76), .C1(n9178), .Y(n9176) );
  MXI2X1 U5785 ( .A(n10468), .B(n10469), .S0(n8735), .Y(n4934) );
  MXI2X1 U5786 ( .A(n10467), .B(n10468), .S0(n8750), .Y(n4933) );
  MXI2X1 U5787 ( .A(n10466), .B(n10467), .S0(n8745), .Y(n4932) );
  MXI2X1 U5788 ( .A(n10465), .B(n10466), .S0(n8745), .Y(n4931) );
  MXI2X1 U5789 ( .A(n10464), .B(n10465), .S0(n8745), .Y(n4930) );
  MXI2X1 U5790 ( .A(n10463), .B(n10464), .S0(n8745), .Y(n4929) );
  MXI2X1 U5791 ( .A(n1944), .B(n10463), .S0(n8745), .Y(n4928) );
  CLKINVX1 U5792 ( .A(n9179), .Y(n4927) );
  AOI222XL U5793 ( .A0(n11223), .A1(n6201), .B0(n9177), .B1(fir_d[1]), .C0(N77), .C1(n9178), .Y(n9179) );
  MXI2X1 U5794 ( .A(n10461), .B(n10462), .S0(n8745), .Y(n4926) );
  MXI2X1 U5795 ( .A(n10460), .B(n10461), .S0(n8746), .Y(n4925) );
  MXI2X1 U5796 ( .A(n10459), .B(n10460), .S0(n8746), .Y(n4924) );
  MXI2X1 U5797 ( .A(n10458), .B(n10459), .S0(n8746), .Y(n4923) );
  MXI2X1 U5798 ( .A(n10457), .B(n10458), .S0(n8746), .Y(n4922) );
  MXI2X1 U5799 ( .A(n10456), .B(n10457), .S0(n8746), .Y(n4921) );
  MXI2X1 U5800 ( .A(n1936), .B(n10456), .S0(n8746), .Y(n4920) );
  CLKINVX1 U5801 ( .A(n9180), .Y(n4919) );
  AOI222XL U5802 ( .A0(n11223), .A1(n6202), .B0(n9177), .B1(fir_d[2]), .C0(N78), .C1(n9178), .Y(n9180) );
  MXI2X1 U5803 ( .A(n10454), .B(n10455), .S0(n8746), .Y(n4918) );
  MXI2X1 U5804 ( .A(n10453), .B(n10454), .S0(n8746), .Y(n4917) );
  MXI2X1 U5805 ( .A(n10452), .B(n10453), .S0(n8746), .Y(n4916) );
  MXI2X1 U5806 ( .A(n10451), .B(n10452), .S0(n8746), .Y(n4915) );
  MXI2X1 U5807 ( .A(n10450), .B(n10451), .S0(n8746), .Y(n4914) );
  MXI2X1 U5808 ( .A(n10449), .B(n10450), .S0(n8746), .Y(n4913) );
  MXI2X1 U5809 ( .A(n1928), .B(n10449), .S0(n8746), .Y(n4912) );
  CLKINVX1 U5810 ( .A(n9181), .Y(n4911) );
  AOI222XL U5811 ( .A0(n11216), .A1(n6203), .B0(n9177), .B1(fir_d[3]), .C0(N79), .C1(n9178), .Y(n9181) );
  MXI2X1 U5812 ( .A(n10447), .B(n10448), .S0(n8747), .Y(n4910) );
  MXI2X1 U5813 ( .A(n10446), .B(n10447), .S0(n8747), .Y(n4909) );
  MXI2X1 U5814 ( .A(n10445), .B(n10446), .S0(n8747), .Y(n4908) );
  MXI2X1 U5815 ( .A(n10444), .B(n10445), .S0(n8747), .Y(n4907) );
  MXI2X1 U5816 ( .A(n10443), .B(n10444), .S0(n8747), .Y(n4906) );
  MXI2X1 U5817 ( .A(n10442), .B(n10443), .S0(n8747), .Y(n4905) );
  MXI2X1 U5818 ( .A(n1920), .B(n10442), .S0(n8747), .Y(n4904) );
  CLKINVX1 U5819 ( .A(n9182), .Y(n4903) );
  AOI222XL U5820 ( .A0(n11222), .A1(n6204), .B0(n9177), .B1(fir_d[4]), .C0(N80), .C1(n9178), .Y(n9182) );
  MXI2X1 U5821 ( .A(n10440), .B(n10441), .S0(n8747), .Y(n4902) );
  MXI2X1 U5822 ( .A(n10439), .B(n10440), .S0(n8747), .Y(n4901) );
  MXI2X1 U5823 ( .A(n10438), .B(n10439), .S0(n8747), .Y(n4900) );
  MXI2X1 U5824 ( .A(n10437), .B(n10438), .S0(n8747), .Y(n4899) );
  MXI2X1 U5825 ( .A(n10436), .B(n10437), .S0(n8747), .Y(n4898) );
  MXI2X1 U5826 ( .A(n10435), .B(n10436), .S0(n8747), .Y(n4897) );
  MXI2X1 U5827 ( .A(n1912), .B(n10435), .S0(n8748), .Y(n4896) );
  CLKINVX1 U5828 ( .A(n9183), .Y(n4895) );
  AOI222XL U5829 ( .A0(n11224), .A1(n6205), .B0(n9177), .B1(fir_d[5]), .C0(N81), .C1(n9178), .Y(n9183) );
  MXI2X1 U5830 ( .A(n10433), .B(n10434), .S0(n8748), .Y(n4894) );
  MXI2X1 U5831 ( .A(n10432), .B(n10433), .S0(n8748), .Y(n4893) );
  MXI2X1 U5832 ( .A(n10431), .B(n10432), .S0(n8748), .Y(n4892) );
  MXI2X1 U5833 ( .A(n10430), .B(n10431), .S0(n8748), .Y(n4891) );
  MXI2X1 U5834 ( .A(n10429), .B(n10430), .S0(n8748), .Y(n4890) );
  MXI2X1 U5835 ( .A(n10428), .B(n10429), .S0(n8748), .Y(n4889) );
  MXI2X1 U5836 ( .A(n1904), .B(n10428), .S0(n8748), .Y(n4888) );
  CLKINVX1 U5837 ( .A(n9184), .Y(n4887) );
  AOI222XL U5838 ( .A0(n11224), .A1(n6206), .B0(n9177), .B1(fir_d[6]), .C0(N82), .C1(n9178), .Y(n9184) );
  MXI2X1 U5839 ( .A(n10426), .B(n10427), .S0(n8748), .Y(n4886) );
  MXI2X1 U5840 ( .A(n10425), .B(n10426), .S0(n8748), .Y(n4885) );
  MXI2X1 U5841 ( .A(n10424), .B(n10425), .S0(n8748), .Y(n4884) );
  MXI2X1 U5842 ( .A(n10423), .B(n10424), .S0(n8748), .Y(n4883) );
  MXI2X1 U5843 ( .A(n10422), .B(n10423), .S0(n8748), .Y(n4882) );
  MXI2X1 U5844 ( .A(n10421), .B(n10422), .S0(n8749), .Y(n4881) );
  MXI2X1 U5845 ( .A(n1896), .B(n10421), .S0(n8749), .Y(n4880) );
  CLKINVX1 U5846 ( .A(n9185), .Y(n4879) );
  AOI222XL U5847 ( .A0(n11215), .A1(n6207), .B0(n9177), .B1(fir_d[7]), .C0(N83), .C1(n9178), .Y(n9185) );
  MXI2X1 U5848 ( .A(n10419), .B(n10420), .S0(n8749), .Y(n4878) );
  MXI2X1 U5849 ( .A(n10418), .B(n10419), .S0(n8749), .Y(n4877) );
  MXI2X1 U5850 ( .A(n10417), .B(n10418), .S0(n8749), .Y(n4876) );
  MXI2X1 U5851 ( .A(n10416), .B(n10417), .S0(n8749), .Y(n4875) );
  MXI2X1 U5852 ( .A(n10415), .B(n10416), .S0(n8749), .Y(n4874) );
  MXI2X1 U5853 ( .A(n10414), .B(n10415), .S0(n8749), .Y(n4873) );
  MXI2X1 U5854 ( .A(n1888), .B(n10414), .S0(n8749), .Y(n4872) );
  CLKINVX1 U5855 ( .A(n9186), .Y(n4871) );
  AOI222XL U5856 ( .A0(n11221), .A1(n6208), .B0(n9177), .B1(fir_d[8]), .C0(N84), .C1(n9178), .Y(n9186) );
  MXI2X1 U5857 ( .A(n10412), .B(n10413), .S0(n8749), .Y(n4870) );
  MXI2X1 U5858 ( .A(n10411), .B(n10412), .S0(n8749), .Y(n4869) );
  MXI2X1 U5859 ( .A(n10410), .B(n10411), .S0(n8749), .Y(n4868) );
  MXI2X1 U5860 ( .A(n10409), .B(n10410), .S0(n8749), .Y(n4867) );
  MXI2X1 U5861 ( .A(n10408), .B(n10409), .S0(n8750), .Y(n4866) );
  MXI2X1 U5862 ( .A(n10407), .B(n10408), .S0(n8750), .Y(n4865) );
  MXI2X1 U5863 ( .A(n1880), .B(n10407), .S0(n8750), .Y(n4864) );
  CLKINVX1 U5864 ( .A(n9187), .Y(n4863) );
  AOI222XL U5865 ( .A0(n11221), .A1(n6209), .B0(n9177), .B1(fir_d[9]), .C0(N85), .C1(n9178), .Y(n9187) );
  MXI2X1 U5866 ( .A(n10405), .B(n10406), .S0(n8750), .Y(n4862) );
  MXI2X1 U5867 ( .A(n10404), .B(n10405), .S0(n8750), .Y(n4861) );
  MXI2X1 U5868 ( .A(n10403), .B(n10404), .S0(n8750), .Y(n4860) );
  MXI2X1 U5869 ( .A(n10402), .B(n10403), .S0(n8755), .Y(n4859) );
  MXI2X1 U5870 ( .A(n10401), .B(n10402), .S0(n8755), .Y(n4858) );
  MXI2X1 U5871 ( .A(n10400), .B(n10401), .S0(n8755), .Y(n4857) );
  MXI2X1 U5872 ( .A(n1872), .B(n10400), .S0(n8735), .Y(n4856) );
  CLKINVX1 U5873 ( .A(n9188), .Y(n4855) );
  AOI222XL U5874 ( .A0(n11221), .A1(n6210), .B0(n9177), .B1(fir_d[10]), .C0(
        N86), .C1(n9178), .Y(n9188) );
  MXI2X1 U5875 ( .A(n10398), .B(n10399), .S0(n8735), .Y(n4854) );
  MXI2X1 U5876 ( .A(n10397), .B(n10398), .S0(n8735), .Y(n4853) );
  MXI2X1 U5877 ( .A(n10396), .B(n10397), .S0(n8735), .Y(n4852) );
  MXI2X1 U5878 ( .A(n10395), .B(n10396), .S0(n8736), .Y(n4851) );
  MXI2X1 U5879 ( .A(n10394), .B(n10395), .S0(n8736), .Y(n4850) );
  MXI2X1 U5880 ( .A(n10393), .B(n10394), .S0(n8736), .Y(n4849) );
  MXI2X1 U5881 ( .A(n1864), .B(n10393), .S0(n8737), .Y(n4848) );
  CLKINVX1 U5882 ( .A(n9189), .Y(n4847) );
  AOI222XL U5883 ( .A0(n11216), .A1(n6211), .B0(n9177), .B1(fir_d[11]), .C0(
        N87), .C1(n9178), .Y(n9189) );
  MXI2X1 U5884 ( .A(n10391), .B(n10392), .S0(n8737), .Y(n4846) );
  MXI2X1 U5885 ( .A(n10390), .B(n10391), .S0(n8737), .Y(n4845) );
  MXI2X1 U5886 ( .A(n10389), .B(n10390), .S0(n8738), .Y(n4844) );
  MXI2X1 U5887 ( .A(n10388), .B(n10389), .S0(n8738), .Y(n4843) );
  MXI2X1 U5888 ( .A(n10387), .B(n10388), .S0(n8738), .Y(n4842) );
  MXI2X1 U5889 ( .A(n10386), .B(n10387), .S0(n8739), .Y(n4841) );
  MXI2X1 U5890 ( .A(n1856), .B(n10386), .S0(n8739), .Y(n4840) );
  CLKINVX1 U5891 ( .A(n9190), .Y(n4839) );
  AOI222XL U5892 ( .A0(n11222), .A1(n6212), .B0(n9177), .B1(fir_d[12]), .C0(
        N88), .C1(n9178), .Y(n9190) );
  MXI2X1 U5893 ( .A(n10384), .B(n10385), .S0(n8739), .Y(n4838) );
  MXI2X1 U5894 ( .A(n10383), .B(n10384), .S0(n8739), .Y(n4837) );
  MXI2X1 U5895 ( .A(n10382), .B(n10383), .S0(n8740), .Y(n4836) );
  MXI2X1 U5896 ( .A(n10381), .B(n10382), .S0(n8740), .Y(n4835) );
  MXI2X1 U5897 ( .A(n10380), .B(n10381), .S0(n8740), .Y(n4834) );
  MXI2X1 U5898 ( .A(n10379), .B(n10380), .S0(n8741), .Y(n4833) );
  MXI2X1 U5899 ( .A(n1848), .B(n10379), .S0(n8741), .Y(n4832) );
  CLKINVX1 U5900 ( .A(n9191), .Y(n4831) );
  AOI222XL U5901 ( .A0(n11222), .A1(n6213), .B0(n9177), .B1(fir_d[13]), .C0(
        N89), .C1(n9178), .Y(n9191) );
  MXI2X1 U5902 ( .A(n10377), .B(n10378), .S0(n8741), .Y(n4830) );
  MXI2X1 U5903 ( .A(n10376), .B(n10377), .S0(n8742), .Y(n4829) );
  MXI2X1 U5904 ( .A(n10375), .B(n10376), .S0(n8742), .Y(n4828) );
  MXI2X1 U5905 ( .A(n10374), .B(n10375), .S0(n8742), .Y(n4827) );
  MXI2X1 U5906 ( .A(n10373), .B(n10374), .S0(n8743), .Y(n4826) );
  MXI2X1 U5907 ( .A(n10372), .B(n10373), .S0(n8743), .Y(n4825) );
  MXI2X1 U5908 ( .A(n1840), .B(n10372), .S0(n8743), .Y(n4824) );
  CLKINVX1 U5909 ( .A(n9192), .Y(n4823) );
  AOI222XL U5910 ( .A0(n11222), .A1(n6214), .B0(n9177), .B1(fir_d[14]), .C0(
        N90), .C1(n9178), .Y(n9192) );
  MXI2X1 U5911 ( .A(n10370), .B(n10371), .S0(n8744), .Y(n4822) );
  MXI2X1 U5912 ( .A(n10369), .B(n10370), .S0(n8744), .Y(n4821) );
  MXI2X1 U5913 ( .A(n10368), .B(n10369), .S0(n8744), .Y(n4820) );
  MXI2X1 U5914 ( .A(n10367), .B(n10368), .S0(n8745), .Y(n4819) );
  MXI2X1 U5915 ( .A(n10366), .B(n10367), .S0(n8745), .Y(n4818) );
  MXI2X1 U5916 ( .A(n10365), .B(n10366), .S0(n8745), .Y(n4817) );
  MXI2X1 U5917 ( .A(n1832), .B(n10365), .S0(n8745), .Y(n4816) );
  CLKINVX1 U5918 ( .A(n9193), .Y(n4815) );
  AOI222XL U5919 ( .A0(n11215), .A1(n6215), .B0(fir_d[15]), .B1(n9177), .C0(
        N91), .C1(n9178), .Y(n9193) );
  NOR2X1 U5920 ( .A(n11222), .B(n11212), .Y(n9178) );
  NOR2X1 U5921 ( .A(n6192), .B(n11215), .Y(n9177) );
  MXI2X1 U5922 ( .A(n10363), .B(n10364), .S0(n8745), .Y(n4814) );
  MXI2X1 U5923 ( .A(n10362), .B(n10363), .S0(n8745), .Y(n4813) );
  MXI2X1 U5924 ( .A(n10361), .B(n10362), .S0(n8745), .Y(n4812) );
  MXI2X1 U5925 ( .A(n10360), .B(n10361), .S0(n8744), .Y(n4811) );
  MXI2X1 U5926 ( .A(n10359), .B(n10360), .S0(n8744), .Y(n4810) );
  MXI2X1 U5927 ( .A(n10358), .B(n10359), .S0(n8744), .Y(n4809) );
  MXI2X1 U5928 ( .A(n1824), .B(n10358), .S0(n8744), .Y(n4808) );
  OAI222XL U5929 ( .A0(n6094), .A1(n9194), .B0(n9195), .B1(n9196), .C0(n10357), 
        .C1(n8759), .Y(n4807) );
  MXI2X1 U5930 ( .A(n10356), .B(n10357), .S0(n8744), .Y(n4806) );
  MXI2X1 U5931 ( .A(n10355), .B(n10356), .S0(n8744), .Y(n4805) );
  MXI2X1 U5932 ( .A(n6094), .B(n10355), .S0(n8744), .Y(n4804) );
  OAI221XL U5933 ( .A0(n9197), .A1(n9198), .B0(n6110), .B1(n9195), .C0(n9199), 
        .Y(n4803) );
  OA22X1 U5934 ( .A0(n9194), .A1(n9196), .B0(n8759), .B1(n10354), .Y(n9199) );
  CLKINVX1 U5935 ( .A(N97), .Y(n9196) );
  MXI2X1 U5936 ( .A(n10353), .B(n10354), .S0(n8744), .Y(n4802) );
  MXI2X1 U5937 ( .A(n10352), .B(n10353), .S0(n8744), .Y(n4801) );
  MXI2X1 U5938 ( .A(n6110), .B(n10352), .S0(n8744), .Y(n4800) );
  OAI221XL U5939 ( .A0(n9197), .A1(n9200), .B0(n6109), .B1(n9195), .C0(n9201), 
        .Y(n4799) );
  OA22X1 U5940 ( .A0(n9202), .A1(n9194), .B0(n8759), .B1(n10351), .Y(n9201) );
  MXI2X1 U5941 ( .A(n10350), .B(n10351), .S0(n8743), .Y(n4798) );
  MXI2X1 U5942 ( .A(n10349), .B(n10350), .S0(n8743), .Y(n4797) );
  MXI2X1 U5943 ( .A(n6109), .B(n10349), .S0(n8743), .Y(n4796) );
  OAI222XL U5944 ( .A0(n6093), .A1(n9194), .B0(n9195), .B1(n9202), .C0(n10348), 
        .C1(n8759), .Y(n4795) );
  CLKINVX1 U5945 ( .A(N98), .Y(n9202) );
  MXI2X1 U5946 ( .A(n10347), .B(n10348), .S0(n8743), .Y(n4794) );
  MXI2X1 U5947 ( .A(n10346), .B(n10347), .S0(n8743), .Y(n4793) );
  MXI2X1 U5948 ( .A(n6093), .B(n10346), .S0(n8743), .Y(n4792) );
  OAI221XL U5949 ( .A0(n9197), .A1(n9203), .B0(n6108), .B1(n9195), .C0(n9204), 
        .Y(n4791) );
  OA22X1 U5950 ( .A0(n9205), .A1(n9194), .B0(n8759), .B1(n10345), .Y(n9204) );
  MXI2X1 U5951 ( .A(n10344), .B(n10345), .S0(n8743), .Y(n4790) );
  MXI2X1 U5952 ( .A(n10343), .B(n10344), .S0(n8743), .Y(n4789) );
  MXI2X1 U5953 ( .A(n6108), .B(n10343), .S0(n8743), .Y(n4788) );
  OAI222XL U5954 ( .A0(n6092), .A1(n9194), .B0(n9195), .B1(n9205), .C0(n10342), 
        .C1(n8759), .Y(n4787) );
  CLKINVX1 U5955 ( .A(N99), .Y(n9205) );
  MXI2X1 U5956 ( .A(n10341), .B(n10342), .S0(n8743), .Y(n4786) );
  MXI2X1 U5957 ( .A(n10340), .B(n10341), .S0(n8742), .Y(n4785) );
  MXI2X1 U5958 ( .A(n6092), .B(n10340), .S0(n8742), .Y(n4784) );
  OAI221XL U5959 ( .A0(n9197), .A1(n9206), .B0(n6107), .B1(n9195), .C0(n9207), 
        .Y(n4783) );
  OA22X1 U5960 ( .A0(n9208), .A1(n9194), .B0(n8759), .B1(n10339), .Y(n9207) );
  MXI2X1 U5961 ( .A(n10338), .B(n10339), .S0(n8742), .Y(n4782) );
  MXI2X1 U5962 ( .A(n10337), .B(n10338), .S0(n8742), .Y(n4781) );
  MXI2X1 U5963 ( .A(n6107), .B(n10337), .S0(n8742), .Y(n4780) );
  OAI222XL U5964 ( .A0(n6091), .A1(n9194), .B0(n9195), .B1(n9208), .C0(n10336), 
        .C1(n8759), .Y(n4779) );
  CLKINVX1 U5965 ( .A(N100), .Y(n9208) );
  MXI2X1 U5966 ( .A(n10335), .B(n10336), .S0(n8742), .Y(n4778) );
  MXI2X1 U5967 ( .A(n10334), .B(n10335), .S0(n8742), .Y(n4777) );
  MXI2X1 U5968 ( .A(n6091), .B(n10334), .S0(n8742), .Y(n4776) );
  OAI221XL U5969 ( .A0(n9197), .A1(n9209), .B0(n6106), .B1(n9195), .C0(n9210), 
        .Y(n4775) );
  OA22X1 U5970 ( .A0(n9211), .A1(n9194), .B0(n8759), .B1(n10333), .Y(n9210) );
  MXI2X1 U5971 ( .A(n10332), .B(n10333), .S0(n8742), .Y(n4774) );
  MXI2X1 U5972 ( .A(n10331), .B(n10332), .S0(n8742), .Y(n4773) );
  MXI2X1 U5973 ( .A(n6106), .B(n10331), .S0(n8741), .Y(n4772) );
  OAI222XL U5974 ( .A0(n6090), .A1(n9194), .B0(n9195), .B1(n9211), .C0(n10330), 
        .C1(n8759), .Y(n4771) );
  CLKINVX1 U5975 ( .A(N101), .Y(n9211) );
  MXI2X1 U5976 ( .A(n10329), .B(n10330), .S0(n8741), .Y(n4770) );
  MXI2X1 U5977 ( .A(n10328), .B(n10329), .S0(n8741), .Y(n4769) );
  MXI2X1 U5978 ( .A(n6090), .B(n10328), .S0(n8741), .Y(n4768) );
  OAI221XL U5979 ( .A0(n9197), .A1(n9212), .B0(n6105), .B1(n9195), .C0(n9213), 
        .Y(n4767) );
  OA22X1 U5980 ( .A0(n9214), .A1(n9194), .B0(n8759), .B1(n10327), .Y(n9213) );
  MXI2X1 U5981 ( .A(n10326), .B(n10327), .S0(n8741), .Y(n4766) );
  MXI2X1 U5982 ( .A(n10325), .B(n10326), .S0(n8741), .Y(n4765) );
  MXI2X1 U5983 ( .A(n6105), .B(n10325), .S0(n8741), .Y(n4764) );
  OAI222XL U5984 ( .A0(n6089), .A1(n9194), .B0(n9195), .B1(n9214), .C0(n10324), 
        .C1(n8759), .Y(n4763) );
  CLKINVX1 U5985 ( .A(N102), .Y(n9214) );
  MXI2X1 U5986 ( .A(n10323), .B(n10324), .S0(n8741), .Y(n4762) );
  MXI2X1 U5987 ( .A(n10322), .B(n10323), .S0(n8741), .Y(n4761) );
  MXI2X1 U5988 ( .A(n6089), .B(n10322), .S0(n8741), .Y(n4760) );
  OAI221XL U5989 ( .A0(n9197), .A1(n9215), .B0(n6104), .B1(n9195), .C0(n9216), 
        .Y(n4759) );
  OA22X1 U5990 ( .A0(n9217), .A1(n9194), .B0(n8759), .B1(n10321), .Y(n9216) );
  MXI2X1 U5991 ( .A(n10320), .B(n10321), .S0(n8740), .Y(n4758) );
  MXI2X1 U5992 ( .A(n10319), .B(n10320), .S0(n8740), .Y(n4757) );
  MXI2X1 U5993 ( .A(n6104), .B(n10319), .S0(n8740), .Y(n4756) );
  OAI222XL U5994 ( .A0(n6088), .A1(n9194), .B0(n9195), .B1(n9217), .C0(n10318), 
        .C1(n8759), .Y(n4755) );
  CLKINVX1 U5995 ( .A(N103), .Y(n9217) );
  MXI2X1 U5996 ( .A(n10317), .B(n10318), .S0(n8740), .Y(n4754) );
  MXI2X1 U5997 ( .A(n10316), .B(n10317), .S0(n8740), .Y(n4753) );
  MXI2X1 U5998 ( .A(n6088), .B(n10316), .S0(n8740), .Y(n4752) );
  OAI221XL U5999 ( .A0(n9197), .A1(n9218), .B0(n6103), .B1(n9195), .C0(n9219), 
        .Y(n4751) );
  OA22X1 U6000 ( .A0(n9220), .A1(n9194), .B0(n8759), .B1(n10315), .Y(n9219) );
  MXI2X1 U6001 ( .A(n10314), .B(n10315), .S0(n8740), .Y(n4750) );
  MXI2X1 U6002 ( .A(n10313), .B(n10314), .S0(n8740), .Y(n4749) );
  MXI2X1 U6003 ( .A(n6103), .B(n10313), .S0(n8740), .Y(n4748) );
  OAI222XL U6004 ( .A0(n6087), .A1(n9194), .B0(n9195), .B1(n9220), .C0(n10312), 
        .C1(n8758), .Y(n4747) );
  CLKINVX1 U6005 ( .A(N104), .Y(n9220) );
  MXI2X1 U6006 ( .A(n10311), .B(n10312), .S0(n8739), .Y(n4746) );
  MXI2X1 U6007 ( .A(n10310), .B(n10311), .S0(n8739), .Y(n4745) );
  MXI2X1 U6008 ( .A(n6087), .B(n10310), .S0(n8739), .Y(n4744) );
  OAI221XL U6009 ( .A0(n9197), .A1(n9221), .B0(n6102), .B1(n9195), .C0(n9222), 
        .Y(n4743) );
  OA22X1 U6010 ( .A0(n9223), .A1(n9194), .B0(n8759), .B1(n10309), .Y(n9222) );
  MXI2X1 U6011 ( .A(n10308), .B(n10309), .S0(n8739), .Y(n4742) );
  MXI2X1 U6012 ( .A(n10307), .B(n10308), .S0(n8739), .Y(n4741) );
  MXI2X1 U6013 ( .A(n6102), .B(n10307), .S0(n8739), .Y(n4740) );
  OAI222XL U6014 ( .A0(n6086), .A1(n9194), .B0(n9195), .B1(n9223), .C0(n10306), 
        .C1(n8759), .Y(n4739) );
  CLKINVX1 U6015 ( .A(N105), .Y(n9223) );
  MXI2X1 U6016 ( .A(n10305), .B(n10306), .S0(n8739), .Y(n4738) );
  MXI2X1 U6017 ( .A(n10304), .B(n10305), .S0(n8739), .Y(n4737) );
  MXI2X1 U6018 ( .A(n6086), .B(n10304), .S0(n8739), .Y(n4736) );
  OAI221XL U6019 ( .A0(n9197), .A1(n9224), .B0(n6101), .B1(n9195), .C0(n9225), 
        .Y(n4735) );
  OA22X1 U6020 ( .A0(n9226), .A1(n9194), .B0(n8759), .B1(n10303), .Y(n9225) );
  MXI2X1 U6021 ( .A(n10302), .B(n10303), .S0(n8738), .Y(n4734) );
  MXI2X1 U6022 ( .A(n10301), .B(n10302), .S0(n8738), .Y(n4733) );
  MXI2X1 U6023 ( .A(n6101), .B(n10301), .S0(n8738), .Y(n4732) );
  OAI222XL U6024 ( .A0(n6085), .A1(n9194), .B0(n9195), .B1(n9226), .C0(n10300), 
        .C1(n8759), .Y(n4731) );
  CLKINVX1 U6025 ( .A(N106), .Y(n9226) );
  MXI2X1 U6026 ( .A(n10299), .B(n10300), .S0(n8738), .Y(n4730) );
  MXI2X1 U6027 ( .A(n10298), .B(n10299), .S0(n8738), .Y(n4729) );
  MXI2X1 U6028 ( .A(n6085), .B(n10298), .S0(n8738), .Y(n4728) );
  OAI221XL U6029 ( .A0(n9197), .A1(n9227), .B0(n6100), .B1(n9195), .C0(n9228), 
        .Y(n4727) );
  OA22X1 U6030 ( .A0(n9229), .A1(n9194), .B0(n8759), .B1(n10297), .Y(n9228) );
  MXI2X1 U6031 ( .A(n10296), .B(n10297), .S0(n8738), .Y(n4726) );
  MXI2X1 U6032 ( .A(n10295), .B(n10296), .S0(n8738), .Y(n4725) );
  MXI2X1 U6033 ( .A(n6100), .B(n10295), .S0(n8738), .Y(n4724) );
  OAI222XL U6034 ( .A0(n6084), .A1(n9194), .B0(n9195), .B1(n9229), .C0(n10294), 
        .C1(n8759), .Y(n4723) );
  CLKINVX1 U6035 ( .A(N107), .Y(n9229) );
  MXI2X1 U6036 ( .A(n10293), .B(n10294), .S0(n8738), .Y(n4722) );
  MXI2X1 U6037 ( .A(n10292), .B(n10293), .S0(n8737), .Y(n4721) );
  MXI2X1 U6038 ( .A(n6084), .B(n10292), .S0(n8737), .Y(n4720) );
  OAI221XL U6039 ( .A0(n9197), .A1(n9230), .B0(n6099), .B1(n9195), .C0(n9231), 
        .Y(n4719) );
  OA22X1 U6040 ( .A0(n9232), .A1(n9194), .B0(n8759), .B1(n10291), .Y(n9231) );
  MXI2X1 U6041 ( .A(n10290), .B(n10291), .S0(n8737), .Y(n4718) );
  MXI2X1 U6042 ( .A(n10289), .B(n10290), .S0(n8737), .Y(n4717) );
  MXI2X1 U6043 ( .A(n6099), .B(n10289), .S0(n8737), .Y(n4716) );
  OAI222XL U6044 ( .A0(n6083), .A1(n9194), .B0(n9195), .B1(n9232), .C0(n10288), 
        .C1(n8759), .Y(n4715) );
  CLKINVX1 U6045 ( .A(N108), .Y(n9232) );
  MXI2X1 U6046 ( .A(n10287), .B(n10288), .S0(n8737), .Y(n4714) );
  MXI2X1 U6047 ( .A(n10286), .B(n10287), .S0(n8737), .Y(n4713) );
  MXI2X1 U6048 ( .A(n6083), .B(n10286), .S0(n8737), .Y(n4712) );
  OAI221XL U6049 ( .A0(n9197), .A1(n9233), .B0(n6098), .B1(n9195), .C0(n9234), 
        .Y(n4711) );
  OA22X1 U6050 ( .A0(n9235), .A1(n9194), .B0(n8759), .B1(n10285), .Y(n9234) );
  MXI2X1 U6051 ( .A(n10284), .B(n10285), .S0(n8737), .Y(n4710) );
  MXI2X1 U6052 ( .A(n10283), .B(n10284), .S0(n8737), .Y(n4709) );
  MXI2X1 U6053 ( .A(n6098), .B(n10283), .S0(n8736), .Y(n4708) );
  OAI222XL U6054 ( .A0(n6082), .A1(n9194), .B0(n9195), .B1(n9235), .C0(n10282), 
        .C1(n8758), .Y(n4707) );
  CLKINVX1 U6055 ( .A(N109), .Y(n9235) );
  MXI2X1 U6056 ( .A(n10281), .B(n10282), .S0(n8736), .Y(n4706) );
  MXI2X1 U6057 ( .A(n10280), .B(n10281), .S0(n8736), .Y(n4705) );
  MXI2X1 U6058 ( .A(n6082), .B(n10280), .S0(n8736), .Y(n4704) );
  OAI221XL U6059 ( .A0(n9197), .A1(n9236), .B0(n6097), .B1(n9195), .C0(n9237), 
        .Y(n4703) );
  OA22X1 U6060 ( .A0(n9238), .A1(n9194), .B0(n8759), .B1(n10279), .Y(n9237) );
  MXI2X1 U6061 ( .A(n10278), .B(n10279), .S0(n8736), .Y(n4702) );
  MXI2X1 U6062 ( .A(n10277), .B(n10278), .S0(n8736), .Y(n4701) );
  MXI2X1 U6063 ( .A(n6097), .B(n10277), .S0(n8736), .Y(n4700) );
  OAI222XL U6064 ( .A0(n6081), .A1(n9194), .B0(n9195), .B1(n9238), .C0(n10276), 
        .C1(n8758), .Y(n4699) );
  CLKINVX1 U6065 ( .A(N110), .Y(n9238) );
  MXI2X1 U6066 ( .A(n10275), .B(n10276), .S0(n8736), .Y(n4698) );
  MXI2X1 U6067 ( .A(n10274), .B(n10275), .S0(n8736), .Y(n4697) );
  MXI2X1 U6068 ( .A(n6081), .B(n10274), .S0(n8736), .Y(n4696) );
  OAI221XL U6069 ( .A0(n9197), .A1(n9239), .B0(n6096), .B1(n9195), .C0(n9240), 
        .Y(n4695) );
  OA22X1 U6070 ( .A0(n9241), .A1(n9194), .B0(n8759), .B1(n10273), .Y(n9240) );
  MXI2X1 U6071 ( .A(n10272), .B(n10273), .S0(n8735), .Y(n4694) );
  MXI2X1 U6072 ( .A(n10271), .B(n10272), .S0(n8735), .Y(n4693) );
  MXI2X1 U6073 ( .A(n6096), .B(n10271), .S0(n8735), .Y(n4692) );
  OAI222XL U6074 ( .A0(n6080), .A1(n9194), .B0(n9195), .B1(n9241), .C0(n10270), 
        .C1(n8758), .Y(n4691) );
  CLKINVX1 U6075 ( .A(N111), .Y(n9241) );
  MXI2X1 U6076 ( .A(n10269), .B(n10270), .S0(n8735), .Y(n4690) );
  MXI2X1 U6077 ( .A(n10268), .B(n10269), .S0(n8735), .Y(n4689) );
  MXI2X1 U6078 ( .A(n6080), .B(n10268), .S0(n8735), .Y(n4688) );
  OAI221XL U6079 ( .A0(n9197), .A1(n9242), .B0(n6095), .B1(n9195), .C0(n9243), 
        .Y(n4687) );
  OA22X1 U6080 ( .A0(n9244), .A1(n9194), .B0(n8759), .B1(n10267), .Y(n9243) );
  NAND3X1 U6081 ( .A(n9245), .B(n8756), .C(n9246), .Y(n9197) );
  MXI2X1 U6082 ( .A(n10266), .B(n10267), .S0(n8735), .Y(n4686) );
  MXI2X1 U6083 ( .A(n10265), .B(n10266), .S0(n8735), .Y(n4685) );
  MXI2X1 U6084 ( .A(n6095), .B(n10265), .S0(n8740), .Y(n4684) );
  OAI222XL U6085 ( .A0(n6079), .A1(n9194), .B0(n9195), .B1(n9244), .C0(n10264), 
        .C1(n8758), .Y(n4683) );
  CLKINVX1 U6086 ( .A(N112), .Y(n9244) );
  NAND2X1 U6087 ( .A(n9247), .B(n8756), .Y(n9195) );
  NAND2X1 U6088 ( .A(mult_add_355_aco_b), .B(n8756), .Y(n9194) );
  MXI2X1 U6089 ( .A(n10263), .B(n10264), .S0(n8755), .Y(n4682) );
  MXI2X1 U6090 ( .A(n10262), .B(n10263), .S0(n8755), .Y(n4681) );
  MXI2X1 U6091 ( .A(n6079), .B(n10262), .S0(n8755), .Y(n4680) );
  CLKINVX1 U6092 ( .A(n9248), .Y(n4679) );
  AOI222XL U6093 ( .A0(n11223), .A1(n6216), .B0(result_r[0]), .B1(n9249), .C0(
        N300), .C1(n9250), .Y(n9248) );
  MXI2X1 U6094 ( .A(n1725), .B(n10261), .S0(n8755), .Y(n4678) );
  CLKINVX1 U6095 ( .A(n9251), .Y(n4677) );
  AOI222XL U6096 ( .A0(n11223), .A1(n6217), .B0(result_r[1]), .B1(n9249), .C0(
        N301), .C1(n9250), .Y(n9251) );
  MXI2X1 U6097 ( .A(n1723), .B(n10260), .S0(n8755), .Y(n4676) );
  CLKINVX1 U6098 ( .A(n9252), .Y(n4675) );
  AOI222XL U6099 ( .A0(n11223), .A1(n6218), .B0(result_r[2]), .B1(n9249), .C0(
        N302), .C1(n9250), .Y(n9252) );
  MXI2X1 U6100 ( .A(n1721), .B(n10259), .S0(n8755), .Y(n4674) );
  CLKINVX1 U6101 ( .A(n9253), .Y(n4673) );
  AOI222XL U6102 ( .A0(n11216), .A1(n6219), .B0(result_r[3]), .B1(n9249), .C0(
        N303), .C1(n9250), .Y(n9253) );
  MXI2X1 U6103 ( .A(n1719), .B(n10258), .S0(n8755), .Y(n4672) );
  CLKINVX1 U6104 ( .A(n9254), .Y(n4671) );
  AOI222XL U6105 ( .A0(n11224), .A1(n6220), .B0(result_r[4]), .B1(n9249), .C0(
        N304), .C1(n9250), .Y(n9254) );
  MXI2X1 U6106 ( .A(n1717), .B(n10257), .S0(n8755), .Y(n4670) );
  CLKINVX1 U6107 ( .A(n9255), .Y(n4669) );
  AOI222XL U6108 ( .A0(n11224), .A1(n6221), .B0(result_r[5]), .B1(n9249), .C0(
        N305), .C1(n9250), .Y(n9255) );
  MXI2X1 U6109 ( .A(n1715), .B(n10256), .S0(n8755), .Y(n4668) );
  CLKINVX1 U6110 ( .A(n9256), .Y(n4667) );
  AOI222XL U6111 ( .A0(n11224), .A1(n6222), .B0(result_r[6]), .B1(n9249), .C0(
        N306), .C1(n9250), .Y(n9256) );
  MXI2X1 U6112 ( .A(n1713), .B(n10255), .S0(n8754), .Y(n4666) );
  CLKINVX1 U6113 ( .A(n9257), .Y(n4665) );
  AOI222XL U6114 ( .A0(n11215), .A1(n6223), .B0(result_r[7]), .B1(n9249), .C0(
        N307), .C1(n9250), .Y(n9257) );
  MXI2X1 U6115 ( .A(n1711), .B(n10254), .S0(n8754), .Y(n4664) );
  CLKINVX1 U6116 ( .A(n9258), .Y(n4663) );
  AOI222XL U6117 ( .A0(n11221), .A1(n6224), .B0(result_r[8]), .B1(n9249), .C0(
        N308), .C1(n9250), .Y(n9258) );
  MXI2X1 U6118 ( .A(n1709), .B(n10253), .S0(n8754), .Y(n4662) );
  CLKINVX1 U6119 ( .A(n9259), .Y(n4661) );
  AOI222XL U6120 ( .A0(n11221), .A1(n6225), .B0(result_r[9]), .B1(n9249), .C0(
        N309), .C1(n9250), .Y(n9259) );
  MXI2X1 U6121 ( .A(n1707), .B(n10252), .S0(n8754), .Y(n4660) );
  CLKINVX1 U6122 ( .A(n9260), .Y(n4659) );
  AOI222XL U6123 ( .A0(n11221), .A1(n6226), .B0(result_r[10]), .B1(n9249), 
        .C0(N310), .C1(n9250), .Y(n9260) );
  MXI2X1 U6124 ( .A(n1705), .B(n10251), .S0(n8754), .Y(n4658) );
  CLKINVX1 U6125 ( .A(n9261), .Y(n4657) );
  AOI222XL U6126 ( .A0(n11216), .A1(n6227), .B0(result_r[11]), .B1(n9249), 
        .C0(N311), .C1(n9250), .Y(n9261) );
  MXI2X1 U6127 ( .A(n1703), .B(n10250), .S0(n8754), .Y(n4656) );
  CLKINVX1 U6128 ( .A(n9262), .Y(n4655) );
  AOI222XL U6129 ( .A0(n11222), .A1(n6228), .B0(result_r[12]), .B1(n9249), 
        .C0(N312), .C1(n9250), .Y(n9262) );
  MXI2X1 U6130 ( .A(n1701), .B(n10249), .S0(n8754), .Y(n4654) );
  CLKINVX1 U6131 ( .A(n9263), .Y(n4653) );
  AOI222XL U6132 ( .A0(n11222), .A1(n6229), .B0(result_r[13]), .B1(n9249), 
        .C0(N313), .C1(n9250), .Y(n9263) );
  MXI2X1 U6133 ( .A(n1699), .B(n10248), .S0(n8754), .Y(n4652) );
  CLKINVX1 U6134 ( .A(n9264), .Y(n4651) );
  AOI222XL U6135 ( .A0(n11222), .A1(n6230), .B0(result_r[14]), .B1(n9249), 
        .C0(N314), .C1(n9250), .Y(n9264) );
  MXI2X1 U6136 ( .A(n1697), .B(n10247), .S0(n8754), .Y(n4650) );
  CLKINVX1 U6137 ( .A(n9265), .Y(n4649) );
  AOI222XL U6138 ( .A0(n11215), .A1(n6231), .B0(result_r[15]), .B1(n9249), 
        .C0(N315), .C1(n9250), .Y(n9265) );
  MXI2X1 U6139 ( .A(n1695), .B(n10246), .S0(n8754), .Y(n4648) );
  CLKINVX1 U6140 ( .A(n9266), .Y(n4647) );
  AOI222XL U6141 ( .A0(n11223), .A1(n6232), .B0(result_r[16]), .B1(n9249), 
        .C0(N316), .C1(n9250), .Y(n9266) );
  MXI2X1 U6142 ( .A(n1693), .B(n10245), .S0(n8754), .Y(n4646) );
  CLKINVX1 U6143 ( .A(n9267), .Y(n4645) );
  AOI222XL U6144 ( .A0(n11223), .A1(n6233), .B0(result_r[17]), .B1(n9249), 
        .C0(N317), .C1(n9250), .Y(n9267) );
  MXI2X1 U6145 ( .A(n1691), .B(n10244), .S0(n8754), .Y(n4644) );
  CLKINVX1 U6146 ( .A(n9268), .Y(n4643) );
  AOI222XL U6147 ( .A0(n11223), .A1(n6234), .B0(result_r[18]), .B1(n9249), 
        .C0(N318), .C1(n9250), .Y(n9268) );
  MXI2X1 U6148 ( .A(n1689), .B(n10243), .S0(n8754), .Y(n4642) );
  CLKINVX1 U6149 ( .A(n9269), .Y(n4641) );
  AOI222XL U6150 ( .A0(n11216), .A1(n6235), .B0(result_r[19]), .B1(n9249), 
        .C0(N319), .C1(n9250), .Y(n9269) );
  MXI2X1 U6151 ( .A(n1687), .B(n10242), .S0(n8753), .Y(n4640) );
  CLKINVX1 U6152 ( .A(n9270), .Y(n4639) );
  AOI222XL U6153 ( .A0(n11224), .A1(n6236), .B0(result_r[20]), .B1(n9249), 
        .C0(N320), .C1(n9250), .Y(n9270) );
  MXI2X1 U6154 ( .A(n1685), .B(n10241), .S0(n8753), .Y(n4638) );
  CLKINVX1 U6155 ( .A(n9271), .Y(n4637) );
  AOI222XL U6156 ( .A0(n11224), .A1(n6237), .B0(result_r[21]), .B1(n9249), 
        .C0(N321), .C1(n9250), .Y(n9271) );
  MXI2X1 U6157 ( .A(n1683), .B(n10240), .S0(n8753), .Y(n4636) );
  CLKINVX1 U6158 ( .A(n9272), .Y(n4635) );
  AOI222XL U6159 ( .A0(n11224), .A1(n6238), .B0(result_r[22]), .B1(n9249), 
        .C0(N322), .C1(n9250), .Y(n9272) );
  MXI2X1 U6160 ( .A(n1681), .B(n10239), .S0(n8753), .Y(n4634) );
  CLKINVX1 U6161 ( .A(n9273), .Y(n4633) );
  AOI222XL U6162 ( .A0(n11215), .A1(n6239), .B0(result_r[23]), .B1(n9249), 
        .C0(N323), .C1(n9250), .Y(n9273) );
  MXI2X1 U6163 ( .A(n1679), .B(n10238), .S0(n8753), .Y(n4632) );
  CLKINVX1 U6164 ( .A(n9274), .Y(n4631) );
  AOI222XL U6165 ( .A0(n11221), .A1(n6240), .B0(result_r[24]), .B1(n9249), 
        .C0(N324), .C1(n9250), .Y(n9274) );
  MXI2X1 U6166 ( .A(n1677), .B(n10237), .S0(n8753), .Y(n4630) );
  CLKINVX1 U6167 ( .A(n9275), .Y(n4629) );
  AOI222XL U6168 ( .A0(n11221), .A1(n6241), .B0(result_r[25]), .B1(n9249), 
        .C0(N325), .C1(n9250), .Y(n9275) );
  MXI2X1 U6169 ( .A(n1675), .B(n10236), .S0(n8753), .Y(n4628) );
  CLKINVX1 U6170 ( .A(n9276), .Y(n4627) );
  AOI222XL U6171 ( .A0(n11221), .A1(n6242), .B0(result_r[26]), .B1(n9249), 
        .C0(N326), .C1(n9250), .Y(n9276) );
  MXI2X1 U6172 ( .A(n1673), .B(n10235), .S0(n8753), .Y(n4626) );
  CLKINVX1 U6173 ( .A(n9277), .Y(n4625) );
  AOI222XL U6174 ( .A0(n11216), .A1(n6243), .B0(result_r[27]), .B1(n9249), 
        .C0(N327), .C1(n9250), .Y(n9277) );
  MXI2X1 U6175 ( .A(n1671), .B(n10234), .S0(n8753), .Y(n4624) );
  CLKINVX1 U6176 ( .A(n9278), .Y(n4623) );
  AOI222XL U6177 ( .A0(n11222), .A1(n6244), .B0(result_r[28]), .B1(n9249), 
        .C0(N328), .C1(n9250), .Y(n9278) );
  MXI2X1 U6178 ( .A(n1669), .B(n10233), .S0(n8753), .Y(n4622) );
  CLKINVX1 U6179 ( .A(n9279), .Y(n4621) );
  AOI222XL U6180 ( .A0(n11222), .A1(n6245), .B0(result_r[29]), .B1(n9249), 
        .C0(N329), .C1(n9250), .Y(n9279) );
  MXI2X1 U6181 ( .A(n1667), .B(n10232), .S0(n8753), .Y(n4620) );
  CLKINVX1 U6182 ( .A(n9280), .Y(n4619) );
  AOI222XL U6183 ( .A0(n11222), .A1(n6246), .B0(result_r[30]), .B1(n9249), 
        .C0(N330), .C1(n9250), .Y(n9280) );
  MXI2X1 U6184 ( .A(n1665), .B(n10231), .S0(n8753), .Y(n4618) );
  CLKINVX1 U6185 ( .A(n9281), .Y(n4617) );
  AOI222XL U6186 ( .A0(n11215), .A1(n6247), .B0(result_r[31]), .B1(n9249), 
        .C0(N331), .C1(n9250), .Y(n9281) );
  MXI2X1 U6187 ( .A(n1663), .B(n10230), .S0(n8753), .Y(n4616) );
  CLKINVX1 U6188 ( .A(n9282), .Y(n4615) );
  AOI222XL U6189 ( .A0(n11223), .A1(n6248), .B0(result_i[0]), .B1(n9249), .C0(
        N332), .C1(n9250), .Y(n9282) );
  MXI2X1 U6190 ( .A(n1661), .B(n10229), .S0(n8752), .Y(n4614) );
  CLKINVX1 U6191 ( .A(n9283), .Y(n4613) );
  AOI222XL U6192 ( .A0(n11223), .A1(n6249), .B0(result_i[1]), .B1(n9249), .C0(
        N333), .C1(n9250), .Y(n9283) );
  MXI2X1 U6193 ( .A(n1659), .B(n10228), .S0(n8752), .Y(n4612) );
  CLKINVX1 U6194 ( .A(n9284), .Y(n4611) );
  AOI222XL U6195 ( .A0(n11223), .A1(n6250), .B0(result_i[2]), .B1(n9249), .C0(
        N334), .C1(n9250), .Y(n9284) );
  MXI2X1 U6196 ( .A(n1657), .B(n10227), .S0(n8752), .Y(n4610) );
  CLKINVX1 U6197 ( .A(n9285), .Y(n4609) );
  AOI222XL U6198 ( .A0(n11216), .A1(n6251), .B0(result_i[3]), .B1(n9249), .C0(
        N335), .C1(n9250), .Y(n9285) );
  MXI2X1 U6199 ( .A(n1655), .B(n10226), .S0(n8752), .Y(n4608) );
  CLKINVX1 U6200 ( .A(n9286), .Y(n4607) );
  AOI222XL U6201 ( .A0(n11224), .A1(n6252), .B0(result_i[4]), .B1(n9249), .C0(
        N336), .C1(n9250), .Y(n9286) );
  MXI2X1 U6202 ( .A(n1653), .B(n10225), .S0(n8752), .Y(n4606) );
  CLKINVX1 U6203 ( .A(n9287), .Y(n4605) );
  AOI222XL U6204 ( .A0(n11224), .A1(n6253), .B0(result_i[5]), .B1(n9249), .C0(
        N337), .C1(n9250), .Y(n9287) );
  MXI2X1 U6205 ( .A(n1651), .B(n10224), .S0(n8752), .Y(n4604) );
  CLKINVX1 U6206 ( .A(n9288), .Y(n4603) );
  AOI222XL U6207 ( .A0(n11224), .A1(n6254), .B0(result_i[6]), .B1(n9249), .C0(
        N338), .C1(n9250), .Y(n9288) );
  MXI2X1 U6208 ( .A(n1649), .B(n10223), .S0(n8752), .Y(n4602) );
  CLKINVX1 U6209 ( .A(n9289), .Y(n4601) );
  AOI222XL U6210 ( .A0(n11215), .A1(n6255), .B0(result_i[7]), .B1(n9249), .C0(
        N339), .C1(n9250), .Y(n9289) );
  MXI2X1 U6211 ( .A(n1647), .B(n10222), .S0(n8752), .Y(n4600) );
  CLKINVX1 U6212 ( .A(n9290), .Y(n4599) );
  AOI222XL U6213 ( .A0(n11221), .A1(n6256), .B0(result_i[8]), .B1(n9249), .C0(
        N340), .C1(n9250), .Y(n9290) );
  MXI2X1 U6214 ( .A(n1645), .B(n10221), .S0(n8752), .Y(n4598) );
  CLKINVX1 U6215 ( .A(n9291), .Y(n4597) );
  AOI222XL U6216 ( .A0(n11221), .A1(n6257), .B0(result_i[9]), .B1(n9249), .C0(
        N341), .C1(n9250), .Y(n9291) );
  MXI2X1 U6217 ( .A(n1643), .B(n10220), .S0(n8752), .Y(n4596) );
  CLKINVX1 U6218 ( .A(n9292), .Y(n4595) );
  AOI222XL U6219 ( .A0(n11221), .A1(n6258), .B0(result_i[10]), .B1(n9249), 
        .C0(N342), .C1(n9250), .Y(n9292) );
  MXI2X1 U6220 ( .A(n1641), .B(n10219), .S0(n8752), .Y(n4594) );
  CLKINVX1 U6221 ( .A(n9293), .Y(n4593) );
  AOI222XL U6222 ( .A0(n11216), .A1(n6259), .B0(result_i[11]), .B1(n9249), 
        .C0(N343), .C1(n9250), .Y(n9293) );
  MXI2X1 U6223 ( .A(n1639), .B(n10218), .S0(n8752), .Y(n4592) );
  CLKINVX1 U6224 ( .A(n9294), .Y(n4591) );
  AOI222XL U6225 ( .A0(n11222), .A1(n6260), .B0(result_i[12]), .B1(n9249), 
        .C0(N344), .C1(n9250), .Y(n9294) );
  MXI2X1 U6226 ( .A(n1637), .B(n10217), .S0(n8752), .Y(n4590) );
  CLKINVX1 U6227 ( .A(n9295), .Y(n4589) );
  AOI222XL U6228 ( .A0(n11222), .A1(n6261), .B0(result_i[13]), .B1(n9249), 
        .C0(N345), .C1(n9250), .Y(n9295) );
  MXI2X1 U6229 ( .A(n1635), .B(n10216), .S0(n8751), .Y(n4588) );
  CLKINVX1 U6230 ( .A(n9296), .Y(n4587) );
  AOI222XL U6231 ( .A0(n11222), .A1(n6262), .B0(result_i[14]), .B1(n9249), 
        .C0(N346), .C1(n9250), .Y(n9296) );
  MXI2X1 U6232 ( .A(n1633), .B(n10215), .S0(n8751), .Y(n4586) );
  CLKINVX1 U6233 ( .A(n9297), .Y(n4585) );
  AOI222XL U6234 ( .A0(n11215), .A1(n6263), .B0(result_i[15]), .B1(n9249), 
        .C0(N347), .C1(n9250), .Y(n9297) );
  MXI2X1 U6235 ( .A(n1631), .B(n10214), .S0(n8751), .Y(n4584) );
  CLKINVX1 U6236 ( .A(n9298), .Y(n4583) );
  AOI222XL U6237 ( .A0(n11223), .A1(n6264), .B0(result_i[16]), .B1(n9249), 
        .C0(N348), .C1(n9250), .Y(n9298) );
  MXI2X1 U6238 ( .A(n1629), .B(n10213), .S0(n8751), .Y(n4582) );
  CLKINVX1 U6239 ( .A(n9299), .Y(n4581) );
  AOI222XL U6240 ( .A0(n11223), .A1(n6265), .B0(result_i[17]), .B1(n9249), 
        .C0(N349), .C1(n9250), .Y(n9299) );
  MXI2X1 U6241 ( .A(n1627), .B(n10212), .S0(n8751), .Y(n4580) );
  CLKINVX1 U6242 ( .A(n9300), .Y(n4579) );
  AOI222XL U6243 ( .A0(n11223), .A1(n6266), .B0(result_i[18]), .B1(n9249), 
        .C0(N350), .C1(n9250), .Y(n9300) );
  MXI2X1 U6244 ( .A(n1625), .B(n10211), .S0(n8751), .Y(n4578) );
  CLKINVX1 U6245 ( .A(n9301), .Y(n4577) );
  AOI222XL U6246 ( .A0(n11216), .A1(n6267), .B0(result_i[19]), .B1(n9249), 
        .C0(N351), .C1(n9250), .Y(n9301) );
  MXI2X1 U6247 ( .A(n1623), .B(n10210), .S0(n8751), .Y(n4576) );
  CLKINVX1 U6248 ( .A(n9302), .Y(n4575) );
  AOI222XL U6249 ( .A0(n11224), .A1(n6268), .B0(result_i[20]), .B1(n9249), 
        .C0(N352), .C1(n9250), .Y(n9302) );
  MXI2X1 U6250 ( .A(n1621), .B(n10209), .S0(n8751), .Y(n4574) );
  CLKINVX1 U6251 ( .A(n9303), .Y(n4573) );
  AOI222XL U6252 ( .A0(n11224), .A1(n6269), .B0(result_i[21]), .B1(n9249), 
        .C0(N353), .C1(n9250), .Y(n9303) );
  MXI2X1 U6253 ( .A(n1619), .B(n10208), .S0(n8751), .Y(n4572) );
  CLKINVX1 U6254 ( .A(n9304), .Y(n4571) );
  AOI222XL U6255 ( .A0(n11224), .A1(n6270), .B0(result_i[22]), .B1(n9249), 
        .C0(N354), .C1(n9250), .Y(n9304) );
  MXI2X1 U6256 ( .A(n1617), .B(n10207), .S0(n8751), .Y(n4570) );
  CLKINVX1 U6257 ( .A(n9305), .Y(n4569) );
  AOI222XL U6258 ( .A0(n11215), .A1(n6271), .B0(result_i[23]), .B1(n9249), 
        .C0(N355), .C1(n9250), .Y(n9305) );
  MXI2X1 U6259 ( .A(n1615), .B(n10206), .S0(n8751), .Y(n4568) );
  CLKINVX1 U6260 ( .A(n9306), .Y(n4567) );
  AOI222XL U6261 ( .A0(n11221), .A1(n6272), .B0(result_i[24]), .B1(n9249), 
        .C0(N356), .C1(n9250), .Y(n9306) );
  MXI2X1 U6262 ( .A(n1613), .B(n10205), .S0(n8751), .Y(n4566) );
  CLKINVX1 U6263 ( .A(n9307), .Y(n4565) );
  AOI222XL U6264 ( .A0(n11221), .A1(n6273), .B0(result_i[25]), .B1(n9249), 
        .C0(N357), .C1(n9250), .Y(n9307) );
  MXI2X1 U6265 ( .A(n1611), .B(n10204), .S0(n8751), .Y(n4564) );
  CLKINVX1 U6266 ( .A(n9308), .Y(n4563) );
  AOI222XL U6267 ( .A0(n11221), .A1(n6274), .B0(result_i[26]), .B1(n9249), 
        .C0(N358), .C1(n9250), .Y(n9308) );
  MXI2X1 U6268 ( .A(n1609), .B(n10203), .S0(n8750), .Y(n4562) );
  CLKINVX1 U6269 ( .A(n9309), .Y(n4561) );
  AOI222XL U6270 ( .A0(n11216), .A1(n6275), .B0(result_i[27]), .B1(n9249), 
        .C0(N359), .C1(n9250), .Y(n9309) );
  MXI2X1 U6271 ( .A(n1607), .B(n10202), .S0(n8750), .Y(n4560) );
  CLKINVX1 U6272 ( .A(n9310), .Y(n4559) );
  AOI222XL U6273 ( .A0(n11222), .A1(n6276), .B0(result_i[28]), .B1(n9249), 
        .C0(N360), .C1(n9250), .Y(n9310) );
  MXI2X1 U6274 ( .A(n1605), .B(n10201), .S0(n8750), .Y(n4558) );
  CLKINVX1 U6275 ( .A(n9311), .Y(n4557) );
  AOI222XL U6276 ( .A0(n11222), .A1(n6277), .B0(result_i[29]), .B1(n9249), 
        .C0(N361), .C1(n9250), .Y(n9311) );
  MXI2X1 U6277 ( .A(n1603), .B(n10200), .S0(n8750), .Y(n4556) );
  CLKINVX1 U6278 ( .A(n9312), .Y(n4555) );
  AOI222XL U6279 ( .A0(n11222), .A1(n6278), .B0(result_i[30]), .B1(n9249), 
        .C0(N362), .C1(n9250), .Y(n9312) );
  MXI2X1 U6280 ( .A(n1601), .B(n10199), .S0(n8750), .Y(n4554) );
  CLKINVX1 U6281 ( .A(n9313), .Y(n4553) );
  AOI222XL U6282 ( .A0(n11215), .A1(n6279), .B0(result_i[31]), .B1(n9249), 
        .C0(N363), .C1(n9250), .Y(n9313) );
  MXI2X1 U6283 ( .A(n1599), .B(n10198), .S0(n8750), .Y(n4552) );
  OAI222XL U6284 ( .A0(n8756), .A1(n6175), .B0(n9314), .B1(n9315), .C0(n9316), 
        .C1(n9317), .Y(n4551) );
  CLKINVX1 U6285 ( .A(N400), .Y(n9314) );
  OAI222XL U6286 ( .A0(n8757), .A1(n6174), .B0(n9318), .B1(n9315), .C0(n9319), 
        .C1(n9317), .Y(n4550) );
  CLKINVX1 U6287 ( .A(N401), .Y(n9318) );
  OAI222XL U6288 ( .A0(n8756), .A1(n6173), .B0(n9320), .B1(n9315), .C0(n9321), 
        .C1(n9317), .Y(n4549) );
  CLKINVX1 U6289 ( .A(N402), .Y(n9320) );
  OAI222XL U6290 ( .A0(n8757), .A1(n6172), .B0(n9322), .B1(n9315), .C0(n9323), 
        .C1(n9317), .Y(n4548) );
  CLKINVX1 U6291 ( .A(N403), .Y(n9322) );
  OAI222XL U6292 ( .A0(n8756), .A1(n6171), .B0(n9324), .B1(n9315), .C0(n9325), 
        .C1(n9317), .Y(n4547) );
  CLKINVX1 U6293 ( .A(N404), .Y(n9324) );
  OAI222XL U6294 ( .A0(n8756), .A1(n6170), .B0(n9326), .B1(n9315), .C0(n9327), 
        .C1(n9317), .Y(n4546) );
  CLKINVX1 U6295 ( .A(N405), .Y(n9326) );
  OAI222XL U6296 ( .A0(n8756), .A1(n6169), .B0(n9328), .B1(n9315), .C0(n9329), 
        .C1(n9317), .Y(n4545) );
  CLKINVX1 U6297 ( .A(N406), .Y(n9328) );
  OAI222XL U6298 ( .A0(n8757), .A1(n6168), .B0(n9330), .B1(n9315), .C0(n9331), 
        .C1(n9317), .Y(n4544) );
  CLKINVX1 U6299 ( .A(N407), .Y(n9330) );
  OAI222XL U6300 ( .A0(n8756), .A1(n6167), .B0(n9332), .B1(n9315), .C0(n9333), 
        .C1(n9317), .Y(n4543) );
  CLKINVX1 U6301 ( .A(N408), .Y(n9332) );
  OAI222XL U6302 ( .A0(n8757), .A1(n6166), .B0(n9334), .B1(n9315), .C0(n9335), 
        .C1(n9317), .Y(n4542) );
  CLKINVX1 U6303 ( .A(N409), .Y(n9334) );
  OAI222XL U6304 ( .A0(n8756), .A1(n6165), .B0(n9336), .B1(n9315), .C0(n9337), 
        .C1(n9317), .Y(n4541) );
  CLKINVX1 U6305 ( .A(N410), .Y(n9336) );
  OAI222XL U6306 ( .A0(n8757), .A1(n6164), .B0(n9338), .B1(n9315), .C0(n9339), 
        .C1(n9317), .Y(n4540) );
  CLKINVX1 U6307 ( .A(N411), .Y(n9338) );
  OAI222XL U6308 ( .A0(n8756), .A1(n6163), .B0(n9340), .B1(n9315), .C0(n9341), 
        .C1(n9317), .Y(n4539) );
  CLKINVX1 U6309 ( .A(N412), .Y(n9340) );
  OAI222XL U6310 ( .A0(n8757), .A1(n6162), .B0(n9342), .B1(n9315), .C0(n9343), 
        .C1(n9317), .Y(n4538) );
  CLKINVX1 U6311 ( .A(N413), .Y(n9342) );
  OAI222XL U6312 ( .A0(n8756), .A1(n6161), .B0(n9344), .B1(n9315), .C0(n9345), 
        .C1(n9317), .Y(n4537) );
  CLKINVX1 U6313 ( .A(N414), .Y(n9344) );
  OAI222XL U6314 ( .A0(n8756), .A1(n6160), .B0(n9346), .B1(n9315), .C0(n9347), 
        .C1(n9317), .Y(n4536) );
  CLKINVX1 U6315 ( .A(N415), .Y(n9346) );
  OAI222XL U6316 ( .A0(n8756), .A1(n6159), .B0(n9348), .B1(n9315), .C0(n9349), 
        .C1(n9317), .Y(n4535) );
  CLKINVX1 U6317 ( .A(N416), .Y(n9348) );
  OAI222XL U6318 ( .A0(n8756), .A1(n6158), .B0(n9350), .B1(n9315), .C0(n9351), 
        .C1(n9317), .Y(n4534) );
  CLKINVX1 U6319 ( .A(N417), .Y(n9350) );
  OAI222XL U6320 ( .A0(n8756), .A1(n6157), .B0(n9352), .B1(n9315), .C0(n9353), 
        .C1(n9317), .Y(n4533) );
  CLKINVX1 U6321 ( .A(N418), .Y(n9352) );
  OAI222XL U6322 ( .A0(n8757), .A1(n6156), .B0(n9354), .B1(n9315), .C0(n9355), 
        .C1(n9317), .Y(n4532) );
  CLKINVX1 U6323 ( .A(N419), .Y(n9354) );
  OAI222XL U6324 ( .A0(n8756), .A1(n6155), .B0(n9356), .B1(n9315), .C0(n9357), 
        .C1(n9317), .Y(n4531) );
  CLKINVX1 U6325 ( .A(N420), .Y(n9356) );
  OAI222XL U6326 ( .A0(n8757), .A1(n6154), .B0(n9358), .B1(n9315), .C0(n9359), 
        .C1(n9317), .Y(n4530) );
  CLKINVX1 U6327 ( .A(N421), .Y(n9358) );
  OAI222XL U6328 ( .A0(n8756), .A1(n6153), .B0(n9360), .B1(n9315), .C0(n9361), 
        .C1(n9317), .Y(n4529) );
  CLKINVX1 U6329 ( .A(N422), .Y(n9360) );
  OAI222XL U6330 ( .A0(n8757), .A1(n6152), .B0(n9362), .B1(n9315), .C0(n9363), 
        .C1(n9317), .Y(n4528) );
  CLKINVX1 U6331 ( .A(N423), .Y(n9362) );
  OAI222XL U6332 ( .A0(n8756), .A1(n6151), .B0(n9364), .B1(n9315), .C0(n9365), 
        .C1(n9317), .Y(n4527) );
  CLKINVX1 U6333 ( .A(N424), .Y(n9364) );
  OAI222XL U6334 ( .A0(n8756), .A1(n6150), .B0(n9366), .B1(n9315), .C0(n9367), 
        .C1(n9317), .Y(n4526) );
  CLKINVX1 U6335 ( .A(N425), .Y(n9366) );
  OAI222XL U6336 ( .A0(n8756), .A1(n6149), .B0(n9368), .B1(n9315), .C0(n9369), 
        .C1(n9317), .Y(n4525) );
  CLKINVX1 U6337 ( .A(N426), .Y(n9368) );
  OAI222XL U6338 ( .A0(n8757), .A1(n6148), .B0(n9370), .B1(n9315), .C0(n9371), 
        .C1(n9317), .Y(n4524) );
  CLKINVX1 U6339 ( .A(N427), .Y(n9370) );
  OAI222XL U6340 ( .A0(n8757), .A1(n6147), .B0(n9372), .B1(n9315), .C0(n9373), 
        .C1(n9317), .Y(n4523) );
  CLKINVX1 U6341 ( .A(N428), .Y(n9372) );
  OAI222XL U6342 ( .A0(n8757), .A1(n6146), .B0(n9374), .B1(n9315), .C0(n9375), 
        .C1(n9317), .Y(n4522) );
  CLKINVX1 U6343 ( .A(N429), .Y(n9374) );
  OAI222XL U6344 ( .A0(n8756), .A1(n6145), .B0(n9376), .B1(n9315), .C0(n9377), 
        .C1(n9317), .Y(n4521) );
  CLKINVX1 U6345 ( .A(N430), .Y(n9376) );
  OAI222XL U6346 ( .A0(n8756), .A1(n6144), .B0(n9378), .B1(n9315), .C0(n9379), 
        .C1(n9317), .Y(n4520) );
  CLKINVX1 U6347 ( .A(N431), .Y(n9378) );
  CLKINVX1 U6348 ( .A(n9382), .Y(n4519) );
  AOI221XL U6349 ( .A0(n9383), .A1(N448), .B0(n9384), .B1(N368), .C0(n9385), 
        .Y(n9382) );
  OAI22XL U6350 ( .A0(n9386), .A1(n9317), .B0(n8758), .B1(n6127), .Y(n9385) );
  CLKINVX1 U6351 ( .A(n9387), .Y(n4518) );
  AOI221XL U6352 ( .A0(n9383), .A1(N463), .B0(n9384), .B1(N383), .C0(n9388), 
        .Y(n9387) );
  OAI22XL U6353 ( .A0(n9389), .A1(n9317), .B0(n8758), .B1(n6112), .Y(n9388) );
  OAI221XL U6354 ( .A0(n9317), .A1(n9390), .B0(n6143), .B1(n8757), .C0(n9391), 
        .Y(n4517) );
  AOI22X1 U6355 ( .A0(N432), .A1(n9383), .B0(N528), .B1(n9384), .Y(n9391) );
  OAI221XL U6356 ( .A0(n9317), .A1(n9392), .B0(n6142), .B1(n8758), .C0(n9393), 
        .Y(n4516) );
  OAI221XL U6357 ( .A0(n9317), .A1(n9394), .B0(n6141), .B1(n8758), .C0(n9395), 
        .Y(n4515) );
  OAI221XL U6358 ( .A0(n9317), .A1(n9396), .B0(n6140), .B1(n8758), .C0(n9397), 
        .Y(n4514) );
  OAI221XL U6359 ( .A0(n9317), .A1(n9398), .B0(n6139), .B1(n8757), .C0(n9399), 
        .Y(n4513) );
  OAI221XL U6360 ( .A0(n9317), .A1(n9400), .B0(n6138), .B1(n8757), .C0(n9401), 
        .Y(n4512) );
  OAI221XL U6361 ( .A0(n9317), .A1(n9402), .B0(n6137), .B1(n8757), .C0(n9403), 
        .Y(n4511) );
  OAI221XL U6362 ( .A0(n9317), .A1(n9404), .B0(n6136), .B1(n8757), .C0(n9405), 
        .Y(n4510) );
  OAI221XL U6363 ( .A0(n9317), .A1(n9406), .B0(n6135), .B1(n8758), .C0(n9407), 
        .Y(n4509) );
  OAI221XL U6364 ( .A0(n9317), .A1(n9408), .B0(n6134), .B1(n8757), .C0(n9409), 
        .Y(n4508) );
  OAI221XL U6365 ( .A0(n9317), .A1(n9410), .B0(n6133), .B1(n8757), .C0(n9411), 
        .Y(n4507) );
  OAI221XL U6366 ( .A0(n9317), .A1(n9412), .B0(n6132), .B1(n8757), .C0(n9413), 
        .Y(n4506) );
  OAI221XL U6367 ( .A0(n9317), .A1(n9414), .B0(n6131), .B1(n8757), .C0(n9415), 
        .Y(n4505) );
  OAI221XL U6368 ( .A0(n9317), .A1(n9416), .B0(n6130), .B1(n8757), .C0(n9417), 
        .Y(n4504) );
  OAI221XL U6369 ( .A0(n9317), .A1(n9418), .B0(n6129), .B1(n8757), .C0(n9419), 
        .Y(n4503) );
  OAI221XL U6370 ( .A0(n9317), .A1(n9420), .B0(n6128), .B1(n8757), .C0(n9421), 
        .Y(n4502) );
  AOI22X1 U6371 ( .A0(N447), .A1(n9383), .B0(N543), .B1(n9384), .Y(n9421) );
  CLKINVX1 U6372 ( .A(n9422), .Y(n4501) );
  AOI221XL U6373 ( .A0(n9383), .A1(N449), .B0(n9384), .B1(N369), .C0(n9423), 
        .Y(n9422) );
  OAI22XL U6374 ( .A0(n9424), .A1(n9317), .B0(n8758), .B1(n6126), .Y(n9423) );
  CLKINVX1 U6375 ( .A(n9425), .Y(n4500) );
  AOI221XL U6376 ( .A0(n9383), .A1(N450), .B0(n9384), .B1(N370), .C0(n9426), 
        .Y(n9425) );
  OAI22XL U6377 ( .A0(n9427), .A1(n9317), .B0(n8758), .B1(n6125), .Y(n9426) );
  CLKINVX1 U6378 ( .A(n9428), .Y(n4499) );
  AOI221XL U6379 ( .A0(n9383), .A1(N451), .B0(n9384), .B1(N371), .C0(n9429), 
        .Y(n9428) );
  OAI22XL U6380 ( .A0(n9430), .A1(n9317), .B0(n8758), .B1(n6124), .Y(n9429) );
  CLKINVX1 U6381 ( .A(n9431), .Y(n4498) );
  AOI221XL U6382 ( .A0(n9383), .A1(N452), .B0(n9384), .B1(N372), .C0(n9432), 
        .Y(n9431) );
  OAI22XL U6383 ( .A0(n9433), .A1(n9317), .B0(n8758), .B1(n6123), .Y(n9432) );
  CLKINVX1 U6384 ( .A(n9434), .Y(n4497) );
  AOI221XL U6385 ( .A0(n9383), .A1(N453), .B0(n9384), .B1(N373), .C0(n9435), 
        .Y(n9434) );
  OAI22XL U6386 ( .A0(n9436), .A1(n9317), .B0(n8758), .B1(n6122), .Y(n9435) );
  CLKINVX1 U6387 ( .A(n9437), .Y(n4496) );
  AOI221XL U6388 ( .A0(n9383), .A1(N454), .B0(n9384), .B1(N374), .C0(n9438), 
        .Y(n9437) );
  OAI22XL U6389 ( .A0(n9439), .A1(n9317), .B0(n8758), .B1(n6121), .Y(n9438) );
  CLKINVX1 U6390 ( .A(n9440), .Y(n4495) );
  AOI221XL U6391 ( .A0(n9383), .A1(N455), .B0(n9384), .B1(N375), .C0(n9441), 
        .Y(n9440) );
  OAI22XL U6392 ( .A0(n9442), .A1(n9317), .B0(n8758), .B1(n6120), .Y(n9441) );
  CLKINVX1 U6393 ( .A(n9443), .Y(n4494) );
  AOI221XL U6394 ( .A0(n9383), .A1(N456), .B0(n9384), .B1(N376), .C0(n9444), 
        .Y(n9443) );
  OAI22XL U6395 ( .A0(n9445), .A1(n9317), .B0(n8758), .B1(n6119), .Y(n9444) );
  CLKINVX1 U6396 ( .A(n9446), .Y(n4493) );
  AOI221XL U6397 ( .A0(n9383), .A1(N457), .B0(n9384), .B1(N377), .C0(n9447), 
        .Y(n9446) );
  OAI22XL U6398 ( .A0(n9448), .A1(n9317), .B0(n8758), .B1(n6118), .Y(n9447) );
  CLKINVX1 U6399 ( .A(n9449), .Y(n4492) );
  AOI221XL U6400 ( .A0(n9383), .A1(N458), .B0(n9384), .B1(N378), .C0(n9450), 
        .Y(n9449) );
  OAI22XL U6401 ( .A0(n9451), .A1(n9317), .B0(n8758), .B1(n6117), .Y(n9450) );
  CLKINVX1 U6402 ( .A(n9452), .Y(n4491) );
  AOI221XL U6403 ( .A0(n9383), .A1(N459), .B0(n9384), .B1(N379), .C0(n9453), 
        .Y(n9452) );
  OAI22XL U6404 ( .A0(n9454), .A1(n9317), .B0(n8758), .B1(n6116), .Y(n9453) );
  CLKINVX1 U6405 ( .A(n9455), .Y(n4490) );
  AOI221XL U6406 ( .A0(n9383), .A1(N460), .B0(n9384), .B1(N380), .C0(n9456), 
        .Y(n9455) );
  OAI22XL U6407 ( .A0(n9457), .A1(n9317), .B0(n8758), .B1(n6115), .Y(n9456) );
  CLKINVX1 U6408 ( .A(n9458), .Y(n4489) );
  AOI221XL U6409 ( .A0(n9383), .A1(N461), .B0(n9384), .B1(N381), .C0(n9459), 
        .Y(n9458) );
  OAI22XL U6410 ( .A0(n9460), .A1(n9317), .B0(n8758), .B1(n6114), .Y(n9459) );
  CLKINVX1 U6411 ( .A(n9461), .Y(n4488) );
  AOI221XL U6412 ( .A0(n9383), .A1(N462), .B0(n9384), .B1(N382), .C0(n9462), 
        .Y(n9461) );
  OAI22XL U6413 ( .A0(n9463), .A1(n9317), .B0(n8758), .B1(n6113), .Y(n9462) );
  NOR2X1 U6414 ( .A(n8792), .B(n11216), .Y(n9384) );
  NOR2X1 U6415 ( .A(n8781), .B(n11221), .Y(n9383) );
  OAI221XL U6416 ( .A0(n6144), .A1(n9466), .B0(n10197), .B1(n8838), .C0(n9467), 
        .Y(n4487) );
  OAI221XL U6417 ( .A0(n6145), .A1(n9466), .B0(n10196), .B1(n8838), .C0(n9470), 
        .Y(n4486) );
  OAI221XL U6418 ( .A0(n6146), .A1(n9466), .B0(n10195), .B1(n8837), .C0(n9471), 
        .Y(n4485) );
  OAI221XL U6419 ( .A0(n6147), .A1(n9466), .B0(n10194), .B1(n8828), .C0(n9472), 
        .Y(n4484) );
  OAI221XL U6420 ( .A0(n6148), .A1(n9466), .B0(n10193), .B1(n8829), .C0(n9473), 
        .Y(n4483) );
  OAI221XL U6421 ( .A0(n6149), .A1(n9466), .B0(n10192), .B1(n8830), .C0(n9474), 
        .Y(n4482) );
  OAI221XL U6422 ( .A0(n6150), .A1(n9466), .B0(n10191), .B1(n8831), .C0(n9475), 
        .Y(n4481) );
  OAI221XL U6423 ( .A0(n6151), .A1(n9466), .B0(n10190), .B1(n8832), .C0(n9476), 
        .Y(n4480) );
  OAI221XL U6424 ( .A0(n6152), .A1(n9466), .B0(n10189), .B1(n8838), .C0(n9477), 
        .Y(n4479) );
  OAI221XL U6425 ( .A0(n6153), .A1(n9466), .B0(n10188), .B1(n8838), .C0(n9478), 
        .Y(n4478) );
  OAI221XL U6426 ( .A0(n6154), .A1(n9466), .B0(n10187), .B1(n8838), .C0(n9479), 
        .Y(n4477) );
  OAI221XL U6427 ( .A0(n6155), .A1(n9466), .B0(n10186), .B1(n8838), .C0(n9480), 
        .Y(n4476) );
  OAI221XL U6428 ( .A0(n6156), .A1(n9466), .B0(n10185), .B1(n8838), .C0(n9481), 
        .Y(n4475) );
  OAI221XL U6429 ( .A0(n6157), .A1(n9466), .B0(n10184), .B1(n8838), .C0(n9482), 
        .Y(n4474) );
  OAI221XL U6430 ( .A0(n6158), .A1(n9466), .B0(n10183), .B1(n8838), .C0(n9483), 
        .Y(n4473) );
  OAI221XL U6431 ( .A0(n6159), .A1(n9466), .B0(n10182), .B1(n8838), .C0(n9484), 
        .Y(n4472) );
  OAI221XL U6432 ( .A0(n6112), .A1(n9466), .B0(n10181), .B1(n8838), .C0(n9485), 
        .Y(n4471) );
  OAI221XL U6433 ( .A0(n6113), .A1(n9466), .B0(n10180), .B1(n8838), .C0(n9486), 
        .Y(n4470) );
  OAI221XL U6434 ( .A0(n6114), .A1(n9466), .B0(n10179), .B1(n8838), .C0(n9487), 
        .Y(n4469) );
  OAI221XL U6435 ( .A0(n6115), .A1(n9466), .B0(n10178), .B1(n8838), .C0(n9488), 
        .Y(n4468) );
  OAI221XL U6436 ( .A0(n6116), .A1(n9466), .B0(n10177), .B1(n8838), .C0(n9489), 
        .Y(n4467) );
  OAI221XL U6437 ( .A0(n6117), .A1(n9466), .B0(n10176), .B1(n8838), .C0(n9490), 
        .Y(n4466) );
  OAI221XL U6438 ( .A0(n6118), .A1(n9466), .B0(n10175), .B1(n8838), .C0(n9491), 
        .Y(n4465) );
  OAI221XL U6439 ( .A0(n6119), .A1(n9466), .B0(n10174), .B1(n8838), .C0(n9492), 
        .Y(n4464) );
  OAI221XL U6440 ( .A0(n6120), .A1(n9466), .B0(n10173), .B1(n8838), .C0(n9493), 
        .Y(n4463) );
  OAI221XL U6441 ( .A0(n6121), .A1(n9466), .B0(n10172), .B1(n8838), .C0(n9494), 
        .Y(n4462) );
  OAI221XL U6442 ( .A0(n6122), .A1(n9466), .B0(n10171), .B1(n8838), .C0(n9495), 
        .Y(n4461) );
  OAI221XL U6443 ( .A0(n6123), .A1(n9466), .B0(n10170), .B1(n8838), .C0(n9496), 
        .Y(n4460) );
  OAI221XL U6444 ( .A0(n6124), .A1(n9466), .B0(n10169), .B1(n8838), .C0(n9497), 
        .Y(n4459) );
  AOI22X1 U6445 ( .A0(n9468), .A1(N451), .B0(N387), .B1(n9469), .Y(n9497) );
  OAI221XL U6446 ( .A0(n6125), .A1(n9466), .B0(n10168), .B1(n8838), .C0(n9498), 
        .Y(n4458) );
  AOI22X1 U6447 ( .A0(n9468), .A1(N450), .B0(N386), .B1(n9469), .Y(n9498) );
  OAI221XL U6448 ( .A0(n6126), .A1(n9466), .B0(n10167), .B1(n8838), .C0(n9499), 
        .Y(n4457) );
  AOI22X1 U6449 ( .A0(n9468), .A1(N449), .B0(N385), .B1(n9469), .Y(n9499) );
  OAI221XL U6450 ( .A0(n6127), .A1(n9466), .B0(n10166), .B1(n8838), .C0(n9500), 
        .Y(n4456) );
  AOI22X1 U6451 ( .A0(n9468), .A1(N448), .B0(N384), .B1(n9469), .Y(n9500) );
  NOR2X1 U6452 ( .A(n8781), .B(n8840), .Y(n9469) );
  NOR2X1 U6453 ( .A(n8792), .B(n8839), .Y(n9468) );
  NAND3X1 U6454 ( .A(n8792), .B(n8781), .C(n8837), .Y(n9466) );
  MXI2X1 U6455 ( .A(n10165), .B(n10197), .S0(n8837), .Y(n4455) );
  MXI2X1 U6456 ( .A(n10164), .B(n10196), .S0(n8837), .Y(n4454) );
  MXI2X1 U6457 ( .A(n10163), .B(n10195), .S0(n8837), .Y(n4453) );
  MXI2X1 U6458 ( .A(n10162), .B(n10194), .S0(n8837), .Y(n4452) );
  MXI2X1 U6459 ( .A(n10161), .B(n10193), .S0(n8837), .Y(n4451) );
  MXI2X1 U6460 ( .A(n10160), .B(n10192), .S0(n8837), .Y(n4450) );
  MXI2X1 U6461 ( .A(n10159), .B(n10191), .S0(n8837), .Y(n4449) );
  MXI2X1 U6462 ( .A(n10158), .B(n10190), .S0(n8837), .Y(n4448) );
  MXI2X1 U6463 ( .A(n10157), .B(n10189), .S0(n8837), .Y(n4447) );
  MXI2X1 U6464 ( .A(n10156), .B(n10188), .S0(n8837), .Y(n4446) );
  MXI2X1 U6465 ( .A(n10155), .B(n10187), .S0(n8837), .Y(n4445) );
  MXI2X1 U6466 ( .A(n10154), .B(n10186), .S0(n8837), .Y(n4444) );
  MXI2X1 U6467 ( .A(n10153), .B(n10185), .S0(n8836), .Y(n4443) );
  MXI2X1 U6468 ( .A(n10152), .B(n10184), .S0(n8836), .Y(n4442) );
  MXI2X1 U6469 ( .A(n10151), .B(n10183), .S0(n8836), .Y(n4441) );
  MXI2X1 U6470 ( .A(n10150), .B(n10182), .S0(n8836), .Y(n4440) );
  MXI2X1 U6471 ( .A(n10149), .B(n10181), .S0(n8836), .Y(n4439) );
  MXI2X1 U6472 ( .A(n10148), .B(n10180), .S0(n8836), .Y(n4438) );
  MXI2X1 U6473 ( .A(n10147), .B(n10179), .S0(n8836), .Y(n4437) );
  MXI2X1 U6474 ( .A(n10146), .B(n10178), .S0(n8836), .Y(n4436) );
  MXI2X1 U6475 ( .A(n10145), .B(n10177), .S0(n8836), .Y(n4435) );
  MXI2X1 U6476 ( .A(n10144), .B(n10176), .S0(n8836), .Y(n4434) );
  MXI2X1 U6477 ( .A(n10143), .B(n10175), .S0(n8836), .Y(n4433) );
  MXI2X1 U6478 ( .A(n10142), .B(n10174), .S0(n8836), .Y(n4432) );
  MXI2X1 U6479 ( .A(n10141), .B(n10173), .S0(n8836), .Y(n4431) );
  MXI2X1 U6480 ( .A(n10140), .B(n10172), .S0(n8835), .Y(n4430) );
  MXI2X1 U6481 ( .A(n10139), .B(n10171), .S0(n8835), .Y(n4429) );
  MXI2X1 U6482 ( .A(n10138), .B(n10170), .S0(n8835), .Y(n4428) );
  MXI2X1 U6483 ( .A(n10137), .B(n10169), .S0(n8835), .Y(n4427) );
  MXI2X1 U6484 ( .A(n10136), .B(n10168), .S0(n8835), .Y(n4426) );
  MXI2X1 U6485 ( .A(n10135), .B(n10167), .S0(n8835), .Y(n4425) );
  MXI2X1 U6486 ( .A(n10134), .B(n10166), .S0(n8835), .Y(n4424) );
  MXI2X1 U6487 ( .A(n10133), .B(n10165), .S0(n8835), .Y(n4423) );
  MXI2X1 U6488 ( .A(n10132), .B(n10164), .S0(n8835), .Y(n4422) );
  MXI2X1 U6489 ( .A(n10131), .B(n10163), .S0(n8835), .Y(n4421) );
  MXI2X1 U6490 ( .A(n10130), .B(n10162), .S0(n8835), .Y(n4420) );
  MXI2X1 U6491 ( .A(n10129), .B(n10161), .S0(n8835), .Y(n4419) );
  MXI2X1 U6492 ( .A(n10128), .B(n10160), .S0(n8835), .Y(n4418) );
  MXI2X1 U6493 ( .A(n10127), .B(n10159), .S0(n8834), .Y(n4417) );
  MXI2X1 U6494 ( .A(n10126), .B(n10158), .S0(n8834), .Y(n4416) );
  MXI2X1 U6495 ( .A(n10125), .B(n10157), .S0(n8834), .Y(n4415) );
  MXI2X1 U6496 ( .A(n10124), .B(n10156), .S0(n8834), .Y(n4414) );
  MXI2X1 U6497 ( .A(n10123), .B(n10155), .S0(n8834), .Y(n4413) );
  MXI2X1 U6498 ( .A(n10122), .B(n10154), .S0(n8834), .Y(n4412) );
  MXI2X1 U6499 ( .A(n10121), .B(n10153), .S0(n8834), .Y(n4411) );
  MXI2X1 U6500 ( .A(n10120), .B(n10152), .S0(n8834), .Y(n4410) );
  MXI2X1 U6501 ( .A(n10119), .B(n10151), .S0(n8834), .Y(n4409) );
  MXI2X1 U6502 ( .A(n10118), .B(n10150), .S0(n8834), .Y(n4408) );
  MXI2X1 U6503 ( .A(n10117), .B(n10149), .S0(n8834), .Y(n4407) );
  MXI2X1 U6504 ( .A(n10116), .B(n10148), .S0(n8834), .Y(n4406) );
  MXI2X1 U6505 ( .A(n10115), .B(n10147), .S0(n8834), .Y(n4405) );
  MXI2X1 U6506 ( .A(n10114), .B(n10146), .S0(n8833), .Y(n4404) );
  MXI2X1 U6507 ( .A(n10113), .B(n10145), .S0(n8833), .Y(n4403) );
  MXI2X1 U6508 ( .A(n10112), .B(n10144), .S0(n8833), .Y(n4402) );
  MXI2X1 U6509 ( .A(n10111), .B(n10143), .S0(n8833), .Y(n4401) );
  MXI2X1 U6510 ( .A(n101101), .B(n10142), .S0(n8833), .Y(n4400) );
  MXI2X1 U6511 ( .A(n10109), .B(n10141), .S0(n8833), .Y(n4399) );
  MXI2X1 U6512 ( .A(n10108), .B(n10140), .S0(n8833), .Y(n4398) );
  MXI2X1 U6513 ( .A(n10107), .B(n10139), .S0(n8833), .Y(n4397) );
  MXI2X1 U6514 ( .A(n10106), .B(n10138), .S0(n8833), .Y(n4396) );
  MXI2X1 U6515 ( .A(n10105), .B(n10137), .S0(n8833), .Y(n4395) );
  MXI2X1 U6516 ( .A(n10104), .B(n10136), .S0(n8833), .Y(n4394) );
  MXI2X1 U6517 ( .A(n10103), .B(n10135), .S0(n8833), .Y(n4393) );
  MXI2X1 U6518 ( .A(n10102), .B(n10134), .S0(n8833), .Y(n4392) );
  MXI2X1 U6519 ( .A(n10101), .B(n10133), .S0(n8832), .Y(n4391) );
  MXI2X1 U6520 ( .A(n10100), .B(n10132), .S0(n8832), .Y(n4390) );
  MXI2X1 U6521 ( .A(n10099), .B(n10131), .S0(n8832), .Y(n4389) );
  MXI2X1 U6522 ( .A(n10098), .B(n10130), .S0(n8832), .Y(n4388) );
  MXI2X1 U6523 ( .A(n10097), .B(n10129), .S0(n8832), .Y(n4387) );
  MXI2X1 U6524 ( .A(n10096), .B(n10128), .S0(n8832), .Y(n4386) );
  MXI2X1 U6525 ( .A(n10095), .B(n10127), .S0(n8832), .Y(n4385) );
  MXI2X1 U6526 ( .A(n10094), .B(n10126), .S0(n8832), .Y(n4384) );
  MXI2X1 U6527 ( .A(n10093), .B(n10125), .S0(n8832), .Y(n4383) );
  MXI2X1 U6528 ( .A(n10092), .B(n10124), .S0(n8832), .Y(n4382) );
  MXI2X1 U6529 ( .A(n10091), .B(n10123), .S0(n8832), .Y(n4381) );
  MXI2X1 U6530 ( .A(n10090), .B(n10122), .S0(n8832), .Y(n4380) );
  MXI2X1 U6531 ( .A(n10089), .B(n10121), .S0(n8832), .Y(n4379) );
  MXI2X1 U6532 ( .A(n10088), .B(n10120), .S0(n8831), .Y(n4378) );
  MXI2X1 U6533 ( .A(n10087), .B(n10119), .S0(n8831), .Y(n4377) );
  MXI2X1 U6534 ( .A(n10086), .B(n10118), .S0(n8831), .Y(n4376) );
  MXI2X1 U6535 ( .A(n10085), .B(n10117), .S0(n8831), .Y(n4375) );
  MXI2X1 U6536 ( .A(n10084), .B(n10116), .S0(n8831), .Y(n4374) );
  MXI2X1 U6537 ( .A(n10083), .B(n10115), .S0(n8831), .Y(n4373) );
  MXI2X1 U6538 ( .A(n10082), .B(n10114), .S0(n8831), .Y(n4372) );
  MXI2X1 U6539 ( .A(n10081), .B(n10113), .S0(n8831), .Y(n4371) );
  MXI2X1 U6540 ( .A(n10080), .B(n10112), .S0(n8831), .Y(n4370) );
  MXI2X1 U6541 ( .A(n10079), .B(n10111), .S0(n8831), .Y(n4369) );
  MXI2X1 U6542 ( .A(n10078), .B(n101101), .S0(n8831), .Y(n4368) );
  MXI2X1 U6543 ( .A(n10077), .B(n10109), .S0(n8831), .Y(n4367) );
  MXI2X1 U6544 ( .A(n10076), .B(n10108), .S0(n8831), .Y(n4366) );
  MXI2X1 U6545 ( .A(n10075), .B(n10107), .S0(n8830), .Y(n4365) );
  MXI2X1 U6546 ( .A(n10074), .B(n10106), .S0(n8830), .Y(n4364) );
  MXI2X1 U6547 ( .A(n10073), .B(n10105), .S0(n8830), .Y(n4363) );
  MXI2X1 U6548 ( .A(n10072), .B(n10104), .S0(n8830), .Y(n4362) );
  MXI2X1 U6549 ( .A(n10071), .B(n10103), .S0(n8830), .Y(n4361) );
  MXI2X1 U6550 ( .A(n10070), .B(n10102), .S0(n8830), .Y(n4360) );
  MXI2X1 U6551 ( .A(n10069), .B(n10101), .S0(n8830), .Y(n4359) );
  MXI2X1 U6552 ( .A(n10068), .B(n10100), .S0(n8830), .Y(n4358) );
  MXI2X1 U6553 ( .A(n10067), .B(n10099), .S0(n8830), .Y(n4357) );
  MXI2X1 U6554 ( .A(n10066), .B(n10098), .S0(n8830), .Y(n4356) );
  MXI2X1 U6555 ( .A(n10065), .B(n10097), .S0(n8830), .Y(n4355) );
  MXI2X1 U6556 ( .A(n10064), .B(n10096), .S0(n8830), .Y(n4354) );
  MXI2X1 U6557 ( .A(n10063), .B(n10095), .S0(n8830), .Y(n4353) );
  MXI2X1 U6558 ( .A(n10062), .B(n10094), .S0(n8829), .Y(n4352) );
  MXI2X1 U6559 ( .A(n10061), .B(n10093), .S0(n8829), .Y(n4351) );
  MXI2X1 U6560 ( .A(n10060), .B(n10092), .S0(n8829), .Y(n4350) );
  MXI2X1 U6561 ( .A(n10059), .B(n10091), .S0(n8829), .Y(n4349) );
  MXI2X1 U6562 ( .A(n10058), .B(n10090), .S0(n8829), .Y(n4348) );
  MXI2X1 U6563 ( .A(n10057), .B(n10089), .S0(n8829), .Y(n4347) );
  MXI2X1 U6564 ( .A(n10056), .B(n10088), .S0(n8829), .Y(n4346) );
  MXI2X1 U6565 ( .A(n10055), .B(n10087), .S0(n8829), .Y(n4345) );
  MXI2X1 U6566 ( .A(n10054), .B(n10086), .S0(n8829), .Y(n4344) );
  MXI2X1 U6567 ( .A(n10053), .B(n10085), .S0(n8829), .Y(n4343) );
  MXI2X1 U6568 ( .A(n10052), .B(n10084), .S0(n8829), .Y(n4342) );
  MXI2X1 U6569 ( .A(n10051), .B(n10083), .S0(n8829), .Y(n4341) );
  MXI2X1 U6570 ( .A(n10050), .B(n10082), .S0(n8829), .Y(n4340) );
  MXI2X1 U6571 ( .A(n10049), .B(n10081), .S0(n8828), .Y(n4339) );
  MXI2X1 U6572 ( .A(n10048), .B(n10080), .S0(n8828), .Y(n4338) );
  MXI2X1 U6573 ( .A(n10047), .B(n10079), .S0(n8828), .Y(n4337) );
  MXI2X1 U6574 ( .A(n10046), .B(n10078), .S0(n8828), .Y(n4336) );
  MXI2X1 U6575 ( .A(n10045), .B(n10077), .S0(n8828), .Y(n4335) );
  MXI2X1 U6576 ( .A(n10044), .B(n10076), .S0(n8828), .Y(n4334) );
  MXI2X1 U6577 ( .A(n10043), .B(n10075), .S0(n8828), .Y(n4333) );
  MXI2X1 U6578 ( .A(n10042), .B(n10074), .S0(n8828), .Y(n4332) );
  MXI2X1 U6579 ( .A(n10041), .B(n10073), .S0(n8828), .Y(n4331) );
  MXI2X1 U6580 ( .A(n10040), .B(n10072), .S0(n8828), .Y(n4330) );
  MXI2X1 U6581 ( .A(n10039), .B(n10071), .S0(n8828), .Y(n4329) );
  MXI2X1 U6582 ( .A(n10038), .B(n10070), .S0(n8828), .Y(n4328) );
  MXI2X1 U6583 ( .A(n10037), .B(n10069), .S0(n8828), .Y(n4327) );
  MXI2X1 U6584 ( .A(n10036), .B(n10068), .S0(n8827), .Y(n4326) );
  MXI2X1 U6585 ( .A(n10035), .B(n10067), .S0(n8827), .Y(n4325) );
  MXI2X1 U6586 ( .A(n10034), .B(n10066), .S0(n8827), .Y(n4324) );
  MXI2X1 U6587 ( .A(n10033), .B(n10065), .S0(n8827), .Y(n4323) );
  MXI2X1 U6588 ( .A(n10032), .B(n10064), .S0(n8827), .Y(n4322) );
  MXI2X1 U6589 ( .A(n10031), .B(n10063), .S0(n8827), .Y(n4321) );
  MXI2X1 U6590 ( .A(n10030), .B(n10062), .S0(n8827), .Y(n4320) );
  MXI2X1 U6591 ( .A(n10029), .B(n10061), .S0(n8827), .Y(n4319) );
  MXI2X1 U6592 ( .A(n10028), .B(n10060), .S0(n8827), .Y(n4318) );
  MXI2X1 U6593 ( .A(n10027), .B(n10059), .S0(n8827), .Y(n4317) );
  MXI2X1 U6594 ( .A(n10026), .B(n10058), .S0(n8827), .Y(n4316) );
  MXI2X1 U6595 ( .A(n10025), .B(n10057), .S0(n8827), .Y(n4315) );
  MXI2X1 U6596 ( .A(n10024), .B(n10056), .S0(n8827), .Y(n4314) );
  MXI2X1 U6597 ( .A(n10023), .B(n10055), .S0(n8826), .Y(n4313) );
  MXI2X1 U6598 ( .A(n10022), .B(n10054), .S0(n8826), .Y(n4312) );
  MXI2X1 U6599 ( .A(n10021), .B(n10053), .S0(n8826), .Y(n4311) );
  MXI2X1 U6600 ( .A(n10020), .B(n10052), .S0(n8826), .Y(n4310) );
  MXI2X1 U6601 ( .A(n10019), .B(n10051), .S0(n8826), .Y(n4309) );
  MXI2X1 U6602 ( .A(n10018), .B(n10050), .S0(n8826), .Y(n4308) );
  MXI2X1 U6603 ( .A(n10017), .B(n10049), .S0(n8826), .Y(n4307) );
  MXI2X1 U6604 ( .A(n10016), .B(n10048), .S0(n8826), .Y(n4306) );
  MXI2X1 U6605 ( .A(n10015), .B(n10047), .S0(n8826), .Y(n4305) );
  MXI2X1 U6606 ( .A(n10014), .B(n10046), .S0(n8826), .Y(n4304) );
  MXI2X1 U6607 ( .A(n10013), .B(n10045), .S0(n8826), .Y(n4303) );
  MXI2X1 U6608 ( .A(n10012), .B(n10044), .S0(n8826), .Y(n4302) );
  MXI2X1 U6609 ( .A(n10011), .B(n10043), .S0(n8826), .Y(n4301) );
  MXI2X1 U6610 ( .A(n10010), .B(n10042), .S0(n8825), .Y(n4300) );
  MXI2X1 U6611 ( .A(n10009), .B(n10041), .S0(n8825), .Y(n4299) );
  MXI2X1 U6612 ( .A(n10008), .B(n10040), .S0(n8825), .Y(n4298) );
  MXI2X1 U6613 ( .A(n10007), .B(n10039), .S0(n8825), .Y(n4297) );
  MXI2X1 U6614 ( .A(n10006), .B(n10038), .S0(n8825), .Y(n4296) );
  MXI2X1 U6615 ( .A(n10005), .B(n10037), .S0(n8825), .Y(n4295) );
  MXI2X1 U6616 ( .A(n10004), .B(n10036), .S0(n8825), .Y(n4294) );
  MXI2X1 U6617 ( .A(n10003), .B(n10035), .S0(n8825), .Y(n4293) );
  MXI2X1 U6618 ( .A(n10002), .B(n10034), .S0(n8825), .Y(n4292) );
  MXI2X1 U6619 ( .A(n10001), .B(n10033), .S0(n8825), .Y(n4291) );
  MXI2X1 U6620 ( .A(n10000), .B(n10032), .S0(n8825), .Y(n4290) );
  MXI2X1 U6621 ( .A(n9999), .B(n10031), .S0(n8825), .Y(n4289) );
  MXI2X1 U6622 ( .A(n9998), .B(n10030), .S0(n8825), .Y(n4288) );
  MXI2X1 U6623 ( .A(n9997), .B(n10029), .S0(n8824), .Y(n4287) );
  MXI2X1 U6624 ( .A(n9996), .B(n10028), .S0(n8824), .Y(n4286) );
  MXI2X1 U6625 ( .A(n9995), .B(n10027), .S0(n8824), .Y(n4285) );
  MXI2X1 U6626 ( .A(n9994), .B(n10026), .S0(n8824), .Y(n4284) );
  MXI2X1 U6627 ( .A(n9993), .B(n10025), .S0(n8824), .Y(n4283) );
  MXI2X1 U6628 ( .A(n9992), .B(n10024), .S0(n8824), .Y(n4282) );
  MXI2X1 U6629 ( .A(n9991), .B(n10023), .S0(n8824), .Y(n4281) );
  MXI2X1 U6630 ( .A(n9990), .B(n10022), .S0(n8824), .Y(n4280) );
  MXI2X1 U6631 ( .A(n9989), .B(n10021), .S0(n8824), .Y(n4279) );
  MXI2X1 U6632 ( .A(n9988), .B(n10020), .S0(n8824), .Y(n4278) );
  MXI2X1 U6633 ( .A(n9987), .B(n10019), .S0(n8824), .Y(n4277) );
  MXI2X1 U6634 ( .A(n9986), .B(n10018), .S0(n8824), .Y(n4276) );
  MXI2X1 U6635 ( .A(n9985), .B(n10017), .S0(n8824), .Y(n4275) );
  MXI2X1 U6636 ( .A(n9984), .B(n10016), .S0(n8823), .Y(n4274) );
  MXI2X1 U6637 ( .A(n9983), .B(n10015), .S0(n8823), .Y(n4273) );
  MXI2X1 U6638 ( .A(n9982), .B(n10014), .S0(n8823), .Y(n4272) );
  MXI2X1 U6639 ( .A(n9981), .B(n10013), .S0(n8823), .Y(n4271) );
  MXI2X1 U6640 ( .A(n9980), .B(n10012), .S0(n8823), .Y(n4270) );
  MXI2X1 U6641 ( .A(n9979), .B(n10011), .S0(n8823), .Y(n4269) );
  MXI2X1 U6642 ( .A(n9978), .B(n10010), .S0(n8823), .Y(n4268) );
  MXI2X1 U6643 ( .A(n9977), .B(n10009), .S0(n8823), .Y(n4267) );
  MXI2X1 U6644 ( .A(n9976), .B(n10008), .S0(n8823), .Y(n4266) );
  MXI2X1 U6645 ( .A(n9975), .B(n10007), .S0(n8823), .Y(n4265) );
  MXI2X1 U6646 ( .A(n9974), .B(n10006), .S0(n8823), .Y(n4264) );
  MXI2X1 U6647 ( .A(n9973), .B(n10005), .S0(n8823), .Y(n4263) );
  MXI2X1 U6648 ( .A(n9972), .B(n10004), .S0(n8823), .Y(n4262) );
  MXI2X1 U6649 ( .A(n9971), .B(n10003), .S0(n8822), .Y(n4261) );
  MXI2X1 U6650 ( .A(n9970), .B(n10002), .S0(n8822), .Y(n4260) );
  MXI2X1 U6651 ( .A(n9969), .B(n10001), .S0(n8822), .Y(n4259) );
  MXI2X1 U6652 ( .A(n9968), .B(n10000), .S0(n8822), .Y(n4258) );
  MXI2X1 U6653 ( .A(n9967), .B(n9999), .S0(n8822), .Y(n4257) );
  MXI2X1 U6654 ( .A(n9966), .B(n9998), .S0(n8822), .Y(n4256) );
  MXI2X1 U6655 ( .A(n9965), .B(n9997), .S0(n8822), .Y(n4255) );
  MXI2X1 U6656 ( .A(n9964), .B(n9996), .S0(n8822), .Y(n4254) );
  MXI2X1 U6657 ( .A(n9963), .B(n9995), .S0(n8822), .Y(n4253) );
  MXI2X1 U6658 ( .A(n9962), .B(n9994), .S0(n8822), .Y(n4252) );
  MXI2X1 U6659 ( .A(n9961), .B(n9993), .S0(n8822), .Y(n4251) );
  MXI2X1 U6660 ( .A(n9960), .B(n9992), .S0(n8822), .Y(n4250) );
  MXI2X1 U6661 ( .A(n9959), .B(n9991), .S0(n8822), .Y(n4249) );
  MXI2X1 U6662 ( .A(n9958), .B(n9990), .S0(n8821), .Y(n4248) );
  MXI2X1 U6663 ( .A(n9957), .B(n9989), .S0(n8821), .Y(n4247) );
  MXI2X1 U6664 ( .A(n9956), .B(n9988), .S0(n8821), .Y(n4246) );
  MXI2X1 U6665 ( .A(n9955), .B(n9987), .S0(n8821), .Y(n4245) );
  MXI2X1 U6666 ( .A(n9954), .B(n9986), .S0(n8821), .Y(n4244) );
  MXI2X1 U6667 ( .A(n9953), .B(n9985), .S0(n8821), .Y(n4243) );
  MXI2X1 U6668 ( .A(n9952), .B(n9984), .S0(n8821), .Y(n4242) );
  MXI2X1 U6669 ( .A(n9951), .B(n9983), .S0(n8821), .Y(n4241) );
  MXI2X1 U6670 ( .A(n9950), .B(n9982), .S0(n8821), .Y(n4240) );
  MXI2X1 U6671 ( .A(n9949), .B(n9981), .S0(n8821), .Y(n4239) );
  MXI2X1 U6672 ( .A(n9948), .B(n9980), .S0(n8821), .Y(n4238) );
  MXI2X1 U6673 ( .A(n9947), .B(n9979), .S0(n8821), .Y(n4237) );
  MXI2X1 U6674 ( .A(n9946), .B(n9978), .S0(n8821), .Y(n4236) );
  MXI2X1 U6675 ( .A(n9945), .B(n9977), .S0(n8820), .Y(n4235) );
  MXI2X1 U6676 ( .A(n9944), .B(n9976), .S0(n8820), .Y(n4234) );
  MXI2X1 U6677 ( .A(n9943), .B(n9975), .S0(n8820), .Y(n4233) );
  MXI2X1 U6678 ( .A(n9942), .B(n9974), .S0(n8820), .Y(n4232) );
  MXI2X1 U6679 ( .A(n9941), .B(n9973), .S0(n8820), .Y(n4231) );
  MXI2X1 U6680 ( .A(n9940), .B(n9972), .S0(n8820), .Y(n4230) );
  MXI2X1 U6681 ( .A(n9939), .B(n9971), .S0(n8820), .Y(n4229) );
  MXI2X1 U6682 ( .A(n9938), .B(n9970), .S0(n8820), .Y(n4228) );
  MXI2X1 U6683 ( .A(n9937), .B(n9969), .S0(n8820), .Y(n4227) );
  MXI2X1 U6684 ( .A(n9936), .B(n9968), .S0(n8820), .Y(n4226) );
  MXI2X1 U6685 ( .A(n9935), .B(n9967), .S0(n8820), .Y(n4225) );
  MXI2X1 U6686 ( .A(n9934), .B(n9966), .S0(n8820), .Y(n4224) );
  MXI2X1 U6687 ( .A(n9933), .B(n9965), .S0(n8820), .Y(n4223) );
  MXI2X1 U6688 ( .A(n9932), .B(n9964), .S0(n8819), .Y(n4222) );
  MXI2X1 U6689 ( .A(n9931), .B(n9963), .S0(n8819), .Y(n4221) );
  MXI2X1 U6690 ( .A(n9930), .B(n9962), .S0(n8819), .Y(n4220) );
  MXI2X1 U6691 ( .A(n9929), .B(n9961), .S0(n8819), .Y(n4219) );
  MXI2X1 U6692 ( .A(n9928), .B(n9960), .S0(n8819), .Y(n4218) );
  MXI2X1 U6693 ( .A(n9927), .B(n9959), .S0(n8819), .Y(n4217) );
  MXI2X1 U6694 ( .A(n9926), .B(n9958), .S0(n8819), .Y(n4216) );
  MXI2X1 U6695 ( .A(n9925), .B(n9957), .S0(n8819), .Y(n4215) );
  MXI2X1 U6696 ( .A(n9924), .B(n9956), .S0(n8819), .Y(n4214) );
  MXI2X1 U6697 ( .A(n9923), .B(n9955), .S0(n8819), .Y(n4213) );
  MXI2X1 U6698 ( .A(n9922), .B(n9954), .S0(n8819), .Y(n4212) );
  MXI2X1 U6699 ( .A(n9921), .B(n9953), .S0(n8819), .Y(n4211) );
  MXI2X1 U6700 ( .A(n9920), .B(n9952), .S0(n8819), .Y(n4210) );
  MXI2X1 U6701 ( .A(n9919), .B(n9951), .S0(n8818), .Y(n4209) );
  MXI2X1 U6702 ( .A(n9918), .B(n9950), .S0(n8818), .Y(n4208) );
  MXI2X1 U6703 ( .A(n9917), .B(n9949), .S0(n8818), .Y(n4207) );
  MXI2X1 U6704 ( .A(n9916), .B(n9948), .S0(n8818), .Y(n4206) );
  MXI2X1 U6705 ( .A(n9915), .B(n9947), .S0(n8818), .Y(n4205) );
  MXI2X1 U6706 ( .A(n9914), .B(n9946), .S0(n8818), .Y(n4204) );
  MXI2X1 U6707 ( .A(n9913), .B(n9945), .S0(n8818), .Y(n4203) );
  MXI2X1 U6708 ( .A(n9912), .B(n9944), .S0(n8818), .Y(n4202) );
  MXI2X1 U6709 ( .A(n9911), .B(n9943), .S0(n8818), .Y(n4201) );
  MXI2X1 U6710 ( .A(n9910), .B(n9942), .S0(n8818), .Y(n4200) );
  MXI2X1 U6711 ( .A(n9909), .B(n9941), .S0(n8818), .Y(n4199) );
  MXI2X1 U6712 ( .A(n9908), .B(n9940), .S0(n8818), .Y(n4198) );
  MXI2X1 U6713 ( .A(n9907), .B(n9939), .S0(n8818), .Y(n4197) );
  MXI2X1 U6714 ( .A(n9906), .B(n9938), .S0(n8817), .Y(n4196) );
  MXI2X1 U6715 ( .A(n9905), .B(n9937), .S0(n8817), .Y(n4195) );
  MXI2X1 U6716 ( .A(n9904), .B(n9936), .S0(n8817), .Y(n4194) );
  MXI2X1 U6717 ( .A(n9903), .B(n9935), .S0(n8817), .Y(n4193) );
  MXI2X1 U6718 ( .A(n9902), .B(n9934), .S0(n8817), .Y(n4192) );
  MXI2X1 U6719 ( .A(n9901), .B(n9933), .S0(n8817), .Y(n4191) );
  MXI2X1 U6720 ( .A(n9900), .B(n9932), .S0(n8817), .Y(n4190) );
  MXI2X1 U6721 ( .A(n9899), .B(n9931), .S0(n8817), .Y(n4189) );
  MXI2X1 U6722 ( .A(n9898), .B(n9930), .S0(n8817), .Y(n4188) );
  MXI2X1 U6723 ( .A(n9897), .B(n9929), .S0(n8817), .Y(n4187) );
  MXI2X1 U6724 ( .A(n9896), .B(n9928), .S0(n8817), .Y(n4186) );
  MXI2X1 U6725 ( .A(n9895), .B(n9927), .S0(n8817), .Y(n4185) );
  MXI2X1 U6726 ( .A(n9894), .B(n9926), .S0(n8817), .Y(n4184) );
  MXI2X1 U6727 ( .A(n9893), .B(n9925), .S0(n8816), .Y(n4183) );
  MXI2X1 U6728 ( .A(n9892), .B(n9924), .S0(n8816), .Y(n4182) );
  MXI2X1 U6729 ( .A(n9891), .B(n9923), .S0(n8816), .Y(n4181) );
  MXI2X1 U6730 ( .A(n9890), .B(n9922), .S0(n8816), .Y(n4180) );
  MXI2X1 U6731 ( .A(n9889), .B(n9921), .S0(n8816), .Y(n4179) );
  MXI2X1 U6732 ( .A(n9888), .B(n9920), .S0(n8816), .Y(n4178) );
  MXI2X1 U6733 ( .A(n9887), .B(n9919), .S0(n8816), .Y(n4177) );
  MXI2X1 U6734 ( .A(n9886), .B(n9918), .S0(n8816), .Y(n4176) );
  MXI2X1 U6735 ( .A(n9885), .B(n9917), .S0(n8816), .Y(n4175) );
  MXI2X1 U6736 ( .A(n9884), .B(n9916), .S0(n8816), .Y(n4174) );
  MXI2X1 U6737 ( .A(n9883), .B(n9915), .S0(n8816), .Y(n4173) );
  MXI2X1 U6738 ( .A(n9882), .B(n9914), .S0(n8816), .Y(n4172) );
  MXI2X1 U6739 ( .A(n9881), .B(n9913), .S0(n8816), .Y(n4171) );
  MXI2X1 U6740 ( .A(n9880), .B(n9912), .S0(n8815), .Y(n4170) );
  MXI2X1 U6741 ( .A(n9879), .B(n9911), .S0(n8815), .Y(n4169) );
  MXI2X1 U6742 ( .A(n9878), .B(n9910), .S0(n8815), .Y(n4168) );
  MXI2X1 U6743 ( .A(n9877), .B(n9909), .S0(n8815), .Y(n4167) );
  MXI2X1 U6744 ( .A(n9876), .B(n9908), .S0(n8815), .Y(n4166) );
  MXI2X1 U6745 ( .A(n9875), .B(n9907), .S0(n8815), .Y(n4165) );
  MXI2X1 U6746 ( .A(n9874), .B(n9906), .S0(n8815), .Y(n4164) );
  MXI2X1 U6747 ( .A(n9873), .B(n9905), .S0(n8815), .Y(n4163) );
  MXI2X1 U6748 ( .A(n9872), .B(n9904), .S0(n8815), .Y(n4162) );
  MXI2X1 U6749 ( .A(n9871), .B(n9903), .S0(n8815), .Y(n4161) );
  MXI2X1 U6750 ( .A(n9870), .B(n9902), .S0(n8815), .Y(n4160) );
  MXI2X1 U6751 ( .A(n9869), .B(n9901), .S0(n8815), .Y(n4159) );
  MXI2X1 U6752 ( .A(n9868), .B(n9900), .S0(n8815), .Y(n4158) );
  MXI2X1 U6753 ( .A(n9867), .B(n9899), .S0(n8814), .Y(n4157) );
  MXI2X1 U6754 ( .A(n9866), .B(n9898), .S0(n8814), .Y(n4156) );
  MXI2X1 U6755 ( .A(n9865), .B(n9897), .S0(n8814), .Y(n4155) );
  MXI2X1 U6756 ( .A(n9864), .B(n9896), .S0(n8814), .Y(n4154) );
  MXI2X1 U6757 ( .A(n9863), .B(n9895), .S0(n8814), .Y(n4153) );
  MXI2X1 U6758 ( .A(n9862), .B(n9894), .S0(n8814), .Y(n4152) );
  MXI2X1 U6759 ( .A(n9861), .B(n9893), .S0(n8814), .Y(n4151) );
  MXI2X1 U6760 ( .A(n9860), .B(n9892), .S0(n8814), .Y(n4150) );
  MXI2X1 U6761 ( .A(n9859), .B(n9891), .S0(n8814), .Y(n4149) );
  MXI2X1 U6762 ( .A(n9858), .B(n9890), .S0(n8814), .Y(n4148) );
  MXI2X1 U6763 ( .A(n9857), .B(n9889), .S0(n8814), .Y(n4147) );
  MXI2X1 U6764 ( .A(n9856), .B(n9888), .S0(n8814), .Y(n4146) );
  MXI2X1 U6765 ( .A(n9855), .B(n9887), .S0(n8814), .Y(n4145) );
  MXI2X1 U6766 ( .A(n9854), .B(n9886), .S0(n8813), .Y(n4144) );
  MXI2X1 U6767 ( .A(n9853), .B(n9885), .S0(n8813), .Y(n4143) );
  MXI2X1 U6768 ( .A(n9852), .B(n9884), .S0(n8813), .Y(n4142) );
  MXI2X1 U6769 ( .A(n9851), .B(n9883), .S0(n8813), .Y(n4141) );
  MXI2X1 U6770 ( .A(n9850), .B(n9882), .S0(n8813), .Y(n4140) );
  MXI2X1 U6771 ( .A(n9849), .B(n9881), .S0(n8813), .Y(n4139) );
  MXI2X1 U6772 ( .A(n9848), .B(n9880), .S0(n8813), .Y(n4138) );
  MXI2X1 U6773 ( .A(n9847), .B(n9879), .S0(n8813), .Y(n4137) );
  MXI2X1 U6774 ( .A(n9846), .B(n9878), .S0(n8813), .Y(n4136) );
  MXI2X1 U6775 ( .A(n9845), .B(n9877), .S0(n8813), .Y(n4135) );
  MXI2X1 U6776 ( .A(n9844), .B(n9876), .S0(n8813), .Y(n4134) );
  MXI2X1 U6777 ( .A(n9843), .B(n9875), .S0(n8813), .Y(n4133) );
  MXI2X1 U6778 ( .A(n9842), .B(n9874), .S0(n8813), .Y(n4132) );
  MXI2X1 U6779 ( .A(n9841), .B(n9873), .S0(n8812), .Y(n4131) );
  MXI2X1 U6780 ( .A(n9840), .B(n9872), .S0(n8812), .Y(n4130) );
  MXI2X1 U6781 ( .A(n9839), .B(n9871), .S0(n8812), .Y(n4129) );
  MXI2X1 U6782 ( .A(n9838), .B(n9870), .S0(n8812), .Y(n4128) );
  MXI2X1 U6783 ( .A(n9837), .B(n9869), .S0(n8812), .Y(n4127) );
  MXI2X1 U6784 ( .A(n9836), .B(n9868), .S0(n8812), .Y(n4126) );
  MXI2X1 U6785 ( .A(n9835), .B(n9867), .S0(n8812), .Y(n4125) );
  MXI2X1 U6786 ( .A(n9834), .B(n9866), .S0(n8812), .Y(n4124) );
  MXI2X1 U6787 ( .A(n9833), .B(n9865), .S0(n8812), .Y(n4123) );
  MXI2X1 U6788 ( .A(n9832), .B(n9864), .S0(n8812), .Y(n4122) );
  MXI2X1 U6789 ( .A(n9831), .B(n9863), .S0(n8812), .Y(n4121) );
  MXI2X1 U6790 ( .A(n9830), .B(n9862), .S0(n8812), .Y(n4120) );
  MXI2X1 U6791 ( .A(n9829), .B(n9861), .S0(n8812), .Y(n4119) );
  MXI2X1 U6792 ( .A(n9828), .B(n9860), .S0(n8811), .Y(n4118) );
  MXI2X1 U6793 ( .A(n9827), .B(n9859), .S0(n8811), .Y(n4117) );
  MXI2X1 U6794 ( .A(n9826), .B(n9858), .S0(n8811), .Y(n4116) );
  MXI2X1 U6795 ( .A(n9825), .B(n9857), .S0(n8811), .Y(n4115) );
  MXI2X1 U6796 ( .A(n9824), .B(n9856), .S0(n8811), .Y(n4114) );
  MXI2X1 U6797 ( .A(n9823), .B(n9855), .S0(n8811), .Y(n4113) );
  MXI2X1 U6798 ( .A(n9822), .B(n9854), .S0(n8811), .Y(n4112) );
  MXI2X1 U6799 ( .A(n9821), .B(n9853), .S0(n8811), .Y(n4111) );
  MXI2X1 U6800 ( .A(n9820), .B(n9852), .S0(n8811), .Y(n4110) );
  MXI2X1 U6801 ( .A(n9819), .B(n9851), .S0(n8811), .Y(n4109) );
  MXI2X1 U6802 ( .A(n9818), .B(n9850), .S0(n8811), .Y(n4108) );
  MXI2X1 U6803 ( .A(n9817), .B(n9849), .S0(n8811), .Y(n4107) );
  MXI2X1 U6804 ( .A(n9816), .B(n9848), .S0(n8811), .Y(n4106) );
  MXI2X1 U6805 ( .A(n9815), .B(n9847), .S0(n8810), .Y(n4105) );
  MXI2X1 U6806 ( .A(n9814), .B(n9846), .S0(n8810), .Y(n4104) );
  MXI2X1 U6807 ( .A(n9813), .B(n9845), .S0(n8810), .Y(n4103) );
  MXI2X1 U6808 ( .A(n9812), .B(n9844), .S0(n8810), .Y(n4102) );
  MXI2X1 U6809 ( .A(n9811), .B(n9843), .S0(n8810), .Y(n4101) );
  MXI2X1 U6810 ( .A(n9810), .B(n9842), .S0(n8810), .Y(n4100) );
  MXI2X1 U6811 ( .A(n9809), .B(n9841), .S0(n8810), .Y(n4099) );
  MXI2X1 U6812 ( .A(n9808), .B(n9840), .S0(n8810), .Y(n4098) );
  MXI2X1 U6813 ( .A(n9807), .B(n9839), .S0(n8810), .Y(n4097) );
  MXI2X1 U6814 ( .A(n9806), .B(n9838), .S0(n8810), .Y(n4096) );
  MXI2X1 U6815 ( .A(n9805), .B(n9837), .S0(n8810), .Y(n4095) );
  MXI2X1 U6816 ( .A(n9804), .B(n9836), .S0(n8810), .Y(n4094) );
  MXI2X1 U6817 ( .A(n9803), .B(n9835), .S0(n8810), .Y(n4093) );
  MXI2X1 U6818 ( .A(n9802), .B(n9834), .S0(n8809), .Y(n4092) );
  MXI2X1 U6819 ( .A(n9801), .B(n9833), .S0(n8809), .Y(n4091) );
  MXI2X1 U6820 ( .A(n9800), .B(n9832), .S0(n8809), .Y(n4090) );
  MXI2X1 U6821 ( .A(n9799), .B(n9831), .S0(n8809), .Y(n4089) );
  MXI2X1 U6822 ( .A(n9798), .B(n9830), .S0(n8809), .Y(n4088) );
  MXI2X1 U6823 ( .A(n9797), .B(n9829), .S0(n8809), .Y(n4087) );
  MXI2X1 U6824 ( .A(n9796), .B(n9828), .S0(n8809), .Y(n4086) );
  MXI2X1 U6825 ( .A(n9795), .B(n9827), .S0(n8809), .Y(n4085) );
  MXI2X1 U6826 ( .A(n9794), .B(n9826), .S0(n8809), .Y(n4084) );
  MXI2X1 U6827 ( .A(n9793), .B(n9825), .S0(n8809), .Y(n4083) );
  MXI2X1 U6828 ( .A(n9792), .B(n9824), .S0(n8809), .Y(n4082) );
  MXI2X1 U6829 ( .A(n9791), .B(n9823), .S0(n8809), .Y(n4081) );
  MXI2X1 U6830 ( .A(n9790), .B(n9822), .S0(n8809), .Y(n4080) );
  MXI2X1 U6831 ( .A(n9789), .B(n9821), .S0(n8808), .Y(n4079) );
  MXI2X1 U6832 ( .A(n9788), .B(n9820), .S0(n8808), .Y(n4078) );
  MXI2X1 U6833 ( .A(n9787), .B(n9819), .S0(n8808), .Y(n4077) );
  MXI2X1 U6834 ( .A(n9786), .B(n9818), .S0(n8808), .Y(n4076) );
  MXI2X1 U6835 ( .A(n9785), .B(n9817), .S0(n8808), .Y(n4075) );
  MXI2X1 U6836 ( .A(n9784), .B(n9816), .S0(n8808), .Y(n4074) );
  MXI2X1 U6837 ( .A(n9783), .B(n9815), .S0(n8808), .Y(n4073) );
  MXI2X1 U6838 ( .A(n9782), .B(n9814), .S0(n8808), .Y(n4072) );
  MXI2X1 U6839 ( .A(n9781), .B(n9813), .S0(n8808), .Y(n4071) );
  MXI2X1 U6840 ( .A(n9780), .B(n9812), .S0(n8808), .Y(n4070) );
  MXI2X1 U6841 ( .A(n9779), .B(n9811), .S0(n8808), .Y(n4069) );
  MXI2X1 U6842 ( .A(n9778), .B(n9810), .S0(n8808), .Y(n4068) );
  MXI2X1 U6843 ( .A(n9777), .B(n9809), .S0(n8808), .Y(n4067) );
  MXI2X1 U6844 ( .A(n9776), .B(n9808), .S0(n8807), .Y(n4066) );
  MXI2X1 U6845 ( .A(n9775), .B(n9807), .S0(n8807), .Y(n4065) );
  MXI2X1 U6846 ( .A(n9774), .B(n9806), .S0(n8807), .Y(n4064) );
  MXI2X1 U6847 ( .A(n9773), .B(n9805), .S0(n8807), .Y(n4063) );
  MXI2X1 U6848 ( .A(n9772), .B(n9804), .S0(n8807), .Y(n4062) );
  MXI2X1 U6849 ( .A(n9771), .B(n9803), .S0(n8807), .Y(n4061) );
  MXI2X1 U6850 ( .A(n9770), .B(n9802), .S0(n8807), .Y(n4060) );
  MXI2X1 U6851 ( .A(n9769), .B(n9801), .S0(n8807), .Y(n4059) );
  MXI2X1 U6852 ( .A(n9768), .B(n9800), .S0(n8807), .Y(n4058) );
  MXI2X1 U6853 ( .A(n9767), .B(n9799), .S0(n8807), .Y(n4057) );
  MXI2X1 U6854 ( .A(n9766), .B(n9798), .S0(n8807), .Y(n4056) );
  MXI2X1 U6855 ( .A(n9765), .B(n9797), .S0(n8807), .Y(n4055) );
  MXI2X1 U6856 ( .A(n9764), .B(n9796), .S0(n8807), .Y(n4054) );
  MXI2X1 U6857 ( .A(n9763), .B(n9795), .S0(n8806), .Y(n4053) );
  MXI2X1 U6858 ( .A(n9762), .B(n9794), .S0(n8806), .Y(n4052) );
  MXI2X1 U6859 ( .A(n9761), .B(n9793), .S0(n8806), .Y(n4051) );
  MXI2X1 U6860 ( .A(n9760), .B(n9792), .S0(n8806), .Y(n4050) );
  MXI2X1 U6861 ( .A(n9759), .B(n9791), .S0(n8806), .Y(n4049) );
  MXI2X1 U6862 ( .A(n9758), .B(n9790), .S0(n8806), .Y(n4048) );
  MXI2X1 U6863 ( .A(n9757), .B(n9789), .S0(n8806), .Y(n4047) );
  MXI2X1 U6864 ( .A(n9756), .B(n9788), .S0(n8806), .Y(n4046) );
  MXI2X1 U6865 ( .A(n9755), .B(n9787), .S0(n8806), .Y(n4045) );
  MXI2X1 U6866 ( .A(n9754), .B(n9786), .S0(n8806), .Y(n4044) );
  MXI2X1 U6867 ( .A(n9753), .B(n9785), .S0(n8806), .Y(n4043) );
  MXI2X1 U6868 ( .A(n9752), .B(n9784), .S0(n8806), .Y(n4042) );
  MXI2X1 U6869 ( .A(n9751), .B(n9783), .S0(n8806), .Y(n4041) );
  MXI2X1 U6870 ( .A(n9750), .B(n9782), .S0(n8805), .Y(n4040) );
  MXI2X1 U6871 ( .A(n9749), .B(n9781), .S0(n8805), .Y(n4039) );
  MXI2X1 U6872 ( .A(n9748), .B(n9780), .S0(n8805), .Y(n4038) );
  MXI2X1 U6873 ( .A(n9747), .B(n9779), .S0(n8805), .Y(n4037) );
  MXI2X1 U6874 ( .A(n9746), .B(n9778), .S0(n8805), .Y(n4036) );
  MXI2X1 U6875 ( .A(n9745), .B(n9777), .S0(n8805), .Y(n4035) );
  MXI2X1 U6876 ( .A(n9744), .B(n9776), .S0(n8805), .Y(n4034) );
  MXI2X1 U6877 ( .A(n9743), .B(n9775), .S0(n8805), .Y(n4033) );
  MXI2X1 U6878 ( .A(n9742), .B(n9774), .S0(n8805), .Y(n4032) );
  MXI2X1 U6879 ( .A(n9741), .B(n9773), .S0(n8805), .Y(n4031) );
  MXI2X1 U6880 ( .A(n9740), .B(n9772), .S0(n8805), .Y(n4030) );
  MXI2X1 U6881 ( .A(n9739), .B(n9771), .S0(n8805), .Y(n4029) );
  MXI2X1 U6882 ( .A(n9738), .B(n9770), .S0(n8805), .Y(n4028) );
  MXI2X1 U6883 ( .A(n9737), .B(n9769), .S0(n8834), .Y(n4027) );
  MXI2X1 U6884 ( .A(n9736), .B(n9768), .S0(n8835), .Y(n4026) );
  MXI2X1 U6885 ( .A(n9735), .B(n9767), .S0(n8836), .Y(n4025) );
  MXI2X1 U6886 ( .A(n9734), .B(n9766), .S0(n8833), .Y(n4024) );
  MXI2X1 U6887 ( .A(n9733), .B(n9765), .S0(n8822), .Y(n4023) );
  MXI2X1 U6888 ( .A(n9732), .B(n9764), .S0(n8823), .Y(n4022) );
  MXI2X1 U6889 ( .A(n9731), .B(n9763), .S0(n8824), .Y(n4021) );
  MXI2X1 U6890 ( .A(n9730), .B(n9762), .S0(n8825), .Y(n4020) );
  MXI2X1 U6891 ( .A(n9729), .B(n9761), .S0(n8826), .Y(n4019) );
  MXI2X1 U6892 ( .A(n9728), .B(n9760), .S0(n8827), .Y(n4018) );
  MXI2X1 U6893 ( .A(n9727), .B(n9759), .S0(n8810), .Y(n4017) );
  MXI2X1 U6894 ( .A(n9726), .B(n9758), .S0(n8811), .Y(n4016) );
  MXI2X1 U6895 ( .A(n9725), .B(n9757), .S0(n8812), .Y(n4015) );
  MXI2X1 U6896 ( .A(n9724), .B(n9756), .S0(n8804), .Y(n4014) );
  MXI2X1 U6897 ( .A(n9723), .B(n9755), .S0(n8804), .Y(n4013) );
  MXI2X1 U6898 ( .A(n9722), .B(n9754), .S0(n8804), .Y(n4012) );
  MXI2X1 U6899 ( .A(n9721), .B(n9753), .S0(n8804), .Y(n4011) );
  MXI2X1 U6900 ( .A(n9720), .B(n9752), .S0(n8804), .Y(n40101) );
  MXI2X1 U6901 ( .A(n9719), .B(n9751), .S0(n8804), .Y(n4009) );
  MXI2X1 U6902 ( .A(n9718), .B(n9750), .S0(n8804), .Y(n4008) );
  MXI2X1 U6903 ( .A(n9717), .B(n9749), .S0(n8804), .Y(n4007) );
  MXI2X1 U6904 ( .A(n9716), .B(n9748), .S0(n8804), .Y(n4006) );
  MXI2X1 U6905 ( .A(n9715), .B(n9747), .S0(n8804), .Y(n4005) );
  MXI2X1 U6906 ( .A(n9714), .B(n9746), .S0(n8804), .Y(n4004) );
  MXI2X1 U6907 ( .A(n9713), .B(n9745), .S0(n8804), .Y(n4003) );
  MXI2X1 U6908 ( .A(n9712), .B(n9744), .S0(n8804), .Y(n4002) );
  MXI2X1 U6909 ( .A(n9711), .B(n9743), .S0(n8803), .Y(n4001) );
  MXI2X1 U6910 ( .A(n9710), .B(n9742), .S0(n8803), .Y(n4000) );
  MXI2X1 U6911 ( .A(n9709), .B(n9741), .S0(n8803), .Y(n3999) );
  MXI2X1 U6912 ( .A(n9708), .B(n9740), .S0(n8803), .Y(n3998) );
  MXI2X1 U6913 ( .A(n9707), .B(n9739), .S0(n8803), .Y(n3997) );
  MXI2X1 U6914 ( .A(n9706), .B(n9738), .S0(n8803), .Y(n3996) );
  MXI2X1 U6915 ( .A(n9705), .B(n9737), .S0(n8803), .Y(n3995) );
  MXI2X1 U6916 ( .A(n9704), .B(n9736), .S0(n8803), .Y(n3994) );
  MXI2X1 U6917 ( .A(n9703), .B(n9735), .S0(n8803), .Y(n3993) );
  MXI2X1 U6918 ( .A(n9702), .B(n9734), .S0(n8803), .Y(n3992) );
  MXI2X1 U6919 ( .A(n9701), .B(n9733), .S0(n8803), .Y(n3991) );
  MXI2X1 U6920 ( .A(n9700), .B(n9732), .S0(n8803), .Y(n3990) );
  MXI2X1 U6921 ( .A(n9699), .B(n9731), .S0(n8803), .Y(n3989) );
  MXI2X1 U6922 ( .A(n9698), .B(n9730), .S0(n8813), .Y(n3988) );
  MXI2X1 U6923 ( .A(n9697), .B(n9729), .S0(n8814), .Y(n3987) );
  MXI2X1 U6924 ( .A(n9696), .B(n9728), .S0(n8815), .Y(n3986) );
  MXI2X1 U6925 ( .A(n9695), .B(n9727), .S0(n8816), .Y(n3985) );
  MXI2X1 U6926 ( .A(n9694), .B(n9726), .S0(n8817), .Y(n3984) );
  MXI2X1 U6927 ( .A(n9693), .B(n9725), .S0(n8818), .Y(n3983) );
  MXI2X1 U6928 ( .A(n9692), .B(n9724), .S0(n8819), .Y(n3982) );
  MXI2X1 U6929 ( .A(n9691), .B(n9723), .S0(n8820), .Y(n3981) );
  MXI2X1 U6930 ( .A(n9690), .B(n9722), .S0(n8821), .Y(n3980) );
  MXI2X1 U6931 ( .A(n9689), .B(n9721), .S0(n8805), .Y(n3979) );
  MXI2X1 U6932 ( .A(n9688), .B(n9720), .S0(n8806), .Y(n3978) );
  MXI2X1 U6933 ( .A(n9687), .B(n9719), .S0(n8807), .Y(n3977) );
  MXI2X1 U6934 ( .A(n9686), .B(n9718), .S0(n8808), .Y(n3976) );
  CLKINVX1 U6935 ( .A(data_valid), .Y(n9158) );
  OAI31XL U6936 ( .A0(n9174), .A1(n6068), .A2(n6067), .B0(n10475), .Y(n3462)
         );
  NAND2X1 U6937 ( .A(n9685), .B(n9501), .Y(n3461) );
  NAND4X1 U6938 ( .A(n9170), .B(n6191), .C(n6189), .D(n6193), .Y(n9501) );
  NOR2BX1 U6939 ( .AN(n9167), .B(n6072), .Y(n9170) );
  NOR3X1 U6940 ( .A(n6074), .B(n6075), .C(n6073), .Y(n9167) );
  NAND2X1 U6941 ( .A(n9502), .B(n9503), .Y(multiplier_r_6) );
  NAND2BX1 U6942 ( .AN(multiplier_r[14]), .B(n9504), .Y(multiplier_i_9) );
  NAND2BX1 U6943 ( .AN(multiplier_r[11]), .B(n9502), .Y(multiplier_r[14]) );
  NAND2X1 U6944 ( .A(n9505), .B(n9157), .Y(multiplier_r[11]) );
  NAND2BX1 U6945 ( .AN(multiplier_r_8), .B(n9505), .Y(multiplier_i_6) );
  NAND2BX1 U6946 ( .AN(multiplier_r[12]), .B(n9502), .Y(multiplier_r_8) );
  NAND2X1 U6947 ( .A(n9504), .B(n9506), .Y(multiplier_r[12]) );
  NAND2X1 U6948 ( .A(multiplier_r[16]), .B(n9505), .Y(multiplier_i_31) );
  NOR2X1 U6949 ( .A(n9507), .B(multiplier_r[13]), .Y(multiplier_r[16]) );
  NAND2X1 U6950 ( .A(n9502), .B(n9508), .Y(multiplier_r[13]) );
  NAND2BX1 U6951 ( .AN(multiplier_i_8), .B(n9157), .Y(multiplier_i_0) );
  NAND2X1 U6952 ( .A(n9502), .B(n9506), .Y(multiplier_i_8) );
  NAND2X1 U6953 ( .A(n9504), .B(n9503), .Y(multiplier_i[14]) );
  CLKINVX1 U6954 ( .A(multiplier_r_31), .Y(n9503) );
  NAND2X1 U6955 ( .A(n9505), .B(n9506), .Y(multiplier_r_31) );
  CLKINVX1 U6956 ( .A(n10480), .Y(n9506) );
  NOR2X1 U6957 ( .A(n9509), .B(n6072), .Y(n10480) );
  NAND2X1 U6958 ( .A(n9157), .B(n9502), .Y(multiplier_i[12]) );
  NAND3BX1 U6959 ( .AN(n6072), .B(n6075), .C(n6073), .Y(n9502) );
  NAND2X1 U6960 ( .A(n9505), .B(n9508), .Y(multiplier_i[11]) );
  CLKINVX1 U6961 ( .A(multiplier_r[15]), .Y(n9508) );
  NAND2X1 U6962 ( .A(n9157), .B(n9504), .Y(multiplier_r[15]) );
  OAI211X1 U6963 ( .A0(n6073), .A1(counter[0]), .B0(n9163), .C0(n9507), .Y(
        n9504) );
  CLKINVX1 U6964 ( .A(n9510), .Y(n9163) );
  NAND3X1 U6965 ( .A(n6075), .B(counter[2]), .C(n9507), .Y(n9157) );
  AND2X1 U6966 ( .A(n6072), .B(counter[1]), .Y(n9507) );
  CLKMX2X2 U6967 ( .A(n9511), .B(n9509), .S0(n6072), .Y(n9505) );
  OR2X1 U6968 ( .A(n9512), .B(n6073), .Y(n9509) );
  NAND2X1 U6969 ( .A(n9510), .B(counter[1]), .Y(n9511) );
  AOI21X1 U6970 ( .A0(n9513), .A1(n9514), .B0(data[15]), .Y(hd08_35) );
  XOR2X1 U6971 ( .A(n9515), .B(n9516), .Y(hd08_9_) );
  XOR2X1 U6972 ( .A(data[7]), .B(data[4]), .Y(n9516) );
  XNOR2X1 U6973 ( .A(n9517), .B(n9518), .Y(hd08_8_) );
  XNOR2X1 U6974 ( .A(data[6]), .B(n9519), .Y(n9518) );
  XOR2X1 U6975 ( .A(n9520), .B(n9521), .Y(hd08_7_) );
  XNOR2X1 U6976 ( .A(data[2]), .B(n9522), .Y(n9521) );
  XOR2X1 U6977 ( .A(n9523), .B(n9524), .Y(hd08_6_) );
  XNOR2X1 U6978 ( .A(data[1]), .B(data[4]), .Y(n9524) );
  OAI21XL U6979 ( .A0(data[0]), .A1(n9519), .B0(n9523), .Y(hd08_5_) );
  XOR2X1 U6980 ( .A(n9514), .B(n9525), .Y(hd08_20_) );
  XNOR2X1 U6981 ( .A(data[14]), .B(data[15]), .Y(n9525) );
  OAI21XL U6982 ( .A0(data[13]), .A1(n9526), .B0(n9513), .Y(n9514) );
  XOR2X1 U6983 ( .A(n9526), .B(n9527), .Y(hd08_19_) );
  XNOR2X1 U6984 ( .A(n9513), .B(data[13]), .Y(n9527) );
  OA21XL U6985 ( .A0(n9528), .A1(n9529), .B0(n9530), .Y(n9526) );
  AO21X1 U6986 ( .A0(n9529), .A1(n9528), .B0(data[15]), .Y(n9530) );
  XOR2X1 U6987 ( .A(n9528), .B(n9531), .Y(hd08_18_) );
  XNOR2X1 U6988 ( .A(data[15]), .B(n9529), .Y(n9531) );
  OA21XL U6989 ( .A0(data[12]), .A1(n9532), .B0(n9533), .Y(n9528) );
  OAI21XL U6990 ( .A0(n9534), .A1(n9535), .B0(data[15]), .Y(n9533) );
  XOR2X1 U6991 ( .A(n9532), .B(n9536), .Y(hd08_17_) );
  XNOR2X1 U6992 ( .A(data[15]), .B(n9534), .Y(n9536) );
  CLKINVX1 U6993 ( .A(n9535), .Y(n9532) );
  OAI22XL U6994 ( .A0(data[11]), .A1(n9537), .B0(n9538), .B1(n9513), .Y(n9535)
         );
  AND2X1 U6995 ( .A(data[11]), .B(n9537), .Y(n9538) );
  XOR2X1 U6996 ( .A(n9537), .B(n9539), .Y(hd08_16_) );
  XNOR2X1 U6997 ( .A(n9513), .B(data[11]), .Y(n9539) );
  CLKINVX1 U6998 ( .A(data[14]), .Y(n9513) );
  OA21XL U6999 ( .A0(data[10]), .A1(n9540), .B0(n9541), .Y(n9537) );
  OAI21XL U7000 ( .A0(n9542), .A1(n9543), .B0(data[13]), .Y(n9541) );
  XOR2X1 U7001 ( .A(n9540), .B(n9544), .Y(hd08_15_) );
  XNOR2X1 U7002 ( .A(n9529), .B(data[10]), .Y(n9544) );
  CLKINVX1 U7003 ( .A(data[13]), .Y(n9529) );
  CLKINVX1 U7004 ( .A(n9543), .Y(n9540) );
  OAI21XL U7005 ( .A0(n9545), .A1(n9534), .B0(n9546), .Y(n9543) );
  AO21X1 U7006 ( .A0(n9534), .A1(n9545), .B0(data[9]), .Y(n9546) );
  XOR2X1 U7007 ( .A(n9545), .B(n9547), .Y(hd08_14_) );
  XNOR2X1 U7008 ( .A(data[9]), .B(n9534), .Y(n9547) );
  CLKINVX1 U7009 ( .A(data[12]), .Y(n9534) );
  AOI2BB2X1 U7010 ( .B0(n9548), .B1(data[11]), .A0N(data[8]), .A1N(n9549), .Y(
        n9545) );
  NOR2X1 U7011 ( .A(data[11]), .B(n9548), .Y(n9549) );
  XNOR2X1 U7012 ( .A(n9548), .B(n9550), .Y(hd08_13_) );
  XOR2X1 U7013 ( .A(data[8]), .B(data[11]), .Y(n9550) );
  OAI21XL U7014 ( .A0(n9551), .A1(n9542), .B0(n9552), .Y(n9548) );
  AO21X1 U7015 ( .A0(n9542), .A1(n9551), .B0(data[7]), .Y(n9552) );
  XOR2X1 U7016 ( .A(n9551), .B(n9553), .Y(hd08_12_) );
  XNOR2X1 U7017 ( .A(data[7]), .B(n9542), .Y(n9553) );
  CLKINVX1 U7018 ( .A(data[10]), .Y(n9542) );
  OA21XL U7019 ( .A0(data[6]), .A1(n9554), .B0(n9555), .Y(n9551) );
  OAI2BB1X1 U7020 ( .A0N(data[6]), .A1N(n9554), .B0(data[9]), .Y(n9555) );
  XOR2X1 U7021 ( .A(n9554), .B(n9556), .Y(hd08_11_) );
  XOR2X1 U7022 ( .A(data[9]), .B(data[6]), .Y(n9556) );
  AOI22X1 U7023 ( .A0(n9522), .A1(n9557), .B0(n9558), .B1(data[8]), .Y(n9554)
         );
  OR2X1 U7024 ( .A(n9557), .B(n9522), .Y(n9558) );
  XNOR2X1 U7025 ( .A(n9557), .B(n9559), .Y(hd08_10_) );
  XNOR2X1 U7026 ( .A(data[8]), .B(n9522), .Y(n9559) );
  OAI21XL U7027 ( .A0(data[4]), .A1(n9515), .B0(n9560), .Y(n9557) );
  OAI2BB1X1 U7028 ( .A0N(data[4]), .A1N(n9515), .B0(data[7]), .Y(n9560) );
  AOI22X1 U7029 ( .A0(n9519), .A1(n9517), .B0(n9561), .B1(data[6]), .Y(n9515)
         );
  OR2X1 U7030 ( .A(n9517), .B(n9519), .Y(n9561) );
  OAI21XL U7031 ( .A0(n9520), .A1(n9522), .B0(n9562), .Y(n9517) );
  AO21X1 U7032 ( .A0(n9522), .A1(n9520), .B0(data[2]), .Y(n9562) );
  CLKINVX1 U7033 ( .A(data[5]), .Y(n9522) );
  AOI21X1 U7034 ( .A0(n9523), .A1(data[4]), .B0(n9563), .Y(n9520) );
  AOI2BB1X1 U7035 ( .A0N(data[4]), .A1N(n9523), .B0(data[1]), .Y(n9563) );
  NAND2X1 U7036 ( .A(data[0]), .B(n9519), .Y(n9523) );
  CLKINVX1 U7037 ( .A(data[3]), .Y(n9519) );
  CLKINVX1 U7038 ( .A(n9564), .Y(fir_d[9]) );
  CLKINVX1 U7039 ( .A(n9565), .Y(fir_d[8]) );
  CLKINVX1 U7040 ( .A(n9566), .Y(fir_d[7]) );
  CLKINVX1 U7041 ( .A(n9567), .Y(fir_d[6]) );
  CLKINVX1 U7042 ( .A(n9568), .Y(fir_d[5]) );
  CLKINVX1 U7043 ( .A(n9569), .Y(fir_d[4]) );
  CLKINVX1 U7044 ( .A(n9570), .Y(fir_d[3]) );
  CLKINVX1 U7045 ( .A(n9571), .Y(fir_d[2]) );
  CLKINVX1 U7046 ( .A(n9572), .Y(fir_d[1]) );
  CLKINVX1 U7047 ( .A(n9573), .Y(fir_d[15]) );
  CLKINVX1 U7048 ( .A(n9574), .Y(fir_d[14]) );
  CLKINVX1 U7049 ( .A(n9575), .Y(fir_d[13]) );
  CLKINVX1 U7050 ( .A(n9576), .Y(fir_d[12]) );
  CLKINVX1 U7051 ( .A(n9577), .Y(fir_d[11]) );
  CLKINVX1 U7052 ( .A(n9578), .Y(fir_d[10]) );
  CLKINVX1 U7053 ( .A(n9579), .Y(fir_d[0]) );
  OAI22XL U7054 ( .A0(n6166), .A1(n8781), .B0(n6134), .B1(n8794), .Y(U3_U8_Z_9) );
  OAI22XL U7055 ( .A0(n6167), .A1(n8781), .B0(n6135), .B1(n8794), .Y(U3_U8_Z_8) );
  OAI22XL U7056 ( .A0(n6168), .A1(n8781), .B0(n6136), .B1(n8794), .Y(U3_U8_Z_7) );
  OAI22XL U7057 ( .A0(n6169), .A1(n8781), .B0(n6137), .B1(n8794), .Y(U3_U8_Z_6) );
  OAI22XL U7058 ( .A0(n6170), .A1(n8781), .B0(n6138), .B1(n8794), .Y(U3_U8_Z_5) );
  OAI22XL U7059 ( .A0(n6171), .A1(n8781), .B0(n6139), .B1(n8794), .Y(U3_U8_Z_4) );
  OAI22XL U7060 ( .A0(n6144), .A1(n8781), .B0(n6112), .B1(n8794), .Y(
        U3_U8_Z_31) );
  OAI22XL U7061 ( .A0(n6145), .A1(n8781), .B0(n6113), .B1(n8794), .Y(
        U3_U8_Z_30) );
  OAI22XL U7062 ( .A0(n6172), .A1(n8781), .B0(n6140), .B1(n8794), .Y(U3_U8_Z_3) );
  OAI22XL U7063 ( .A0(n6146), .A1(n8781), .B0(n6114), .B1(n8794), .Y(
        U3_U8_Z_29) );
  OAI22XL U7064 ( .A0(n6147), .A1(n8781), .B0(n6115), .B1(n8794), .Y(
        U3_U8_Z_28) );
  OAI22XL U7065 ( .A0(n6148), .A1(n8781), .B0(n6116), .B1(n8794), .Y(
        U3_U8_Z_27) );
  OAI22XL U7066 ( .A0(n6149), .A1(n8782), .B0(n6117), .B1(n8794), .Y(
        U3_U8_Z_26) );
  OAI22XL U7067 ( .A0(n6150), .A1(n8782), .B0(n6118), .B1(n8794), .Y(
        U3_U8_Z_25) );
  OAI22XL U7068 ( .A0(n6151), .A1(n8782), .B0(n6119), .B1(n8794), .Y(
        U3_U8_Z_24) );
  OAI22XL U7069 ( .A0(n6152), .A1(n8782), .B0(n6120), .B1(n8794), .Y(
        U3_U8_Z_23) );
  OAI22XL U7070 ( .A0(n6153), .A1(n8782), .B0(n6121), .B1(n8794), .Y(
        U3_U8_Z_22) );
  OAI22XL U7071 ( .A0(n6154), .A1(n8782), .B0(n6122), .B1(n8794), .Y(
        U3_U8_Z_21) );
  OAI22XL U7072 ( .A0(n6155), .A1(n8782), .B0(n6123), .B1(n8794), .Y(
        U3_U8_Z_20) );
  OAI22XL U7073 ( .A0(n6173), .A1(n8782), .B0(n6141), .B1(n8795), .Y(U3_U8_Z_2) );
  OAI22XL U7074 ( .A0(n6156), .A1(n8782), .B0(n6124), .B1(n8795), .Y(
        U3_U8_Z_19) );
  OAI22XL U7075 ( .A0(n6157), .A1(n8782), .B0(n6125), .B1(n8795), .Y(
        U3_U8_Z_18) );
  OAI22XL U7076 ( .A0(n6158), .A1(n8782), .B0(n6126), .B1(n8795), .Y(
        U3_U8_Z_17) );
  OAI22XL U7077 ( .A0(n6159), .A1(n8782), .B0(n6127), .B1(n8795), .Y(
        U3_U8_Z_16) );
  OAI22XL U7078 ( .A0(n6160), .A1(n8782), .B0(n6128), .B1(n8795), .Y(
        U3_U8_Z_15) );
  OAI22XL U7079 ( .A0(n6161), .A1(n8782), .B0(n6129), .B1(n8795), .Y(
        U3_U8_Z_14) );
  OAI22XL U7080 ( .A0(n6162), .A1(n8782), .B0(n6130), .B1(n8795), .Y(
        U3_U8_Z_13) );
  OAI22XL U7081 ( .A0(n6163), .A1(n8782), .B0(n6131), .B1(n8795), .Y(
        U3_U8_Z_12) );
  OAI22XL U7082 ( .A0(n6164), .A1(n8783), .B0(n6132), .B1(n8796), .Y(
        U3_U8_Z_11) );
  OAI22XL U7083 ( .A0(n6165), .A1(n8782), .B0(n6133), .B1(n8795), .Y(
        U3_U8_Z_10) );
  OAI22XL U7084 ( .A0(n6174), .A1(n8782), .B0(n6142), .B1(n8795), .Y(U3_U8_Z_1) );
  OAI22XL U7085 ( .A0(n6175), .A1(n8782), .B0(n6143), .B1(n8795), .Y(U3_U8_Z_0) );
  OAI22XL U7086 ( .A0(n8788), .A1(n9408), .B0(n9335), .B1(n8795), .Y(U3_U7_Z_9) );
  OAI22XL U7087 ( .A0(n8787), .A1(n9406), .B0(n9333), .B1(n8795), .Y(U3_U7_Z_8) );
  OAI22XL U7088 ( .A0(n8787), .A1(n9404), .B0(n9331), .B1(n8795), .Y(U3_U7_Z_7) );
  OAI22XL U7089 ( .A0(n8787), .A1(n9402), .B0(n9329), .B1(n8795), .Y(U3_U7_Z_6) );
  OAI22XL U7090 ( .A0(n8787), .A1(n9400), .B0(n9327), .B1(n8795), .Y(U3_U7_Z_5) );
  OAI22XL U7091 ( .A0(n8787), .A1(n9398), .B0(n9325), .B1(n8795), .Y(U3_U7_Z_4) );
  OAI22XL U7092 ( .A0(n8787), .A1(n9389), .B0(n9379), .B1(n8795), .Y(
        U3_U7_Z_31) );
  OAI22XL U7093 ( .A0(n8787), .A1(n9463), .B0(n9377), .B1(n8795), .Y(
        U3_U7_Z_30) );
  OAI22XL U7094 ( .A0(n8787), .A1(n9396), .B0(n9323), .B1(n8796), .Y(U3_U7_Z_3) );
  OAI22XL U7095 ( .A0(n8787), .A1(n9460), .B0(n9375), .B1(n8796), .Y(
        U3_U7_Z_29) );
  OAI22XL U7096 ( .A0(n8786), .A1(n9457), .B0(n9373), .B1(n8796), .Y(
        U3_U7_Z_28) );
  OAI22XL U7097 ( .A0(n8786), .A1(n9454), .B0(n9371), .B1(n8796), .Y(
        U3_U7_Z_27) );
  OAI22XL U7098 ( .A0(n8787), .A1(n9451), .B0(n9369), .B1(n8796), .Y(
        U3_U7_Z_26) );
  OAI22XL U7099 ( .A0(n8787), .A1(n9448), .B0(n9367), .B1(n8796), .Y(
        U3_U7_Z_25) );
  OAI22XL U7100 ( .A0(n8786), .A1(n9445), .B0(n9365), .B1(n8796), .Y(
        U3_U7_Z_24) );
  OAI22XL U7101 ( .A0(n8787), .A1(n9442), .B0(n9363), .B1(n8796), .Y(
        U3_U7_Z_23) );
  OAI22XL U7102 ( .A0(n8786), .A1(n9439), .B0(n9361), .B1(n8796), .Y(
        U3_U7_Z_22) );
  OAI22XL U7103 ( .A0(n8786), .A1(n9436), .B0(n9359), .B1(n8796), .Y(
        U3_U7_Z_21) );
  OAI22XL U7104 ( .A0(n8787), .A1(n9433), .B0(n9357), .B1(n8796), .Y(
        U3_U7_Z_20) );
  OAI22XL U7105 ( .A0(n8786), .A1(n9394), .B0(n9321), .B1(n8796), .Y(U3_U7_Z_2) );
  OAI22XL U7106 ( .A0(n8787), .A1(n9430), .B0(n9355), .B1(n8796), .Y(
        U3_U7_Z_19) );
  OAI22XL U7107 ( .A0(n8787), .A1(n9427), .B0(n9353), .B1(n8796), .Y(
        U3_U7_Z_18) );
  OAI22XL U7108 ( .A0(n8786), .A1(n9424), .B0(n9351), .B1(n8796), .Y(
        U3_U7_Z_17) );
  OAI22XL U7109 ( .A0(n8786), .A1(n9386), .B0(n9349), .B1(n8796), .Y(
        U3_U7_Z_16) );
  OAI22XL U7110 ( .A0(n8787), .A1(n9420), .B0(n9347), .B1(n8796), .Y(
        U3_U7_Z_15) );
  OAI22XL U7111 ( .A0(n8786), .A1(n9418), .B0(n9345), .B1(n8796), .Y(
        U3_U7_Z_14) );
  OAI22XL U7112 ( .A0(n8786), .A1(n9416), .B0(n9343), .B1(n8796), .Y(
        U3_U7_Z_13) );
  OAI22XL U7113 ( .A0(n8787), .A1(n9414), .B0(n9341), .B1(n8797), .Y(
        U3_U7_Z_12) );
  OAI22XL U7114 ( .A0(n8787), .A1(n9412), .B0(n9339), .B1(n8797), .Y(
        U3_U7_Z_11) );
  OAI22XL U7115 ( .A0(n8786), .A1(n9410), .B0(n9337), .B1(n8797), .Y(
        U3_U7_Z_10) );
  OAI22XL U7116 ( .A0(n8787), .A1(n9392), .B0(n9319), .B1(n8797), .Y(U3_U7_Z_1) );
  OAI22XL U7117 ( .A0(n8786), .A1(n9390), .B0(n9316), .B1(n8797), .Y(U3_U7_Z_0) );
  OAI22XL U7118 ( .A0(n6134), .A1(n8783), .B0(n6166), .B1(n8797), .Y(U3_U6_Z_9) );
  OAI22XL U7119 ( .A0(n6135), .A1(n8783), .B0(n6167), .B1(n8797), .Y(U3_U6_Z_8) );
  OAI22XL U7120 ( .A0(n6136), .A1(n8783), .B0(n6168), .B1(n8797), .Y(U3_U6_Z_7) );
  OAI22XL U7121 ( .A0(n6137), .A1(n8783), .B0(n6169), .B1(n8797), .Y(U3_U6_Z_6) );
  OAI22XL U7122 ( .A0(n6138), .A1(n8783), .B0(n6170), .B1(n8797), .Y(U3_U6_Z_5) );
  OAI22XL U7123 ( .A0(n6139), .A1(n8783), .B0(n6171), .B1(n8797), .Y(U3_U6_Z_4) );
  OAI22XL U7124 ( .A0(n6112), .A1(n8783), .B0(n6144), .B1(n8797), .Y(
        U3_U6_Z_31) );
  OAI22XL U7125 ( .A0(n6113), .A1(n8783), .B0(n6145), .B1(n8797), .Y(
        U3_U6_Z_30) );
  OAI22XL U7126 ( .A0(n6140), .A1(n8783), .B0(n6172), .B1(n8797), .Y(U3_U6_Z_3) );
  OAI22XL U7127 ( .A0(n6114), .A1(n8783), .B0(n6146), .B1(n8797), .Y(
        U3_U6_Z_29) );
  OAI22XL U7128 ( .A0(n6115), .A1(n8783), .B0(n6147), .B1(n8797), .Y(
        U3_U6_Z_28) );
  OAI22XL U7129 ( .A0(n6116), .A1(n8783), .B0(n6148), .B1(n8797), .Y(
        U3_U6_Z_27) );
  OAI22XL U7130 ( .A0(n6117), .A1(n8783), .B0(n6149), .B1(n8797), .Y(
        U3_U6_Z_26) );
  OAI22XL U7131 ( .A0(n6118), .A1(n8783), .B0(n6150), .B1(n8797), .Y(
        U3_U6_Z_25) );
  OAI22XL U7132 ( .A0(n6119), .A1(n8783), .B0(n6151), .B1(n8797), .Y(
        U3_U6_Z_24) );
  OAI22XL U7133 ( .A0(n6120), .A1(n8783), .B0(n6152), .B1(n8798), .Y(
        U3_U6_Z_23) );
  OAI22XL U7134 ( .A0(n6121), .A1(n8783), .B0(n6153), .B1(n8798), .Y(
        U3_U6_Z_22) );
  OAI22XL U7135 ( .A0(n6122), .A1(n8783), .B0(n6154), .B1(n8798), .Y(
        U3_U6_Z_21) );
  OAI22XL U7136 ( .A0(n6123), .A1(n8784), .B0(n6155), .B1(n8798), .Y(
        U3_U6_Z_20) );
  OAI22XL U7137 ( .A0(n6141), .A1(n8784), .B0(n6173), .B1(n8798), .Y(U3_U6_Z_2) );
  OAI22XL U7138 ( .A0(n6124), .A1(n8784), .B0(n6156), .B1(n8798), .Y(
        U3_U6_Z_19) );
  OAI22XL U7139 ( .A0(n6125), .A1(n8784), .B0(n6157), .B1(n8798), .Y(
        U3_U6_Z_18) );
  OAI22XL U7140 ( .A0(n6126), .A1(n8784), .B0(n6158), .B1(n8798), .Y(
        U3_U6_Z_17) );
  OAI22XL U7141 ( .A0(n6127), .A1(n8784), .B0(n6159), .B1(n8798), .Y(
        U3_U6_Z_16) );
  OAI22XL U7142 ( .A0(n6128), .A1(n8784), .B0(n6160), .B1(n8798), .Y(
        U3_U6_Z_15) );
  OAI22XL U7143 ( .A0(n6129), .A1(n8784), .B0(n6161), .B1(n8798), .Y(
        U3_U6_Z_14) );
  OAI22XL U7144 ( .A0(n6130), .A1(n8784), .B0(n6162), .B1(n8798), .Y(
        U3_U6_Z_13) );
  OAI22XL U7145 ( .A0(n6131), .A1(n8784), .B0(n6163), .B1(n8798), .Y(
        U3_U6_Z_12) );
  OAI22XL U7146 ( .A0(n6132), .A1(n8785), .B0(n6164), .B1(n8798), .Y(
        U3_U6_Z_11) );
  OAI22XL U7147 ( .A0(n6133), .A1(n8784), .B0(n6165), .B1(n8798), .Y(
        U3_U6_Z_10) );
  OAI22XL U7148 ( .A0(n6142), .A1(n8784), .B0(n6174), .B1(n8798), .Y(U3_U6_Z_1) );
  OAI22XL U7149 ( .A0(n6143), .A1(n8785), .B0(n6175), .B1(n8794), .Y(U3_U6_Z_0) );
  OAI22XL U7150 ( .A0(n9335), .A1(n8784), .B0(n8793), .B1(n9408), .Y(U3_U5_Z_9) );
  CLKINVX1 U7151 ( .A(BF2I_b_ei_n[9]), .Y(n9408) );
  CLKINVX1 U7152 ( .A(BF2I_b_er_n[9]), .Y(n9335) );
  OAI22XL U7153 ( .A0(n9333), .A1(n8785), .B0(n8793), .B1(n9406), .Y(U3_U5_Z_8) );
  CLKINVX1 U7154 ( .A(BF2I_b_ei_n[8]), .Y(n9406) );
  CLKINVX1 U7155 ( .A(BF2I_b_er_n[8]), .Y(n9333) );
  OAI22XL U7156 ( .A0(n9331), .A1(n8784), .B0(n8793), .B1(n9404), .Y(U3_U5_Z_7) );
  CLKINVX1 U7157 ( .A(BF2I_b_ei_n[7]), .Y(n9404) );
  CLKINVX1 U7158 ( .A(BF2I_b_er_n[7]), .Y(n9331) );
  OAI22XL U7159 ( .A0(n9329), .A1(n8784), .B0(n8793), .B1(n9402), .Y(U3_U5_Z_6) );
  CLKINVX1 U7160 ( .A(BF2I_b_ei_n[6]), .Y(n9402) );
  CLKINVX1 U7161 ( .A(BF2I_b_er_n[6]), .Y(n9329) );
  OAI22XL U7162 ( .A0(n9327), .A1(n8785), .B0(n8793), .B1(n9400), .Y(U3_U5_Z_5) );
  CLKINVX1 U7163 ( .A(BF2I_b_ei_n[5]), .Y(n9400) );
  CLKINVX1 U7164 ( .A(BF2I_b_er_n[5]), .Y(n9327) );
  OAI22XL U7165 ( .A0(n9325), .A1(n8785), .B0(n8793), .B1(n9398), .Y(U3_U5_Z_4) );
  CLKINVX1 U7166 ( .A(BF2I_b_ei_n[4]), .Y(n9398) );
  CLKINVX1 U7167 ( .A(BF2I_b_er_n[4]), .Y(n9325) );
  OAI22XL U7168 ( .A0(n9379), .A1(n8785), .B0(n8793), .B1(n9389), .Y(
        U3_U5_Z_31) );
  CLKINVX1 U7169 ( .A(BF2I_b_ei_n[31]), .Y(n9389) );
  CLKINVX1 U7170 ( .A(BF2I_b_er_n[31]), .Y(n9379) );
  OAI22XL U7171 ( .A0(n9377), .A1(n8785), .B0(n8793), .B1(n9463), .Y(
        U3_U5_Z_30) );
  CLKINVX1 U7172 ( .A(BF2I_b_ei_n[30]), .Y(n9463) );
  CLKINVX1 U7173 ( .A(BF2I_b_er_n[30]), .Y(n9377) );
  OAI22XL U7174 ( .A0(n9323), .A1(n8785), .B0(n8793), .B1(n9396), .Y(U3_U5_Z_3) );
  CLKINVX1 U7175 ( .A(BF2I_b_ei_n[3]), .Y(n9396) );
  CLKINVX1 U7176 ( .A(BF2I_b_er_n[3]), .Y(n9323) );
  OAI22XL U7177 ( .A0(n9375), .A1(n8784), .B0(n8793), .B1(n9460), .Y(
        U3_U5_Z_29) );
  CLKINVX1 U7178 ( .A(BF2I_b_ei_n[29]), .Y(n9460) );
  CLKINVX1 U7179 ( .A(BF2I_b_er_n[29]), .Y(n9375) );
  OAI22XL U7180 ( .A0(n9373), .A1(n8785), .B0(n8793), .B1(n9457), .Y(
        U3_U5_Z_28) );
  CLKINVX1 U7181 ( .A(BF2I_b_ei_n[28]), .Y(n9457) );
  CLKINVX1 U7182 ( .A(BF2I_b_er_n[28]), .Y(n9373) );
  OAI22XL U7183 ( .A0(n9371), .A1(n8785), .B0(n8793), .B1(n9454), .Y(
        U3_U5_Z_27) );
  CLKINVX1 U7184 ( .A(BF2I_b_ei_n[27]), .Y(n9454) );
  CLKINVX1 U7185 ( .A(BF2I_b_er_n[27]), .Y(n9371) );
  OAI22XL U7186 ( .A0(n9369), .A1(n8785), .B0(n8793), .B1(n9451), .Y(
        U3_U5_Z_26) );
  CLKINVX1 U7187 ( .A(BF2I_b_ei_n[26]), .Y(n9451) );
  CLKINVX1 U7188 ( .A(BF2I_b_er_n[26]), .Y(n9369) );
  OAI22XL U7189 ( .A0(n9367), .A1(n8785), .B0(n8793), .B1(n9448), .Y(
        U3_U5_Z_25) );
  CLKINVX1 U7190 ( .A(BF2I_b_ei_n[25]), .Y(n9448) );
  CLKINVX1 U7191 ( .A(BF2I_b_er_n[25]), .Y(n9367) );
  OAI22XL U7192 ( .A0(n9365), .A1(n8784), .B0(n8793), .B1(n9445), .Y(
        U3_U5_Z_24) );
  CLKINVX1 U7193 ( .A(BF2I_b_ei_n[24]), .Y(n9445) );
  CLKINVX1 U7194 ( .A(BF2I_b_er_n[24]), .Y(n9365) );
  OAI22XL U7195 ( .A0(n9363), .A1(n8785), .B0(n8793), .B1(n9442), .Y(
        U3_U5_Z_23) );
  CLKINVX1 U7196 ( .A(BF2I_b_ei_n[23]), .Y(n9442) );
  CLKINVX1 U7197 ( .A(BF2I_b_er_n[23]), .Y(n9363) );
  OAI22XL U7198 ( .A0(n9361), .A1(n8784), .B0(n8793), .B1(n9439), .Y(
        U3_U5_Z_22) );
  CLKINVX1 U7199 ( .A(BF2I_b_ei_n[22]), .Y(n9439) );
  CLKINVX1 U7200 ( .A(BF2I_b_er_n[22]), .Y(n9361) );
  OAI22XL U7201 ( .A0(n9359), .A1(n8785), .B0(n8793), .B1(n9436), .Y(
        U3_U5_Z_21) );
  CLKINVX1 U7202 ( .A(BF2I_b_ei_n[21]), .Y(n9436) );
  CLKINVX1 U7203 ( .A(BF2I_b_er_n[21]), .Y(n9359) );
  OAI22XL U7204 ( .A0(n9357), .A1(n8785), .B0(n8792), .B1(n9433), .Y(
        U3_U5_Z_20) );
  CLKINVX1 U7205 ( .A(BF2I_b_ei_n[20]), .Y(n9433) );
  CLKINVX1 U7206 ( .A(BF2I_b_er_n[20]), .Y(n9357) );
  OAI22XL U7207 ( .A0(n9321), .A1(n8786), .B0(n8792), .B1(n9394), .Y(U3_U5_Z_2) );
  CLKINVX1 U7208 ( .A(BF2I_b_ei_n[2]), .Y(n9394) );
  CLKINVX1 U7209 ( .A(BF2I_b_er_n[2]), .Y(n9321) );
  OAI22XL U7210 ( .A0(n9355), .A1(n8786), .B0(n8792), .B1(n9430), .Y(
        U3_U5_Z_19) );
  CLKINVX1 U7211 ( .A(BF2I_b_ei_n[19]), .Y(n9430) );
  CLKINVX1 U7212 ( .A(BF2I_b_er_n[19]), .Y(n9355) );
  OAI22XL U7213 ( .A0(n9353), .A1(n8785), .B0(n8792), .B1(n9427), .Y(
        U3_U5_Z_18) );
  CLKINVX1 U7214 ( .A(BF2I_b_ei_n[18]), .Y(n9427) );
  CLKINVX1 U7215 ( .A(BF2I_b_er_n[18]), .Y(n9353) );
  OAI22XL U7216 ( .A0(n9351), .A1(n8786), .B0(n8792), .B1(n9424), .Y(
        U3_U5_Z_17) );
  CLKINVX1 U7217 ( .A(BF2I_b_ei_n[17]), .Y(n9424) );
  CLKINVX1 U7218 ( .A(BF2I_b_er_n[17]), .Y(n9351) );
  OAI22XL U7219 ( .A0(n9349), .A1(n8785), .B0(n8792), .B1(n9386), .Y(
        U3_U5_Z_16) );
  CLKINVX1 U7220 ( .A(BF2I_b_ei_n[16]), .Y(n9386) );
  CLKINVX1 U7221 ( .A(BF2I_b_er_n[16]), .Y(n9349) );
  OAI22XL U7222 ( .A0(n9347), .A1(n8785), .B0(n8792), .B1(n9420), .Y(
        U3_U5_Z_15) );
  CLKINVX1 U7223 ( .A(BF2I_b_ei_n[15]), .Y(n9420) );
  CLKINVX1 U7224 ( .A(BF2I_b_er_n[15]), .Y(n9347) );
  OAI22XL U7225 ( .A0(n9345), .A1(n8786), .B0(n8792), .B1(n9418), .Y(
        U3_U5_Z_14) );
  CLKINVX1 U7226 ( .A(BF2I_b_ei_n[14]), .Y(n9418) );
  CLKINVX1 U7227 ( .A(BF2I_b_er_n[14]), .Y(n9345) );
  OAI22XL U7228 ( .A0(n9343), .A1(n8786), .B0(n8792), .B1(n9416), .Y(
        U3_U5_Z_13) );
  CLKINVX1 U7229 ( .A(BF2I_b_ei_n[13]), .Y(n9416) );
  CLKINVX1 U7230 ( .A(BF2I_b_er_n[13]), .Y(n9343) );
  OAI22XL U7231 ( .A0(n9341), .A1(n8785), .B0(n8792), .B1(n9414), .Y(
        U3_U5_Z_12) );
  CLKINVX1 U7232 ( .A(BF2I_b_ei_n[12]), .Y(n9414) );
  CLKINVX1 U7233 ( .A(BF2I_b_er_n[12]), .Y(n9341) );
  OAI22XL U7234 ( .A0(n9339), .A1(n8786), .B0(n8792), .B1(n9412), .Y(
        U3_U5_Z_11) );
  CLKINVX1 U7235 ( .A(BF2I_b_ei_n[11]), .Y(n9412) );
  CLKINVX1 U7236 ( .A(BF2I_b_er_n[11]), .Y(n9339) );
  OAI22XL U7237 ( .A0(n9337), .A1(n8786), .B0(n8792), .B1(n9410), .Y(
        U3_U5_Z_10) );
  CLKINVX1 U7238 ( .A(BF2I_b_ei_n[10]), .Y(n9410) );
  CLKINVX1 U7239 ( .A(BF2I_b_er_n[10]), .Y(n9337) );
  OAI22XL U7240 ( .A0(n9319), .A1(n8784), .B0(n8793), .B1(n9392), .Y(U3_U5_Z_1) );
  CLKINVX1 U7241 ( .A(BF2I_b_ei_n[1]), .Y(n9392) );
  CLKINVX1 U7242 ( .A(BF2I_b_er_n[1]), .Y(n9319) );
  OAI22XL U7243 ( .A0(n9316), .A1(n8781), .B0(n8792), .B1(n9390), .Y(U3_U5_Z_0) );
  CLKINVX1 U7244 ( .A(BF2I_b_ei_n[0]), .Y(n9390) );
  CLKINVX1 U7245 ( .A(n9381), .Y(n9465) );
  NOR2X1 U7246 ( .A(BF2I_b_s), .B(n10473), .Y(n9381) );
  CLKINVX1 U7247 ( .A(n9380), .Y(n9464) );
  NOR2X1 U7248 ( .A(n10473), .B(n6111), .Y(n9380) );
  CLKINVX1 U7249 ( .A(BF2I_b_er_n[0]), .Y(n9316) );
  OAI22XL U7250 ( .A0(n6101), .A1(n9245), .B0(n6085), .B1(n9246), .Y(U3_U3_Z_9) );
  OAI22XL U7251 ( .A0(n6102), .A1(n9245), .B0(n6086), .B1(n9246), .Y(U3_U3_Z_8) );
  OAI22XL U7252 ( .A0(n6103), .A1(n9245), .B0(n6087), .B1(n9246), .Y(U3_U3_Z_7) );
  OAI22XL U7253 ( .A0(n6104), .A1(n9245), .B0(n6088), .B1(n9246), .Y(U3_U3_Z_6) );
  OAI22XL U7254 ( .A0(n6105), .A1(n9245), .B0(n6089), .B1(n9246), .Y(U3_U3_Z_5) );
  OAI22XL U7255 ( .A0(n6106), .A1(n9245), .B0(n6090), .B1(n9246), .Y(U3_U3_Z_4) );
  OAI22XL U7256 ( .A0(n6107), .A1(n9245), .B0(n6091), .B1(n9246), .Y(U3_U3_Z_3) );
  OAI22XL U7257 ( .A0(n6108), .A1(n9245), .B0(n6092), .B1(n9246), .Y(U3_U3_Z_2) );
  OAI22XL U7258 ( .A0(n6095), .A1(n9245), .B0(n6079), .B1(n9246), .Y(
        U3_U3_Z_15) );
  OAI22XL U7259 ( .A0(n6096), .A1(n9245), .B0(n6080), .B1(n9246), .Y(
        U3_U3_Z_14) );
  OAI22XL U7260 ( .A0(n6097), .A1(n9245), .B0(n6081), .B1(n9246), .Y(
        U3_U3_Z_13) );
  OAI22XL U7261 ( .A0(n6098), .A1(n9245), .B0(n6082), .B1(n9246), .Y(
        U3_U3_Z_12) );
  OAI22XL U7262 ( .A0(n6099), .A1(n9245), .B0(n6083), .B1(n9246), .Y(
        U3_U3_Z_11) );
  OAI22XL U7263 ( .A0(n6100), .A1(n9245), .B0(n6084), .B1(n9246), .Y(
        U3_U3_Z_10) );
  OAI22XL U7264 ( .A0(n6109), .A1(n9245), .B0(n6093), .B1(n9246), .Y(U3_U3_Z_1) );
  OAI22XL U7265 ( .A0(n6110), .A1(n9245), .B0(n6094), .B1(n9246), .Y(U3_U3_Z_0) );
  NOR2X1 U7266 ( .A(n10052), .B(n8889), .Y(N999) );
  NOR2X1 U7267 ( .A(n10051), .B(n8889), .Y(N998) );
  NOR2X1 U7268 ( .A(n10050), .B(n8889), .Y(N997) );
  NOR2X1 U7269 ( .A(n10049), .B(n8889), .Y(N996) );
  NOR2X1 U7270 ( .A(n10048), .B(n8889), .Y(N995) );
  NOR2X1 U7271 ( .A(n10047), .B(n8888), .Y(N994) );
  NOR2X1 U7272 ( .A(n10046), .B(n8888), .Y(N993) );
  NOR2X1 U7273 ( .A(n10045), .B(n8888), .Y(N992) );
  NOR2X1 U7274 ( .A(n10044), .B(n8888), .Y(N991) );
  NOR2X1 U7275 ( .A(n10043), .B(n8888), .Y(N990) );
  NOR2X1 U7276 ( .A(n10042), .B(n8888), .Y(N989) );
  NOR2X1 U7277 ( .A(n10041), .B(n8888), .Y(N988) );
  NOR2X1 U7278 ( .A(n10040), .B(n8888), .Y(N987) );
  NOR2X1 U7279 ( .A(n10039), .B(n8888), .Y(N986) );
  NOR2X1 U7280 ( .A(n10038), .B(n8888), .Y(N985) );
  NOR2X1 U7281 ( .A(n9813), .B(n8888), .Y(N984) );
  NOR2X1 U7282 ( .A(n9812), .B(n8888), .Y(N983) );
  NOR2X1 U7283 ( .A(n9811), .B(n8888), .Y(N982) );
  NOR2X1 U7284 ( .A(n9810), .B(n8887), .Y(N981) );
  NOR2X1 U7285 ( .A(n9809), .B(n8887), .Y(N980) );
  NOR2X1 U7286 ( .A(n9808), .B(n8887), .Y(N979) );
  NOR2X1 U7287 ( .A(n9807), .B(n8887), .Y(N978) );
  NOR2X1 U7288 ( .A(n9806), .B(n8887), .Y(N977) );
  NOR2X1 U7289 ( .A(n9805), .B(n8887), .Y(N976) );
  NOR2X1 U7290 ( .A(n9804), .B(n8887), .Y(N975) );
  NOR2X1 U7291 ( .A(n9803), .B(n8887), .Y(N974) );
  NOR2X1 U7292 ( .A(n9802), .B(n8887), .Y(N973) );
  NOR2X1 U7293 ( .A(n9801), .B(n8887), .Y(N972) );
  NOR2X1 U7294 ( .A(n9800), .B(n8887), .Y(N971) );
  NOR2X1 U7295 ( .A(n9799), .B(n8887), .Y(N970) );
  NOR2X1 U7296 ( .A(n9798), .B(n8887), .Y(N969) );
  NOR2X1 U7297 ( .A(n9797), .B(n8886), .Y(N968) );
  NOR2X1 U7298 ( .A(n9796), .B(n8886), .Y(N967) );
  NOR2X1 U7299 ( .A(n9795), .B(n8886), .Y(N966) );
  NOR2X1 U7300 ( .A(n9794), .B(n8886), .Y(N965) );
  NOR2X1 U7301 ( .A(n9793), .B(n8886), .Y(N964) );
  NOR2X1 U7302 ( .A(n9792), .B(n8886), .Y(N963) );
  NOR2X1 U7303 ( .A(n9791), .B(n8886), .Y(N962) );
  NOR2X1 U7304 ( .A(n9790), .B(n8886), .Y(N961) );
  NOR2X1 U7305 ( .A(n9789), .B(n8886), .Y(N960) );
  NOR2X1 U7306 ( .A(n9788), .B(n8886), .Y(N959) );
  NOR2X1 U7307 ( .A(n9787), .B(n8886), .Y(N958) );
  NOR2X1 U7308 ( .A(n9786), .B(n8886), .Y(N957) );
  NOR2X1 U7309 ( .A(n9785), .B(n8886), .Y(N956) );
  NOR2X1 U7310 ( .A(n9784), .B(n8885), .Y(N955) );
  NOR2X1 U7311 ( .A(n9783), .B(n8885), .Y(N954) );
  NOR2X1 U7312 ( .A(n9782), .B(n8885), .Y(N953) );
  NOR2X1 U7313 ( .A(n10133), .B(n8885), .Y(N952) );
  NOR2X1 U7314 ( .A(n10132), .B(n8885), .Y(N951) );
  NOR2X1 U7315 ( .A(n10131), .B(n8885), .Y(N950) );
  NOR2X1 U7316 ( .A(n10130), .B(n8885), .Y(N949) );
  NOR2X1 U7317 ( .A(n10129), .B(n8885), .Y(N948) );
  NOR2X1 U7318 ( .A(n10128), .B(n8885), .Y(N947) );
  NOR2X1 U7319 ( .A(n10127), .B(n8885), .Y(N946) );
  NOR2X1 U7320 ( .A(n10126), .B(n8885), .Y(N945) );
  NOR2X1 U7321 ( .A(n10125), .B(n8885), .Y(N944) );
  NOR2X1 U7322 ( .A(n10124), .B(n8885), .Y(N943) );
  NOR2X1 U7323 ( .A(n10123), .B(n8884), .Y(N942) );
  NOR2X1 U7324 ( .A(n10122), .B(n8884), .Y(N941) );
  NOR2X1 U7325 ( .A(n10121), .B(n8884), .Y(N940) );
  NOR2X1 U7326 ( .A(n10120), .B(n8884), .Y(N939) );
  NOR2X1 U7327 ( .A(n10119), .B(n8884), .Y(N938) );
  NOR2X1 U7328 ( .A(n10118), .B(n8884), .Y(N937) );
  NOR2X1 U7329 ( .A(n10117), .B(n8884), .Y(N936) );
  NOR2X1 U7330 ( .A(n10116), .B(n8884), .Y(N935) );
  NOR2X1 U7331 ( .A(n10115), .B(n8884), .Y(N934) );
  NOR2X1 U7332 ( .A(n10114), .B(n8884), .Y(N933) );
  NOR2X1 U7333 ( .A(n10113), .B(n8884), .Y(N932) );
  NOR2X1 U7334 ( .A(n10112), .B(n8884), .Y(N931) );
  NOR2X1 U7335 ( .A(n10111), .B(n8884), .Y(N930) );
  NOR2X1 U7336 ( .A(n101101), .B(n8883), .Y(N929) );
  NOR2X1 U7337 ( .A(n10109), .B(n8883), .Y(N928) );
  NOR2X1 U7338 ( .A(n10108), .B(n8883), .Y(N927) );
  NOR2X1 U7339 ( .A(n10107), .B(n8883), .Y(N926) );
  NOR2X1 U7340 ( .A(n10106), .B(n8883), .Y(N925) );
  NOR2X1 U7341 ( .A(n10105), .B(n8883), .Y(N924) );
  NOR2X1 U7342 ( .A(n10104), .B(n8883), .Y(N923) );
  NOR2X1 U7343 ( .A(n10103), .B(n8883), .Y(N922) );
  NOR2X1 U7344 ( .A(n10102), .B(n8883), .Y(N921) );
  NOR2X1 U7345 ( .A(n9877), .B(n8883), .Y(N920) );
  NOR2X1 U7346 ( .A(n9876), .B(n8883), .Y(N919) );
  NOR2X1 U7347 ( .A(n9875), .B(n8883), .Y(N918) );
  NOR2X1 U7348 ( .A(n9874), .B(n8883), .Y(N917) );
  NOR2X1 U7349 ( .A(n9873), .B(n8882), .Y(N916) );
  NOR2X1 U7350 ( .A(n9872), .B(n8882), .Y(N915) );
  NOR2X1 U7351 ( .A(n9871), .B(n8882), .Y(N914) );
  NOR2X1 U7352 ( .A(n9870), .B(n8882), .Y(N913) );
  NOR2X1 U7353 ( .A(n9869), .B(n8882), .Y(N912) );
  NOR2X1 U7354 ( .A(n9868), .B(n8882), .Y(N911) );
  NOR2X1 U7355 ( .A(n9867), .B(n8882), .Y(N910) );
  NOR2X1 U7356 ( .A(n9866), .B(n8882), .Y(N909) );
  NOR2X1 U7357 ( .A(n9865), .B(n8882), .Y(N908) );
  NOR2X1 U7358 ( .A(n9864), .B(n8882), .Y(N907) );
  NOR2X1 U7359 ( .A(n9863), .B(n8882), .Y(N906) );
  NOR2X1 U7360 ( .A(n9862), .B(n8882), .Y(N905) );
  NOR2X1 U7361 ( .A(n9861), .B(n8882), .Y(N904) );
  NOR2X1 U7362 ( .A(n9860), .B(n8881), .Y(N903) );
  NOR2X1 U7363 ( .A(n9859), .B(n8881), .Y(N902) );
  NOR2X1 U7364 ( .A(n9858), .B(n8881), .Y(N901) );
  NOR2X1 U7365 ( .A(n9857), .B(n8881), .Y(N900) );
  NOR2X1 U7366 ( .A(n9856), .B(n8881), .Y(N899) );
  NOR2X1 U7367 ( .A(n9855), .B(n8881), .Y(N898) );
  NOR2X1 U7368 ( .A(n9854), .B(n8881), .Y(N897) );
  NOR2X1 U7369 ( .A(n9853), .B(n8881), .Y(N896) );
  NOR2X1 U7370 ( .A(n9852), .B(n8881), .Y(N895) );
  NOR2X1 U7371 ( .A(n9851), .B(n8881), .Y(N894) );
  NOR2X1 U7372 ( .A(n9850), .B(n8881), .Y(N893) );
  NOR2X1 U7373 ( .A(n9849), .B(n8881), .Y(N892) );
  NOR2X1 U7374 ( .A(n9848), .B(n8881), .Y(N891) );
  NOR2X1 U7375 ( .A(n9847), .B(n8880), .Y(N890) );
  NOR2X1 U7376 ( .A(n9846), .B(n8880), .Y(N889) );
  NOR2X1 U7377 ( .A(n10005), .B(n8880), .Y(N888) );
  NOR2X1 U7378 ( .A(n10004), .B(n8880), .Y(N887) );
  NOR2X1 U7379 ( .A(n10003), .B(n8880), .Y(N886) );
  NOR2X1 U7380 ( .A(n10002), .B(n8880), .Y(N885) );
  NOR2X1 U7381 ( .A(n10001), .B(n8880), .Y(N884) );
  NOR2X1 U7382 ( .A(n10000), .B(n8880), .Y(N883) );
  NOR2X1 U7383 ( .A(n9999), .B(n8880), .Y(N882) );
  NOR2X1 U7384 ( .A(n9998), .B(n8880), .Y(N881) );
  NOR2X1 U7385 ( .A(n9997), .B(n8880), .Y(N880) );
  NOR2X1 U7386 ( .A(n9996), .B(n8880), .Y(N879) );
  NOR2X1 U7387 ( .A(n9995), .B(n8880), .Y(N878) );
  NOR2X1 U7388 ( .A(n9994), .B(n8879), .Y(N877) );
  NOR2X1 U7389 ( .A(n9993), .B(n8879), .Y(N876) );
  NOR2X1 U7390 ( .A(n9992), .B(n8879), .Y(N875) );
  NOR2X1 U7391 ( .A(n9991), .B(n8879), .Y(N874) );
  NOR2X1 U7392 ( .A(n9990), .B(n8879), .Y(N873) );
  NOR2X1 U7393 ( .A(n9989), .B(n8879), .Y(N872) );
  NOR2X1 U7394 ( .A(n9988), .B(n8879), .Y(N871) );
  NOR2X1 U7395 ( .A(n9987), .B(n8879), .Y(N870) );
  NOR2X1 U7396 ( .A(n9986), .B(n8879), .Y(N869) );
  NOR2X1 U7397 ( .A(n9985), .B(n8879), .Y(N868) );
  NOR2X1 U7398 ( .A(n9984), .B(n8879), .Y(N867) );
  NOR2X1 U7399 ( .A(n9983), .B(n8879), .Y(N866) );
  NOR2X1 U7400 ( .A(n9982), .B(n8879), .Y(N865) );
  NOR2X1 U7401 ( .A(n9981), .B(n8878), .Y(N864) );
  NOR2X1 U7402 ( .A(n9980), .B(n8878), .Y(N863) );
  NOR2X1 U7403 ( .A(n9979), .B(n8878), .Y(N862) );
  NOR2X1 U7404 ( .A(n9978), .B(n8878), .Y(N861) );
  NOR2X1 U7405 ( .A(n9977), .B(n8878), .Y(N860) );
  NOR2X1 U7406 ( .A(n9976), .B(n8878), .Y(N859) );
  NOR2X1 U7407 ( .A(n9975), .B(n8878), .Y(N858) );
  NOR2X1 U7408 ( .A(n9974), .B(n8878), .Y(N857) );
  NOR2X1 U7409 ( .A(n9749), .B(n8878), .Y(N856) );
  NOR2X1 U7410 ( .A(n9748), .B(n8878), .Y(N855) );
  NOR2X1 U7411 ( .A(n9747), .B(n8878), .Y(N854) );
  NOR2X1 U7412 ( .A(n9746), .B(n8878), .Y(N853) );
  NOR2X1 U7413 ( .A(n9745), .B(n8878), .Y(N852) );
  NOR2X1 U7414 ( .A(n9744), .B(n8877), .Y(N851) );
  NOR2X1 U7415 ( .A(n9743), .B(n8877), .Y(N850) );
  NOR2X1 U7416 ( .A(n9742), .B(n8877), .Y(N849) );
  NOR2X1 U7417 ( .A(n9741), .B(n8877), .Y(N848) );
  NOR2X1 U7418 ( .A(n9740), .B(n8877), .Y(N847) );
  NOR2X1 U7419 ( .A(n9739), .B(n8877), .Y(N846) );
  NOR2X1 U7420 ( .A(n9738), .B(n8877), .Y(N845) );
  NOR2X1 U7421 ( .A(n9737), .B(n8877), .Y(N844) );
  NOR2X1 U7422 ( .A(n9736), .B(n8877), .Y(N843) );
  NOR2X1 U7423 ( .A(n9735), .B(n8877), .Y(N842) );
  NOR2X1 U7424 ( .A(n9734), .B(n8877), .Y(N841) );
  NOR2X1 U7425 ( .A(n9733), .B(n8877), .Y(N840) );
  NOR2X1 U7426 ( .A(n9732), .B(n8877), .Y(N839) );
  NOR2X1 U7427 ( .A(n9731), .B(n8876), .Y(N838) );
  NOR2X1 U7428 ( .A(n9730), .B(n8876), .Y(N837) );
  NOR2X1 U7429 ( .A(n9729), .B(n8876), .Y(N836) );
  NOR2X1 U7430 ( .A(n9728), .B(n8876), .Y(N835) );
  NOR2X1 U7431 ( .A(n9727), .B(n8876), .Y(N834) );
  NOR2X1 U7432 ( .A(n9726), .B(n8876), .Y(N833) );
  NOR2X1 U7433 ( .A(n9725), .B(n8876), .Y(N832) );
  NOR2X1 U7434 ( .A(n9724), .B(n8876), .Y(N831) );
  NOR2X1 U7435 ( .A(n9723), .B(n8876), .Y(N830) );
  NOR2X1 U7436 ( .A(n9722), .B(n8876), .Y(N829) );
  NOR2X1 U7437 ( .A(n9721), .B(n8876), .Y(N828) );
  NOR2X1 U7438 ( .A(n9720), .B(n8876), .Y(N827) );
  NOR2X1 U7439 ( .A(n9719), .B(n8876), .Y(N826) );
  NOR2X1 U7440 ( .A(n9718), .B(n8875), .Y(N825) );
  NOR2X1 U7441 ( .A(n10165), .B(n8875), .Y(N824) );
  NOR2X1 U7442 ( .A(n10164), .B(n8875), .Y(N823) );
  NOR2X1 U7443 ( .A(n10163), .B(n8875), .Y(N822) );
  NOR2X1 U7444 ( .A(n10162), .B(n8875), .Y(N821) );
  NOR2X1 U7445 ( .A(n10161), .B(n8875), .Y(N820) );
  NOR2X1 U7446 ( .A(n10160), .B(n8875), .Y(N819) );
  NOR2X1 U7447 ( .A(n10159), .B(n8875), .Y(N818) );
  NOR2X1 U7448 ( .A(n10158), .B(n8875), .Y(N817) );
  NOR2X1 U7449 ( .A(n10157), .B(n8875), .Y(N816) );
  NOR2X1 U7450 ( .A(n10156), .B(n8875), .Y(N815) );
  NOR2X1 U7451 ( .A(n10155), .B(n8875), .Y(N814) );
  NOR2X1 U7452 ( .A(n10154), .B(n8875), .Y(N813) );
  NOR2X1 U7453 ( .A(n10153), .B(n8874), .Y(N812) );
  NOR2X1 U7454 ( .A(n10152), .B(n8874), .Y(N811) );
  NOR2X1 U7455 ( .A(n10151), .B(n8874), .Y(N810) );
  NOR2X1 U7456 ( .A(n10150), .B(n8874), .Y(N809) );
  NOR2X1 U7457 ( .A(n10149), .B(n8874), .Y(N808) );
  NOR2X1 U7458 ( .A(n10148), .B(n8874), .Y(N807) );
  NOR2X1 U7459 ( .A(n10147), .B(n8874), .Y(N806) );
  NOR2X1 U7460 ( .A(n10146), .B(n8874), .Y(N805) );
  NOR2X1 U7461 ( .A(n10145), .B(n8874), .Y(N804) );
  NOR2X1 U7462 ( .A(n10144), .B(n8874), .Y(N803) );
  NOR2X1 U7463 ( .A(n10143), .B(n8874), .Y(N802) );
  NOR2X1 U7464 ( .A(n10142), .B(n8874), .Y(N801) );
  NOR2X1 U7465 ( .A(n10141), .B(n8874), .Y(N800) );
  NOR2X1 U7466 ( .A(n10140), .B(n8873), .Y(N799) );
  NOR2X1 U7467 ( .A(n10139), .B(n8873), .Y(N798) );
  NOR2X1 U7468 ( .A(n10138), .B(n8873), .Y(N797) );
  NOR2X1 U7469 ( .A(n10137), .B(n8873), .Y(N796) );
  NOR2X1 U7470 ( .A(n10136), .B(n8873), .Y(N795) );
  NOR2X1 U7471 ( .A(n10135), .B(n8873), .Y(N794) );
  NOR2X1 U7472 ( .A(n10134), .B(n8873), .Y(N793) );
  NOR2X1 U7473 ( .A(n9909), .B(n8873), .Y(N792) );
  NOR2X1 U7474 ( .A(n9908), .B(n8873), .Y(N791) );
  NOR2X1 U7475 ( .A(n9907), .B(n8873), .Y(N790) );
  NOR2X1 U7476 ( .A(n9906), .B(n8873), .Y(N789) );
  NOR2X1 U7477 ( .A(n9905), .B(n8873), .Y(N788) );
  NOR2X1 U7478 ( .A(n9904), .B(n8873), .Y(N787) );
  NOR2X1 U7479 ( .A(n9903), .B(n8872), .Y(N786) );
  NOR2X1 U7480 ( .A(n9902), .B(n8872), .Y(N785) );
  NOR2X1 U7481 ( .A(n9901), .B(n8872), .Y(N784) );
  NOR2X1 U7482 ( .A(n9900), .B(n8872), .Y(N783) );
  NOR2X1 U7483 ( .A(n9899), .B(n8872), .Y(N782) );
  NOR2X1 U7484 ( .A(n9898), .B(n8872), .Y(N781) );
  NOR2X1 U7485 ( .A(n9897), .B(n8872), .Y(N780) );
  NOR2X1 U7486 ( .A(n9896), .B(n8872), .Y(N779) );
  NOR2X1 U7487 ( .A(n9895), .B(n8872), .Y(N778) );
  NOR2X1 U7488 ( .A(n9894), .B(n8872), .Y(N777) );
  NOR2X1 U7489 ( .A(n9893), .B(n8872), .Y(N776) );
  NOR2X1 U7490 ( .A(n9892), .B(n8872), .Y(N775) );
  NOR2X1 U7491 ( .A(n9891), .B(n8872), .Y(N774) );
  NOR2X1 U7492 ( .A(n9890), .B(n8871), .Y(N773) );
  NOR2X1 U7493 ( .A(n9889), .B(n8871), .Y(N772) );
  NOR2X1 U7494 ( .A(n9888), .B(n8871), .Y(N771) );
  NOR2X1 U7495 ( .A(n9887), .B(n8871), .Y(N770) );
  NOR2X1 U7496 ( .A(n9886), .B(n8871), .Y(N769) );
  NOR2X1 U7497 ( .A(n9885), .B(n8871), .Y(N768) );
  NOR2X1 U7498 ( .A(n9884), .B(n8871), .Y(N767) );
  NOR2X1 U7499 ( .A(n9883), .B(n8871), .Y(N766) );
  NOR2X1 U7500 ( .A(n9882), .B(n8871), .Y(N765) );
  NOR2X1 U7501 ( .A(n9881), .B(n8871), .Y(N764) );
  NOR2X1 U7502 ( .A(n9880), .B(n8871), .Y(N763) );
  NOR2X1 U7503 ( .A(n9879), .B(n8871), .Y(N762) );
  NOR2X1 U7504 ( .A(n9878), .B(n8871), .Y(N761) );
  NOR2X1 U7505 ( .A(n10037), .B(n8870), .Y(N760) );
  NOR2X1 U7506 ( .A(n10036), .B(n8870), .Y(N759) );
  NOR2X1 U7507 ( .A(n10035), .B(n8870), .Y(N758) );
  NOR2X1 U7508 ( .A(n10034), .B(n8870), .Y(N757) );
  NOR2X1 U7509 ( .A(n10033), .B(n8870), .Y(N756) );
  NOR2X1 U7510 ( .A(n10032), .B(n8870), .Y(N755) );
  NOR2X1 U7511 ( .A(n10031), .B(n8870), .Y(N754) );
  NOR2X1 U7512 ( .A(n10030), .B(n8870), .Y(N753) );
  NOR2X1 U7513 ( .A(n10029), .B(n8870), .Y(N752) );
  NOR2X1 U7514 ( .A(n10028), .B(n8870), .Y(N751) );
  NOR2X1 U7515 ( .A(n10027), .B(n8870), .Y(N750) );
  NOR2X1 U7516 ( .A(n10026), .B(n8870), .Y(N749) );
  NOR2X1 U7517 ( .A(n10025), .B(n8870), .Y(N748) );
  NOR2X1 U7518 ( .A(n10024), .B(n8869), .Y(N747) );
  NOR2X1 U7519 ( .A(n10023), .B(n8869), .Y(N746) );
  NOR2X1 U7520 ( .A(n10022), .B(n8869), .Y(N745) );
  NOR2X1 U7521 ( .A(n10021), .B(n8869), .Y(N744) );
  NOR2X1 U7522 ( .A(n10020), .B(n8869), .Y(N743) );
  NOR2X1 U7523 ( .A(n10019), .B(n8869), .Y(N742) );
  NOR2X1 U7524 ( .A(n10018), .B(n8869), .Y(N741) );
  NOR2X1 U7525 ( .A(n10017), .B(n8869), .Y(N740) );
  NOR2X1 U7526 ( .A(n10016), .B(n8869), .Y(N739) );
  NOR2X1 U7527 ( .A(n10015), .B(n8869), .Y(N738) );
  NOR2X1 U7528 ( .A(n10014), .B(n8869), .Y(N737) );
  NOR2X1 U7529 ( .A(n10013), .B(n8869), .Y(N736) );
  NOR2X1 U7530 ( .A(n10012), .B(n8869), .Y(N735) );
  NOR2X1 U7531 ( .A(n10011), .B(n8868), .Y(N734) );
  NOR2X1 U7532 ( .A(n10010), .B(n8868), .Y(N733) );
  NOR2X1 U7533 ( .A(n10009), .B(n8868), .Y(N732) );
  NOR2X1 U7534 ( .A(n10008), .B(n8868), .Y(N731) );
  NOR2X1 U7535 ( .A(n10007), .B(n8868), .Y(N730) );
  NOR2X1 U7536 ( .A(n10006), .B(n8868), .Y(N729) );
  NOR2X1 U7537 ( .A(n9781), .B(n8868), .Y(N728) );
  NOR2X1 U7538 ( .A(n9780), .B(n8868), .Y(N727) );
  NOR2X1 U7539 ( .A(n9779), .B(n8868), .Y(N726) );
  NOR2X1 U7540 ( .A(n9778), .B(n8868), .Y(N725) );
  NOR2X1 U7541 ( .A(n9777), .B(n8868), .Y(N724) );
  NOR2X1 U7542 ( .A(n9776), .B(n8868), .Y(N723) );
  NOR2X1 U7543 ( .A(n9775), .B(n8868), .Y(N722) );
  NOR2X1 U7544 ( .A(n9774), .B(n8867), .Y(N721) );
  NOR2X1 U7545 ( .A(n9773), .B(n8867), .Y(N720) );
  NOR2X1 U7546 ( .A(n9772), .B(n8867), .Y(N719) );
  NOR2X1 U7547 ( .A(n9771), .B(n8867), .Y(N718) );
  NOR2X1 U7548 ( .A(n9770), .B(n8867), .Y(N717) );
  NOR2X1 U7549 ( .A(n9769), .B(n8867), .Y(N716) );
  NOR2X1 U7550 ( .A(n9768), .B(n8867), .Y(N715) );
  NOR2X1 U7551 ( .A(n9767), .B(n8867), .Y(N714) );
  NOR2X1 U7552 ( .A(n9766), .B(n8867), .Y(N713) );
  NOR2X1 U7553 ( .A(n9765), .B(n8867), .Y(N712) );
  NOR2X1 U7554 ( .A(n9764), .B(n8867), .Y(N711) );
  NOR2X1 U7555 ( .A(n9763), .B(n8867), .Y(N710) );
  NOR2X1 U7556 ( .A(n9762), .B(n8867), .Y(N709) );
  NOR2X1 U7557 ( .A(n9761), .B(n8866), .Y(N708) );
  NOR2X1 U7558 ( .A(n9760), .B(n8866), .Y(N707) );
  NOR2X1 U7559 ( .A(n9759), .B(n8866), .Y(N706) );
  NOR2X1 U7560 ( .A(n9758), .B(n8866), .Y(N705) );
  NOR2X1 U7561 ( .A(n9757), .B(n8866), .Y(N704) );
  NOR2X1 U7562 ( .A(n9756), .B(n8866), .Y(N703) );
  NOR2X1 U7563 ( .A(n9755), .B(n8866), .Y(N702) );
  NOR2X1 U7564 ( .A(n9754), .B(n8866), .Y(N701) );
  NOR2X1 U7565 ( .A(n9753), .B(n8866), .Y(N700) );
  NOR2X1 U7566 ( .A(n9752), .B(n8866), .Y(N699) );
  NOR2X1 U7567 ( .A(n9751), .B(n8866), .Y(N698) );
  NOR2X1 U7568 ( .A(n9750), .B(n8866), .Y(N697) );
  NOR2X1 U7569 ( .A(n10101), .B(n8866), .Y(N696) );
  NOR2X1 U7570 ( .A(n10100), .B(n8865), .Y(N695) );
  NOR2X1 U7571 ( .A(n10099), .B(n8865), .Y(N694) );
  NOR2X1 U7572 ( .A(n10098), .B(n8865), .Y(N693) );
  NOR2X1 U7573 ( .A(n10097), .B(n8865), .Y(N692) );
  NOR2X1 U7574 ( .A(n10096), .B(n8865), .Y(N691) );
  NOR2X1 U7575 ( .A(n10095), .B(n8865), .Y(N690) );
  NOR2X1 U7576 ( .A(n10094), .B(n8865), .Y(N689) );
  NOR2X1 U7577 ( .A(n10093), .B(n8865), .Y(N688) );
  NOR2X1 U7578 ( .A(n10092), .B(n8865), .Y(N687) );
  NOR2X1 U7579 ( .A(n10091), .B(n8865), .Y(N686) );
  NOR2X1 U7580 ( .A(n10090), .B(n8865), .Y(N685) );
  NOR2X1 U7581 ( .A(n10089), .B(n8865), .Y(N684) );
  NOR2X1 U7582 ( .A(n10088), .B(n8865), .Y(N683) );
  NOR2X1 U7583 ( .A(n10087), .B(n8864), .Y(N682) );
  NOR2X1 U7584 ( .A(n10086), .B(n8864), .Y(N681) );
  NOR2X1 U7585 ( .A(n10085), .B(n8864), .Y(N680) );
  NOR2X1 U7586 ( .A(n10084), .B(n8864), .Y(N679) );
  NOR2X1 U7587 ( .A(n10083), .B(n8864), .Y(N678) );
  NOR2X1 U7588 ( .A(n10082), .B(n8864), .Y(N677) );
  NOR2X1 U7589 ( .A(n10081), .B(n8864), .Y(N676) );
  NOR2X1 U7590 ( .A(n10080), .B(n8864), .Y(N675) );
  NOR2X1 U7591 ( .A(n10079), .B(n8864), .Y(N674) );
  NOR2X1 U7592 ( .A(n10078), .B(n8864), .Y(N673) );
  NOR2X1 U7593 ( .A(n10077), .B(n8864), .Y(N672) );
  NOR2X1 U7594 ( .A(n10076), .B(n8864), .Y(N671) );
  NOR2X1 U7595 ( .A(n10075), .B(n8864), .Y(N670) );
  NOR2X1 U7596 ( .A(n10074), .B(n8863), .Y(N669) );
  NOR2X1 U7597 ( .A(n10073), .B(n8863), .Y(N668) );
  NOR2X1 U7598 ( .A(n10072), .B(n8863), .Y(N667) );
  NOR2X1 U7599 ( .A(n10071), .B(n8863), .Y(N666) );
  NOR2X1 U7600 ( .A(n10070), .B(n8863), .Y(N665) );
  NOR2X1 U7601 ( .A(n9845), .B(n8863), .Y(N664) );
  NOR2X1 U7602 ( .A(n9844), .B(n8863), .Y(N663) );
  NOR2X1 U7603 ( .A(n9843), .B(n8863), .Y(N662) );
  NOR2X1 U7604 ( .A(n9842), .B(n8863), .Y(N661) );
  NOR2X1 U7605 ( .A(n9841), .B(n8863), .Y(N660) );
  NOR2X1 U7606 ( .A(n9840), .B(n8863), .Y(N659) );
  NOR2X1 U7607 ( .A(n9839), .B(n8863), .Y(N658) );
  NOR2X1 U7608 ( .A(n9838), .B(n8863), .Y(N657) );
  NOR2X1 U7609 ( .A(n9837), .B(n8862), .Y(N656) );
  NOR2X1 U7610 ( .A(n9836), .B(n8862), .Y(N655) );
  NOR2X1 U7611 ( .A(n9835), .B(n8862), .Y(N654) );
  NOR2X1 U7612 ( .A(n9834), .B(n8862), .Y(N653) );
  NOR2X1 U7613 ( .A(n9833), .B(n8862), .Y(N652) );
  NOR2X1 U7614 ( .A(n9832), .B(n8862), .Y(N651) );
  NOR2X1 U7615 ( .A(n9831), .B(n8862), .Y(N650) );
  NOR2X1 U7616 ( .A(n9830), .B(n8862), .Y(N649) );
  NOR2X1 U7617 ( .A(n9829), .B(n8862), .Y(N648) );
  NOR2X1 U7618 ( .A(n9828), .B(n8862), .Y(N647) );
  NOR2X1 U7619 ( .A(n9827), .B(n8862), .Y(N646) );
  NOR2X1 U7620 ( .A(n9826), .B(n8862), .Y(N645) );
  NOR2X1 U7621 ( .A(n9825), .B(n8862), .Y(N644) );
  NOR2X1 U7622 ( .A(n9824), .B(n8861), .Y(N643) );
  NOR2X1 U7623 ( .A(n9823), .B(n8861), .Y(N642) );
  NOR2X1 U7624 ( .A(n9822), .B(n8861), .Y(N641) );
  NOR2X1 U7625 ( .A(n9821), .B(n8861), .Y(N640) );
  NOR2X1 U7626 ( .A(n9820), .B(n8861), .Y(N639) );
  NOR2X1 U7627 ( .A(n9819), .B(n8861), .Y(N638) );
  NOR2X1 U7628 ( .A(n9818), .B(n8861), .Y(N637) );
  NOR2X1 U7629 ( .A(n9817), .B(n8861), .Y(N636) );
  NOR2X1 U7630 ( .A(n9816), .B(n8861), .Y(N635) );
  NOR2X1 U7631 ( .A(n9815), .B(n8861), .Y(N634) );
  NOR2X1 U7632 ( .A(n9814), .B(n8861), .Y(N633) );
  NOR2X1 U7633 ( .A(n9973), .B(n8861), .Y(N632) );
  NOR2X1 U7634 ( .A(n9972), .B(n8861), .Y(N631) );
  NOR2X1 U7635 ( .A(n9971), .B(n8860), .Y(N630) );
  NOR2X1 U7636 ( .A(n9970), .B(n8860), .Y(N629) );
  NOR2X1 U7637 ( .A(n9969), .B(n8860), .Y(N628) );
  NOR2X1 U7638 ( .A(n9968), .B(n8860), .Y(N627) );
  NOR2X1 U7639 ( .A(n9967), .B(n8860), .Y(N626) );
  NOR2X1 U7640 ( .A(n9966), .B(n8860), .Y(N625) );
  NOR2X1 U7641 ( .A(n9965), .B(n8860), .Y(N624) );
  NOR2X1 U7642 ( .A(n9964), .B(n8860), .Y(N623) );
  NOR2X1 U7643 ( .A(n9963), .B(n8860), .Y(N622) );
  NOR2X1 U7644 ( .A(n9962), .B(n8860), .Y(N621) );
  NOR2X1 U7645 ( .A(n9961), .B(n8860), .Y(N620) );
  NOR2X1 U7646 ( .A(n9960), .B(n8860), .Y(N619) );
  NOR2X1 U7647 ( .A(n9959), .B(n8860), .Y(N618) );
  NOR2X1 U7648 ( .A(n9958), .B(n8859), .Y(N617) );
  NOR2X1 U7649 ( .A(n9957), .B(n8859), .Y(N616) );
  NOR2X1 U7650 ( .A(n9956), .B(n8859), .Y(N615) );
  NOR2X1 U7651 ( .A(n9955), .B(n8859), .Y(N614) );
  NOR2X1 U7652 ( .A(n9954), .B(n8859), .Y(N613) );
  NOR2X1 U7653 ( .A(n9953), .B(n8859), .Y(N612) );
  NOR2X1 U7654 ( .A(n9952), .B(n8859), .Y(N611) );
  NOR2X1 U7655 ( .A(n9951), .B(n8859), .Y(N610) );
  NOR2X1 U7656 ( .A(n9950), .B(n8859), .Y(N609) );
  NOR2X1 U7657 ( .A(n9949), .B(n8859), .Y(N608) );
  NOR2X1 U7658 ( .A(n9948), .B(n8859), .Y(N607) );
  NOR2X1 U7659 ( .A(n9947), .B(n8859), .Y(N606) );
  NOR2X1 U7660 ( .A(n9946), .B(n8859), .Y(N605) );
  NOR2X1 U7661 ( .A(n9945), .B(n8858), .Y(N604) );
  NOR2X1 U7662 ( .A(n9944), .B(n8858), .Y(N603) );
  NOR2X1 U7663 ( .A(n9943), .B(n8858), .Y(N602) );
  NOR2X1 U7664 ( .A(n9942), .B(n8858), .Y(N601) );
  NOR2X1 U7665 ( .A(n9717), .B(n8858), .Y(N600) );
  NOR2X1 U7666 ( .A(n9716), .B(n8858), .Y(N599) );
  NOR2X1 U7667 ( .A(n9715), .B(n8858), .Y(N598) );
  NOR2X1 U7668 ( .A(n9714), .B(n8858), .Y(N597) );
  NOR2X1 U7669 ( .A(n9713), .B(n8858), .Y(N596) );
  NOR2X1 U7670 ( .A(n9712), .B(n8858), .Y(N595) );
  NOR2X1 U7671 ( .A(n9711), .B(n8858), .Y(N594) );
  NOR2X1 U7672 ( .A(n9710), .B(n8858), .Y(N593) );
  NOR2X1 U7673 ( .A(n9709), .B(n8858), .Y(N592) );
  NOR2X1 U7674 ( .A(n9708), .B(n8857), .Y(N591) );
  NOR2X1 U7675 ( .A(n9707), .B(n8857), .Y(N590) );
  NOR2X1 U7676 ( .A(n9706), .B(n8857), .Y(N589) );
  NOR2X1 U7677 ( .A(n9705), .B(n8857), .Y(N588) );
  NOR2X1 U7678 ( .A(n9704), .B(n8857), .Y(N587) );
  NOR2X1 U7679 ( .A(n9703), .B(n8857), .Y(N586) );
  NOR2X1 U7680 ( .A(n9702), .B(n8857), .Y(N585) );
  NOR2X1 U7681 ( .A(n9701), .B(n8857), .Y(N584) );
  NOR2X1 U7682 ( .A(n9700), .B(n8857), .Y(N583) );
  NOR2X1 U7683 ( .A(n9699), .B(n8857), .Y(N582) );
  NOR2X1 U7684 ( .A(n9698), .B(n8857), .Y(N581) );
  NOR2X1 U7685 ( .A(n9697), .B(n8857), .Y(N580) );
  NOR2X1 U7686 ( .A(n9696), .B(n8857), .Y(N579) );
  NOR2X1 U7687 ( .A(n9695), .B(n8856), .Y(N578) );
  NOR2X1 U7688 ( .A(n9694), .B(n8856), .Y(N577) );
  NOR2X1 U7689 ( .A(n9693), .B(n8856), .Y(N576) );
  NOR2X1 U7690 ( .A(n9692), .B(n8856), .Y(N575) );
  NOR2X1 U7691 ( .A(n9691), .B(n8856), .Y(N574) );
  NOR2X1 U7692 ( .A(n9690), .B(n8856), .Y(N573) );
  NOR2X1 U7693 ( .A(n9689), .B(n8856), .Y(N572) );
  NOR2X1 U7694 ( .A(n9688), .B(n8856), .Y(N571) );
  NOR2X1 U7695 ( .A(n9687), .B(n8856), .Y(N570) );
  NOR2X1 U7696 ( .A(n9686), .B(n8856), .Y(N569) );
  NOR2X1 U7697 ( .A(n9246), .B(n9242), .Y(N1394) );
  NOR2X1 U7698 ( .A(n9246), .B(n9239), .Y(N1393) );
  NOR2X1 U7699 ( .A(n9246), .B(n9236), .Y(N1392) );
  NOR2X1 U7700 ( .A(n9246), .B(n9233), .Y(N1391) );
  NOR2X1 U7701 ( .A(n9246), .B(n9230), .Y(N1390) );
  NOR2X1 U7702 ( .A(n9246), .B(n9227), .Y(N1389) );
  NOR2X1 U7703 ( .A(n9246), .B(n9224), .Y(N1388) );
  NOR2X1 U7704 ( .A(n9246), .B(n9221), .Y(N1387) );
  NOR2X1 U7705 ( .A(n9246), .B(n9218), .Y(N1386) );
  NOR2X1 U7706 ( .A(n9246), .B(n9215), .Y(N1385) );
  NOR2X1 U7707 ( .A(n9246), .B(n9212), .Y(N1384) );
  NOR2X1 U7708 ( .A(n9246), .B(n9209), .Y(N1383) );
  NOR2X1 U7709 ( .A(n9246), .B(n9206), .Y(N1382) );
  NOR2X1 U7710 ( .A(n9246), .B(n9203), .Y(N1381) );
  NOR2X1 U7711 ( .A(n9246), .B(n9200), .Y(N1380) );
  NOR2X1 U7712 ( .A(n9246), .B(n9198), .Y(N1379) );
  CLKINVX1 U7713 ( .A(n9247), .Y(n9246) );
  NOR2X1 U7714 ( .A(n6192), .B(n10474), .Y(n9247) );
  NOR2X1 U7715 ( .A(n9245), .B(n9242), .Y(N1378) );
  CLKINVX1 U7716 ( .A(BF2I_a_er_n[15]), .Y(n9242) );
  NOR2X1 U7717 ( .A(n9245), .B(n9239), .Y(N1377) );
  CLKINVX1 U7718 ( .A(BF2I_a_er_n[14]), .Y(n9239) );
  NOR2X1 U7719 ( .A(n9245), .B(n9236), .Y(N1376) );
  CLKINVX1 U7720 ( .A(BF2I_a_er_n[13]), .Y(n9236) );
  NOR2X1 U7721 ( .A(n9245), .B(n9233), .Y(N1375) );
  CLKINVX1 U7722 ( .A(BF2I_a_er_n[12]), .Y(n9233) );
  NOR2X1 U7723 ( .A(n9245), .B(n9230), .Y(N1374) );
  CLKINVX1 U7724 ( .A(BF2I_a_er_n[11]), .Y(n9230) );
  NOR2X1 U7725 ( .A(n9245), .B(n9227), .Y(N1373) );
  CLKINVX1 U7726 ( .A(BF2I_a_er_n[10]), .Y(n9227) );
  NOR2X1 U7727 ( .A(n9245), .B(n9224), .Y(N1372) );
  CLKINVX1 U7728 ( .A(BF2I_a_er_n[9]), .Y(n9224) );
  NOR2X1 U7729 ( .A(n9245), .B(n9221), .Y(N1371) );
  CLKINVX1 U7730 ( .A(BF2I_a_er_n[8]), .Y(n9221) );
  NOR2X1 U7731 ( .A(n9245), .B(n9218), .Y(N1370) );
  CLKINVX1 U7732 ( .A(BF2I_a_er_n[7]), .Y(n9218) );
  NOR2X1 U7733 ( .A(n9245), .B(n9215), .Y(N1369) );
  CLKINVX1 U7734 ( .A(BF2I_a_er_n[6]), .Y(n9215) );
  NOR2X1 U7735 ( .A(n9245), .B(n9212), .Y(N1368) );
  CLKINVX1 U7736 ( .A(BF2I_a_er_n[5]), .Y(n9212) );
  NOR2X1 U7737 ( .A(n9245), .B(n9209), .Y(N1367) );
  CLKINVX1 U7738 ( .A(BF2I_a_er_n[4]), .Y(n9209) );
  NOR2X1 U7739 ( .A(n9245), .B(n9206), .Y(N1366) );
  CLKINVX1 U7740 ( .A(BF2I_a_er_n[3]), .Y(n9206) );
  NOR2X1 U7741 ( .A(n9245), .B(n9203), .Y(N1365) );
  CLKINVX1 U7742 ( .A(BF2I_a_er_n[2]), .Y(n9203) );
  NOR2X1 U7743 ( .A(n9245), .B(n9200), .Y(N1364) );
  CLKINVX1 U7744 ( .A(BF2I_a_er_n[1]), .Y(n9200) );
  CLKINVX1 U7745 ( .A(BF2I_a_er_n[0]), .Y(n9198) );
  NOR2X1 U7746 ( .A(n10474), .B(n11213), .Y(mult_add_355_aco_b) );
  NOR2X1 U7747 ( .A(n11212), .B(n9573), .Y(N1362) );
  NAND2X1 U7748 ( .A(N43), .B(n11218), .Y(n9573) );
  NOR2X1 U7749 ( .A(n11213), .B(n9574), .Y(N1361) );
  MXI2X1 U7750 ( .A(d32[30]), .B(N42), .S0(n11218), .Y(n9574) );
  NOR2X1 U7751 ( .A(n11212), .B(n9575), .Y(N1360) );
  MXI2X1 U7752 ( .A(d32[29]), .B(N41), .S0(n11219), .Y(n9575) );
  NOR2X1 U7753 ( .A(n11213), .B(n9576), .Y(N1359) );
  MXI2X1 U7754 ( .A(d32[28]), .B(N40), .S0(n11218), .Y(n9576) );
  NOR2X1 U7755 ( .A(n11212), .B(n9577), .Y(N1358) );
  MXI2X1 U7756 ( .A(d32[27]), .B(N39), .S0(n11219), .Y(n9577) );
  NOR2X1 U7757 ( .A(n11213), .B(n9578), .Y(N1357) );
  MXI2X1 U7758 ( .A(d32[26]), .B(N38), .S0(n11218), .Y(n9578) );
  NOR2X1 U7759 ( .A(n11212), .B(n9564), .Y(N1356) );
  MXI2X1 U7760 ( .A(d32[25]), .B(N37), .S0(n11219), .Y(n9564) );
  NOR2X1 U7761 ( .A(n11213), .B(n9565), .Y(N1355) );
  MXI2X1 U7762 ( .A(d32[24]), .B(N36), .S0(n11218), .Y(n9565) );
  NOR2X1 U7763 ( .A(n11212), .B(n9566), .Y(N1354) );
  MXI2X1 U7764 ( .A(d32[23]), .B(N35), .S0(n11219), .Y(n9566) );
  NOR2X1 U7765 ( .A(n11213), .B(n9567), .Y(N1353) );
  MXI2X1 U7766 ( .A(d32[22]), .B(N34), .S0(n11218), .Y(n9567) );
  NOR2X1 U7767 ( .A(n11212), .B(n9568), .Y(N1352) );
  MXI2X1 U7768 ( .A(d32[21]), .B(N33), .S0(n11219), .Y(n9568) );
  NOR2X1 U7769 ( .A(n11213), .B(n9569), .Y(N1351) );
  MXI2X1 U7770 ( .A(d32[20]), .B(N32), .S0(n11218), .Y(n9569) );
  NOR2X1 U7771 ( .A(n11212), .B(n9570), .Y(N1350) );
  MXI2X1 U7772 ( .A(d32[19]), .B(N31), .S0(n11219), .Y(n9570) );
  NOR2X1 U7773 ( .A(n11213), .B(n9571), .Y(N1349) );
  MXI2X1 U7774 ( .A(d32[18]), .B(N30), .S0(n11218), .Y(n9571) );
  NOR2X1 U7775 ( .A(n11212), .B(n9572), .Y(N1348) );
  MXI2X1 U7776 ( .A(d32[17]), .B(N29), .S0(n11219), .Y(n9572) );
  NOR2X1 U7777 ( .A(n11213), .B(n9579), .Y(N1347) );
  MXI2X1 U7778 ( .A(d32[16]), .B(N28), .S0(n11218), .Y(n9579) );
  NOR2X1 U7779 ( .A(n9581), .B(n6196), .Y(N1233) );
  NOR2X1 U7780 ( .A(n9581), .B(n6197), .Y(N1232) );
  NOR2X1 U7781 ( .A(n9581), .B(n6198), .Y(N1231) );
  NOR2X1 U7782 ( .A(n9581), .B(n6199), .Y(N1230) );
  CLKINVX1 U7783 ( .A(n6071), .Y(n9581) );
  NOR2X1 U7784 ( .A(n9582), .B(n9685), .Y(n6071) );
  OAI22XL U7785 ( .A0(n2860), .A1(n9583), .B0(n9584), .B1(n9585), .Y(N1224) );
  CLKINVX1 U7786 ( .A(fft_d[31]), .Y(n9585) );
  OAI22XL U7787 ( .A0(n2870), .A1(n9583), .B0(n9584), .B1(n9586), .Y(N1223) );
  CLKINVX1 U7788 ( .A(fft_d[30]), .Y(n9586) );
  OAI22XL U7789 ( .A0(n2880), .A1(n9583), .B0(n9584), .B1(n9587), .Y(N1222) );
  CLKINVX1 U7790 ( .A(fft_d[29]), .Y(n9587) );
  OAI22XL U7791 ( .A0(n2890), .A1(n9583), .B0(n9584), .B1(n9588), .Y(N1221) );
  CLKINVX1 U7792 ( .A(fft_d[28]), .Y(n9588) );
  OAI22XL U7793 ( .A0(n290), .A1(n9583), .B0(n9584), .B1(n9589), .Y(N1220) );
  CLKINVX1 U7794 ( .A(fft_d[27]), .Y(n9589) );
  OAI22XL U7795 ( .A0(n291), .A1(n9583), .B0(n9584), .B1(n9590), .Y(N1219) );
  CLKINVX1 U7796 ( .A(fft_d[26]), .Y(n9590) );
  OAI22XL U7797 ( .A0(n292), .A1(n9583), .B0(n9584), .B1(n9591), .Y(N1218) );
  CLKINVX1 U7798 ( .A(fft_d[25]), .Y(n9591) );
  OAI22XL U7799 ( .A0(n293), .A1(n9583), .B0(n9584), .B1(n9592), .Y(N1217) );
  CLKINVX1 U7800 ( .A(fft_d[24]), .Y(n9592) );
  OAI22XL U7801 ( .A0(n294), .A1(n9583), .B0(n9584), .B1(n9593), .Y(N1216) );
  CLKINVX1 U7802 ( .A(fft_d[23]), .Y(n9593) );
  OAI22XL U7803 ( .A0(n295), .A1(n9583), .B0(n9584), .B1(n9594), .Y(N1215) );
  CLKINVX1 U7804 ( .A(fft_d[22]), .Y(n9594) );
  OAI22XL U7805 ( .A0(n296), .A1(n9583), .B0(n9584), .B1(n9595), .Y(N1214) );
  CLKINVX1 U7806 ( .A(fft_d[21]), .Y(n9595) );
  OAI22XL U7807 ( .A0(n297), .A1(n9583), .B0(n9584), .B1(n9596), .Y(N1213) );
  CLKINVX1 U7808 ( .A(fft_d[20]), .Y(n9596) );
  OAI22XL U7809 ( .A0(n298), .A1(n9583), .B0(n9584), .B1(n9597), .Y(N1212) );
  CLKINVX1 U7810 ( .A(fft_d[19]), .Y(n9597) );
  OAI22XL U7811 ( .A0(n299), .A1(n9583), .B0(n9584), .B1(n9598), .Y(N1211) );
  CLKINVX1 U7812 ( .A(fft_d[18]), .Y(n9598) );
  OAI22XL U7813 ( .A0(n3000), .A1(n9583), .B0(n9584), .B1(n9599), .Y(N1210) );
  CLKINVX1 U7814 ( .A(fft_d[17]), .Y(n9599) );
  OAI22XL U7815 ( .A0(n3010), .A1(n9583), .B0(n9584), .B1(n9600), .Y(N1209) );
  CLKINVX1 U7816 ( .A(fft_d[16]), .Y(n9600) );
  OAI22XL U7817 ( .A0(n3020), .A1(n9583), .B0(n9584), .B1(n9601), .Y(N1208) );
  CLKINVX1 U7818 ( .A(fft_d[15]), .Y(n9601) );
  OAI22XL U7819 ( .A0(n3030), .A1(n9583), .B0(n9584), .B1(n9602), .Y(N1207) );
  CLKINVX1 U7820 ( .A(fft_d[14]), .Y(n9602) );
  OAI22XL U7821 ( .A0(n3040), .A1(n9583), .B0(n9584), .B1(n9603), .Y(N1206) );
  CLKINVX1 U7822 ( .A(fft_d[13]), .Y(n9603) );
  OAI22XL U7823 ( .A0(n3050), .A1(n9583), .B0(n9584), .B1(n9604), .Y(N1205) );
  CLKINVX1 U7824 ( .A(fft_d[12]), .Y(n9604) );
  OAI22XL U7825 ( .A0(n3060), .A1(n9583), .B0(n9584), .B1(n9605), .Y(N1204) );
  CLKINVX1 U7826 ( .A(fft_d[11]), .Y(n9605) );
  OAI22XL U7827 ( .A0(n30700), .A1(n9583), .B0(n9584), .B1(n9606), .Y(N1203)
         );
  CLKINVX1 U7828 ( .A(fft_d[10]), .Y(n9606) );
  OAI22XL U7829 ( .A0(n3080), .A1(n9583), .B0(n9584), .B1(n9607), .Y(N1202) );
  CLKINVX1 U7830 ( .A(fft_d[9]), .Y(n9607) );
  OAI22XL U7831 ( .A0(n3090), .A1(n9583), .B0(n9584), .B1(n9608), .Y(N1201) );
  CLKINVX1 U7832 ( .A(fft_d[8]), .Y(n9608) );
  OAI22XL U7833 ( .A0(n3100), .A1(n9583), .B0(n9584), .B1(n9609), .Y(N1200) );
  CLKINVX1 U7834 ( .A(fft_d[7]), .Y(n9609) );
  OAI22XL U7835 ( .A0(n3110), .A1(n9583), .B0(n9584), .B1(n9610), .Y(N1199) );
  CLKINVX1 U7836 ( .A(fft_d[6]), .Y(n9610) );
  OAI22XL U7837 ( .A0(n3120), .A1(n9583), .B0(n9584), .B1(n9611), .Y(N1198) );
  CLKINVX1 U7838 ( .A(fft_d[5]), .Y(n9611) );
  OAI22XL U7839 ( .A0(n3130), .A1(n9583), .B0(n9584), .B1(n9612), .Y(N1197) );
  CLKINVX1 U7840 ( .A(fft_d[4]), .Y(n9612) );
  OAI22XL U7841 ( .A0(n3140), .A1(n9583), .B0(n9584), .B1(n9613), .Y(N1196) );
  CLKINVX1 U7842 ( .A(fft_d[3]), .Y(n9613) );
  OAI22XL U7843 ( .A0(n3150), .A1(n9583), .B0(n9584), .B1(n9614), .Y(N1195) );
  CLKINVX1 U7844 ( .A(fft_d[2]), .Y(n9614) );
  OAI22XL U7845 ( .A0(n3160), .A1(n9583), .B0(n9584), .B1(n9615), .Y(N1194) );
  CLKINVX1 U7846 ( .A(fft_d[1]), .Y(n9615) );
  OAI22XL U7847 ( .A0(n2850), .A1(n9583), .B0(n9584), .B1(n9616), .Y(N1193) );
  OAI22XL U7848 ( .A0(n6196), .A1(n9583), .B0(counter[0]), .B1(n9617), .Y(
        N1192) );
  OAI2BB2XL U7849 ( .B0(n6197), .B1(n9583), .A0N(n9618), .A1N(n9619), .Y(N1191) );
  OAI21XL U7850 ( .A0(n6075), .A1(n6074), .B0(n9512), .Y(n9619) );
  OAI2BB2XL U7851 ( .B0(n6198), .B1(n9583), .A0N(n9618), .A1N(n9620), .Y(N1190) );
  AO21X1 U7852 ( .A0(counter[2]), .A1(n9512), .B0(n9621), .Y(n9620) );
  OAI2BB2XL U7853 ( .B0(n6199), .B1(n9583), .A0N(n9618), .A1N(n9622), .Y(N1189) );
  OAI21XL U7854 ( .A0(n6072), .A1(n9621), .B0(n9174), .Y(n9622) );
  CLKINVX1 U7855 ( .A(n9617), .Y(n9618) );
  NAND3BX1 U7856 ( .AN(n9623), .B(n9582), .C(n6193), .Y(n9583) );
  NAND3X1 U7857 ( .A(n6072), .B(n6074), .C(n9510), .Y(n9582) );
  NOR2X1 U7858 ( .A(counter[2]), .B(n6075), .Y(n9510) );
  OAI2BB1X1 U7859 ( .A0N(fft_d[31]), .A1N(n2860), .B0(n9624), .Y(n9623) );
  OAI21XL U7860 ( .A0(fft_d[31]), .A1(n2860), .B0(n9625), .Y(n9624) );
  OAI2BB1X1 U7861 ( .A0N(fft_d[30]), .A1N(n2870), .B0(n9626), .Y(n9625) );
  OAI221XL U7862 ( .A0(n2880), .A1(fft_d[29]), .B0(n2870), .B1(fft_d[30]), 
        .C0(n9627), .Y(n9626) );
  CLKINVX1 U7863 ( .A(n9628), .Y(n9627) );
  AOI221XL U7864 ( .A0(fft_d[28]), .A1(n2890), .B0(fft_d[29]), .B1(n2880), 
        .C0(n9629), .Y(n9628) );
  CLKINVX1 U7865 ( .A(n9630), .Y(n9629) );
  OAI221XL U7866 ( .A0(n290), .A1(fft_d[27]), .B0(n2890), .B1(fft_d[28]), .C0(
        n9631), .Y(n9630) );
  CLKINVX1 U7867 ( .A(n9632), .Y(n9631) );
  AOI221XL U7868 ( .A0(fft_d[26]), .A1(n291), .B0(fft_d[27]), .B1(n290), .C0(
        n9633), .Y(n9632) );
  CLKINVX1 U7869 ( .A(n9634), .Y(n9633) );
  OAI221XL U7870 ( .A0(n292), .A1(fft_d[25]), .B0(n291), .B1(fft_d[26]), .C0(
        n9635), .Y(n9634) );
  CLKINVX1 U7871 ( .A(n9636), .Y(n9635) );
  AOI221XL U7872 ( .A0(fft_d[24]), .A1(n293), .B0(fft_d[25]), .B1(n292), .C0(
        n9637), .Y(n9636) );
  CLKINVX1 U7873 ( .A(n9638), .Y(n9637) );
  OAI221XL U7874 ( .A0(n294), .A1(fft_d[23]), .B0(n293), .B1(fft_d[24]), .C0(
        n9639), .Y(n9638) );
  CLKINVX1 U7875 ( .A(n9640), .Y(n9639) );
  AOI221XL U7876 ( .A0(fft_d[22]), .A1(n295), .B0(fft_d[23]), .B1(n294), .C0(
        n9641), .Y(n9640) );
  CLKINVX1 U7877 ( .A(n9642), .Y(n9641) );
  OAI221XL U7878 ( .A0(n296), .A1(fft_d[21]), .B0(n295), .B1(fft_d[22]), .C0(
        n9643), .Y(n9642) );
  CLKINVX1 U7879 ( .A(n9644), .Y(n9643) );
  AOI221XL U7880 ( .A0(fft_d[20]), .A1(n297), .B0(fft_d[21]), .B1(n296), .C0(
        n9645), .Y(n9644) );
  CLKINVX1 U7881 ( .A(n9646), .Y(n9645) );
  OAI221XL U7882 ( .A0(n298), .A1(fft_d[19]), .B0(n297), .B1(fft_d[20]), .C0(
        n9647), .Y(n9646) );
  CLKINVX1 U7883 ( .A(n9648), .Y(n9647) );
  AOI221XL U7884 ( .A0(fft_d[18]), .A1(n299), .B0(fft_d[19]), .B1(n298), .C0(
        n9649), .Y(n9648) );
  CLKINVX1 U7885 ( .A(n9650), .Y(n9649) );
  OAI221XL U7886 ( .A0(n3000), .A1(fft_d[17]), .B0(n299), .B1(fft_d[18]), .C0(
        n9651), .Y(n9650) );
  CLKINVX1 U7887 ( .A(n9652), .Y(n9651) );
  AOI221XL U7888 ( .A0(fft_d[16]), .A1(n3010), .B0(fft_d[17]), .B1(n3000), 
        .C0(n9653), .Y(n9652) );
  CLKINVX1 U7889 ( .A(n9654), .Y(n9653) );
  OAI221XL U7890 ( .A0(n3020), .A1(fft_d[15]), .B0(n3010), .B1(fft_d[16]), 
        .C0(n9655), .Y(n9654) );
  CLKINVX1 U7891 ( .A(n9656), .Y(n9655) );
  AOI221XL U7892 ( .A0(fft_d[14]), .A1(n3030), .B0(fft_d[15]), .B1(n3020), 
        .C0(n9657), .Y(n9656) );
  CLKINVX1 U7893 ( .A(n9658), .Y(n9657) );
  OAI221XL U7894 ( .A0(n3040), .A1(fft_d[13]), .B0(n3030), .B1(fft_d[14]), 
        .C0(n9659), .Y(n9658) );
  CLKINVX1 U7895 ( .A(n9660), .Y(n9659) );
  AOI221XL U7896 ( .A0(fft_d[12]), .A1(n3050), .B0(fft_d[13]), .B1(n3040), 
        .C0(n9661), .Y(n9660) );
  CLKINVX1 U7897 ( .A(n9662), .Y(n9661) );
  OAI221XL U7898 ( .A0(n3060), .A1(fft_d[11]), .B0(n3050), .B1(fft_d[12]), 
        .C0(n9663), .Y(n9662) );
  CLKINVX1 U7899 ( .A(n9664), .Y(n9663) );
  AOI221XL U7900 ( .A0(fft_d[10]), .A1(n30700), .B0(fft_d[11]), .B1(n3060), 
        .C0(n9665), .Y(n9664) );
  CLKINVX1 U7901 ( .A(n9666), .Y(n9665) );
  OAI221XL U7902 ( .A0(n30700), .A1(fft_d[10]), .B0(n3080), .B1(fft_d[9]), 
        .C0(n9667), .Y(n9666) );
  CLKINVX1 U7903 ( .A(n9668), .Y(n9667) );
  AOI221XL U7904 ( .A0(fft_d[8]), .A1(n3090), .B0(fft_d[9]), .B1(n3080), .C0(
        n9669), .Y(n9668) );
  CLKINVX1 U7905 ( .A(n9670), .Y(n9669) );
  OAI221XL U7906 ( .A0(n3100), .A1(fft_d[7]), .B0(n3090), .B1(fft_d[8]), .C0(
        n9671), .Y(n9670) );
  CLKINVX1 U7907 ( .A(n9672), .Y(n9671) );
  AOI221XL U7908 ( .A0(fft_d[6]), .A1(n3110), .B0(fft_d[7]), .B1(n3100), .C0(
        n9673), .Y(n9672) );
  CLKINVX1 U7909 ( .A(n9674), .Y(n9673) );
  OAI221XL U7910 ( .A0(n3120), .A1(fft_d[5]), .B0(n3110), .B1(fft_d[6]), .C0(
        n9675), .Y(n9674) );
  CLKINVX1 U7911 ( .A(n9676), .Y(n9675) );
  AOI221XL U7912 ( .A0(fft_d[4]), .A1(n3130), .B0(fft_d[5]), .B1(n3120), .C0(
        n9677), .Y(n9676) );
  CLKINVX1 U7913 ( .A(n9678), .Y(n9677) );
  OAI221XL U7914 ( .A0(n3140), .A1(fft_d[3]), .B0(n3130), .B1(fft_d[4]), .C0(
        n9679), .Y(n9678) );
  CLKINVX1 U7915 ( .A(n9680), .Y(n9679) );
  AOI221XL U7916 ( .A0(fft_d[2]), .A1(n3150), .B0(fft_d[3]), .B1(n3140), .C0(
        n9681), .Y(n9680) );
  CLKINVX1 U7917 ( .A(n9682), .Y(n9681) );
  OAI221XL U7918 ( .A0(fft_d[1]), .A1(n9683), .B0(n3150), .B1(fft_d[2]), .C0(
        n9684), .Y(n9682) );
  AO21X1 U7919 ( .A0(n9683), .A1(fft_d[1]), .B0(n3160), .Y(n9684) );
  NOR2BX1 U7920 ( .AN(n2850), .B(n9616), .Y(n9683) );
  CLKINVX1 U7921 ( .A(fft_d[0]), .Y(n9616) );
  NOR2X1 U7922 ( .A(n10197), .B(n8856), .Y(N1080) );
  NOR2X1 U7923 ( .A(n10196), .B(n8856), .Y(N1079) );
  NOR2X1 U7924 ( .A(n10195), .B(n8856), .Y(N1078) );
  NOR2X1 U7925 ( .A(n10194), .B(n8855), .Y(N1077) );
  NOR2X1 U7926 ( .A(n10193), .B(n8855), .Y(N1076) );
  NOR2X1 U7927 ( .A(n10192), .B(n8855), .Y(N1075) );
  NOR2X1 U7928 ( .A(n10191), .B(n8855), .Y(N1074) );
  NOR2X1 U7929 ( .A(n10190), .B(n8855), .Y(N1073) );
  NOR2X1 U7930 ( .A(n10189), .B(n8855), .Y(N1072) );
  NOR2X1 U7931 ( .A(n10188), .B(n8855), .Y(N1071) );
  NOR2X1 U7932 ( .A(n10187), .B(n8855), .Y(N1070) );
  NOR2X1 U7933 ( .A(n10186), .B(n8855), .Y(N1069) );
  NOR2X1 U7934 ( .A(n10185), .B(n8855), .Y(N1068) );
  NOR2X1 U7935 ( .A(n10184), .B(n8855), .Y(N1067) );
  NOR2X1 U7936 ( .A(n10183), .B(n8855), .Y(N1066) );
  NOR2X1 U7937 ( .A(n10182), .B(n8855), .Y(N1065) );
  NOR2X1 U7938 ( .A(n10181), .B(n8854), .Y(N1064) );
  NOR2X1 U7939 ( .A(n10180), .B(n8854), .Y(N1063) );
  NOR2X1 U7940 ( .A(n10179), .B(n8854), .Y(N1062) );
  NOR2X1 U7941 ( .A(n10178), .B(n8854), .Y(N1061) );
  NOR2X1 U7942 ( .A(n10177), .B(n8854), .Y(N1060) );
  NOR2X1 U7943 ( .A(n10176), .B(n8854), .Y(N1059) );
  NOR2X1 U7944 ( .A(n10175), .B(n8854), .Y(N1058) );
  NOR2X1 U7945 ( .A(n10174), .B(n8854), .Y(N1057) );
  NOR2X1 U7946 ( .A(n10173), .B(n8854), .Y(N1056) );
  NOR2X1 U7947 ( .A(n10172), .B(n8854), .Y(N1055) );
  NOR2X1 U7948 ( .A(n10171), .B(n8854), .Y(N1054) );
  NOR2X1 U7949 ( .A(n10170), .B(n8854), .Y(N1053) );
  NOR2X1 U7950 ( .A(n10169), .B(n8854), .Y(N1052) );
  NOR2X1 U7951 ( .A(n10168), .B(n8853), .Y(N1051) );
  NOR2X1 U7952 ( .A(n10167), .B(n8853), .Y(N1050) );
  NOR2X1 U7953 ( .A(n10166), .B(n8853), .Y(N1049) );
  NOR2X1 U7954 ( .A(n9941), .B(n8853), .Y(N1048) );
  NOR2X1 U7955 ( .A(n9940), .B(n8853), .Y(N1047) );
  NOR2X1 U7956 ( .A(n9939), .B(n8853), .Y(N1046) );
  NOR2X1 U7957 ( .A(n9938), .B(n8853), .Y(N1045) );
  NOR2X1 U7958 ( .A(n9937), .B(n8853), .Y(N1044) );
  NOR2X1 U7959 ( .A(n9936), .B(n8853), .Y(N1043) );
  NOR2X1 U7960 ( .A(n9935), .B(n8853), .Y(N1042) );
  NOR2X1 U7961 ( .A(n9934), .B(n8853), .Y(N1041) );
  NOR2X1 U7962 ( .A(n9933), .B(n8853), .Y(N1040) );
  NOR2X1 U7963 ( .A(n9932), .B(n8853), .Y(N1039) );
  NOR2X1 U7964 ( .A(n9931), .B(n8852), .Y(N1038) );
  NOR2X1 U7965 ( .A(n9930), .B(n8852), .Y(N1037) );
  NOR2X1 U7966 ( .A(n9929), .B(n8852), .Y(N1036) );
  NOR2X1 U7967 ( .A(n9928), .B(n8852), .Y(N1035) );
  NOR2X1 U7968 ( .A(n9927), .B(n8852), .Y(N1034) );
  NOR2X1 U7969 ( .A(n9926), .B(n8852), .Y(N1033) );
  NOR2X1 U7970 ( .A(n9925), .B(n8852), .Y(N1032) );
  NOR2X1 U7971 ( .A(n9924), .B(n8852), .Y(N1031) );
  NOR2X1 U7972 ( .A(n9923), .B(n8852), .Y(N1030) );
  NOR2X1 U7973 ( .A(n9922), .B(n8852), .Y(N1029) );
  NOR2X1 U7974 ( .A(n9921), .B(n8852), .Y(N1028) );
  NOR2X1 U7975 ( .A(n9920), .B(n8852), .Y(N1027) );
  NOR2X1 U7976 ( .A(n9919), .B(n8852), .Y(N1026) );
  NOR2X1 U7977 ( .A(n9918), .B(n8851), .Y(N1025) );
  NOR2X1 U7978 ( .A(n9917), .B(n8851), .Y(N1024) );
  NOR2X1 U7979 ( .A(n9916), .B(n8851), .Y(N1023) );
  NOR2X1 U7980 ( .A(n9915), .B(n8851), .Y(N1022) );
  NOR2X1 U7981 ( .A(n9914), .B(n8851), .Y(N1021) );
  NOR2X1 U7982 ( .A(n9913), .B(n8851), .Y(N1020) );
  NOR2X1 U7983 ( .A(n9912), .B(n8851), .Y(N1019) );
  NOR2X1 U7984 ( .A(n9911), .B(n8851), .Y(N1018) );
  NOR2X1 U7985 ( .A(n9910), .B(n8851), .Y(N1017) );
  NOR2X1 U7986 ( .A(n10069), .B(n8851), .Y(N1016) );
  NOR2X1 U7987 ( .A(n10068), .B(n8851), .Y(N1015) );
  NOR2X1 U7988 ( .A(n10067), .B(n8851), .Y(N1014) );
  NOR2X1 U7989 ( .A(n10066), .B(n8851), .Y(N1013) );
  NOR2X1 U7990 ( .A(n10065), .B(n8850), .Y(N1012) );
  NOR2X1 U7991 ( .A(n10064), .B(n8850), .Y(N1011) );
  NOR2X1 U7992 ( .A(n10063), .B(n8850), .Y(N1010) );
  NOR2X1 U7993 ( .A(n10062), .B(n8850), .Y(N1009) );
  NOR2X1 U7994 ( .A(n10061), .B(n8850), .Y(N1008) );
  NOR2X1 U7995 ( .A(n10060), .B(n8850), .Y(N1007) );
  NOR2X1 U7996 ( .A(n10059), .B(n8850), .Y(N1006) );
  NOR2X1 U7997 ( .A(n10058), .B(n8850), .Y(N1005) );
  NOR2X1 U7998 ( .A(n10057), .B(n8850), .Y(N1004) );
  NOR2X1 U7999 ( .A(n10056), .B(n8850), .Y(N1003) );
  NOR2X1 U8000 ( .A(n10055), .B(n8850), .Y(N1002) );
  NOR2X1 U8001 ( .A(n10054), .B(n8850), .Y(N1001) );
  NOR2X1 U8002 ( .A(n10053), .B(n8850), .Y(N1000) );
  CLKINVX1 U8003 ( .A(n10478), .Y(n9580) );
  NOR3X1 U8004 ( .A(n9174), .B(n10476), .C(n6190), .Y(n10478) );
  NAND2X1 U8005 ( .A(n6072), .B(n9621), .Y(n9174) );
  NOR2X1 U8006 ( .A(counter[2]), .B(n9512), .Y(n9621) );
  NAND2X1 U8007 ( .A(n6075), .B(n6074), .Y(n9512) );
  SDFFRX2 fir_valid_reg ( .D(n6185), .SI(fft_valid), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(fir_valid), .QN(n10471) );
  SDFFRXL FIR_STATE_reg ( .D(n6186), .SI(n10472), .SE(test_se), .CK(clk), .RN(
        n9127), .Q(n10994), .QN(n10470) );
  SDFFRXL counter_reg_4_ ( .D(n6181), .SI(counter[3]), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(n6189), .QN(n6068) );
  SDFFRXL counter_reg_5_ ( .D(n6180), .SI(n6189), .SE(test_se), .CK(clk), .RN(
        n9127), .Q(n6191), .QN(n6067) );
  SDFFRXL BF2I_a_s_reg ( .D(counter[3]), .SI(n6215), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(n6192), .QN(n6078) );
  SDFFRXL BF2I_a07_r_reg_0_ ( .D(n4935), .SI(n10995), .SE(test_se), .CK(clk), 
        .RN(n9049), .Q(n6200), .QN(n10469) );
  SDFFRXL BF2I_a06_r_reg_0_ ( .D(n4934), .SI(n11011), .SE(test_se), .CK(clk), 
        .RN(n9049), .Q(n11010), .QN(n10468) );
  SDFFRXL BF2I_a05_r_reg_0_ ( .D(n4933), .SI(n11027), .SE(test_se), .CK(clk), 
        .RN(n9049), .Q(n11026), .QN(n10467) );
  SDFFRXL BF2I_a04_r_reg_0_ ( .D(n4932), .SI(n11043), .SE(test_se), .CK(clk), 
        .RN(n9049), .Q(n11042), .QN(n10466) );
  SDFFRXL BF2I_a03_r_reg_0_ ( .D(n4931), .SI(n11059), .SE(test_se), .CK(clk), 
        .RN(n9049), .Q(n11058), .QN(n10465) );
  SDFFRXL BF2I_a02_r_reg_0_ ( .D(n4930), .SI(n11075), .SE(test_se), .CK(clk), 
        .RN(n9049), .Q(n11074), .QN(n10464) );
  SDFFRXL BF2I_a01_r_reg_0_ ( .D(n4929), .SI(BF2I_a_xr_n[15]), .SE(test_se), 
        .CK(clk), .RN(n9049), .Q(n11090), .QN(n10463) );
  SDFFRXL BF2I_a07_r_reg_1_ ( .D(n4927), .SI(n6200), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n6201), .QN(n10462) );
  SDFFRXL BF2I_a06_r_reg_1_ ( .D(n4926), .SI(n11010), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11009), .QN(n10461) );
  SDFFRXL BF2I_a05_r_reg_1_ ( .D(n4925), .SI(n11026), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11025), .QN(n10460) );
  SDFFRXL BF2I_a04_r_reg_1_ ( .D(n4924), .SI(n11042), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11041), .QN(n10459) );
  SDFFRXL BF2I_a03_r_reg_1_ ( .D(n4923), .SI(n11058), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11057), .QN(n10458) );
  SDFFRXL BF2I_a02_r_reg_1_ ( .D(n4922), .SI(n11074), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11073), .QN(n10457) );
  SDFFRXL BF2I_a01_r_reg_1_ ( .D(n4921), .SI(n11090), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11089), .QN(n10456) );
  SDFFRXL BF2I_a07_r_reg_2_ ( .D(n4919), .SI(n6201), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(n6202), .QN(n10455) );
  SDFFRXL BF2I_a06_r_reg_2_ ( .D(n4918), .SI(n11009), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(n11008), .QN(n10454) );
  SDFFRXL BF2I_a05_r_reg_2_ ( .D(n4917), .SI(n11025), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11024), .QN(n10453) );
  SDFFRXL BF2I_a04_r_reg_2_ ( .D(n4916), .SI(n11041), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11040), .QN(n10452) );
  SDFFRXL BF2I_a03_r_reg_2_ ( .D(n4915), .SI(n11057), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11056), .QN(n10451) );
  SDFFRXL BF2I_a02_r_reg_2_ ( .D(n4914), .SI(n11073), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11072), .QN(n10450) );
  SDFFRXL BF2I_a01_r_reg_2_ ( .D(n4913), .SI(n11089), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11088), .QN(n10449) );
  SDFFRXL BF2I_a07_r_reg_3_ ( .D(n4911), .SI(n6202), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(n6203), .QN(n10448) );
  SDFFRXL BF2I_a06_r_reg_3_ ( .D(n4910), .SI(n11008), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(n11007), .QN(n10447) );
  SDFFRXL BF2I_a05_r_reg_3_ ( .D(n4909), .SI(n11024), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(n11023), .QN(n10446) );
  SDFFRXL BF2I_a04_r_reg_3_ ( .D(n4908), .SI(n11040), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(n11039), .QN(n10445) );
  SDFFRXL BF2I_a03_r_reg_3_ ( .D(n4907), .SI(n11056), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(n11055), .QN(n10444) );
  SDFFRXL BF2I_a02_r_reg_3_ ( .D(n4906), .SI(n11072), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(n11071), .QN(n10443) );
  SDFFRXL BF2I_a01_r_reg_3_ ( .D(n4905), .SI(n11088), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n11087), .QN(n10442) );
  SDFFRXL BF2I_a07_r_reg_4_ ( .D(n4903), .SI(n6203), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n6204), .QN(n10441) );
  SDFFRXL BF2I_a06_r_reg_4_ ( .D(n4902), .SI(n11007), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n11006), .QN(n10440) );
  SDFFRXL BF2I_a05_r_reg_4_ ( .D(n4901), .SI(n11023), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n11022), .QN(n10439) );
  SDFFRXL BF2I_a04_r_reg_4_ ( .D(n4900), .SI(n11039), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n11038), .QN(n10438) );
  SDFFRXL BF2I_a03_r_reg_4_ ( .D(n4899), .SI(n11055), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n11054), .QN(n10437) );
  SDFFRXL BF2I_a02_r_reg_4_ ( .D(n4898), .SI(n11071), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n11070), .QN(n10436) );
  SDFFRXL BF2I_a01_r_reg_4_ ( .D(n4897), .SI(n11087), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n11086), .QN(n10435) );
  SDFFRXL BF2I_a07_r_reg_5_ ( .D(n4895), .SI(n6204), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(n6205), .QN(n10434) );
  SDFFRXL BF2I_a06_r_reg_5_ ( .D(n4894), .SI(n11006), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11005), .QN(n10433) );
  SDFFRXL BF2I_a05_r_reg_5_ ( .D(n4893), .SI(n11022), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11021), .QN(n10432) );
  SDFFRXL BF2I_a04_r_reg_5_ ( .D(n4892), .SI(n11038), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11037), .QN(n10431) );
  SDFFRXL BF2I_a03_r_reg_5_ ( .D(n4891), .SI(n11054), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11053), .QN(n10430) );
  SDFFRXL BF2I_a02_r_reg_5_ ( .D(n4890), .SI(n11070), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11069), .QN(n10429) );
  SDFFRXL BF2I_a01_r_reg_5_ ( .D(n4889), .SI(n11086), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11085), .QN(n10428) );
  SDFFRXL BF2I_a07_r_reg_6_ ( .D(n4887), .SI(n6205), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(n6206), .QN(n10427) );
  SDFFRXL BF2I_a06_r_reg_6_ ( .D(n4886), .SI(n11005), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(n11004), .QN(n10426) );
  SDFFRXL BF2I_a05_r_reg_6_ ( .D(n4885), .SI(n11021), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(n11020), .QN(n10425) );
  SDFFRXL BF2I_a04_r_reg_6_ ( .D(n4884), .SI(n11037), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(n11036), .QN(n10424) );
  SDFFRXL BF2I_a03_r_reg_6_ ( .D(n4883), .SI(n11053), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(n11052), .QN(n10423) );
  SDFFRXL BF2I_a02_r_reg_6_ ( .D(n4882), .SI(n11069), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n11068), .QN(n10422) );
  SDFFRXL BF2I_a01_r_reg_6_ ( .D(n4881), .SI(n11085), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n11084), .QN(n10421) );
  SDFFRXL BF2I_a07_r_reg_7_ ( .D(n4879), .SI(n6206), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n6207), .QN(n10420) );
  SDFFRXL BF2I_a06_r_reg_7_ ( .D(n4878), .SI(n11004), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n11003), .QN(n10419) );
  SDFFRXL BF2I_a05_r_reg_7_ ( .D(n4877), .SI(n11020), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n11019), .QN(n10418) );
  SDFFRXL BF2I_a04_r_reg_7_ ( .D(n4876), .SI(n11036), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n11035), .QN(n10417) );
  SDFFRXL BF2I_a03_r_reg_7_ ( .D(n4875), .SI(n11052), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n11051), .QN(n10416) );
  SDFFRXL BF2I_a02_r_reg_7_ ( .D(n4874), .SI(n11068), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n11067), .QN(n10415) );
  SDFFRXL BF2I_a01_r_reg_7_ ( .D(n4873), .SI(n11084), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n11083), .QN(n10414) );
  SDFFRXL BF2I_a07_r_reg_8_ ( .D(n4871), .SI(n6207), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n6208), .QN(n10413) );
  SDFFRXL BF2I_a06_r_reg_8_ ( .D(n4870), .SI(n11003), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11002), .QN(n10412) );
  SDFFRXL BF2I_a05_r_reg_8_ ( .D(n4869), .SI(n11019), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11018), .QN(n10411) );
  SDFFRXL BF2I_a04_r_reg_8_ ( .D(n4868), .SI(n11035), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11034), .QN(n10410) );
  SDFFRXL BF2I_a03_r_reg_8_ ( .D(n4867), .SI(n11051), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11050), .QN(n10409) );
  SDFFRXL BF2I_a02_r_reg_8_ ( .D(n4866), .SI(n11067), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11066), .QN(n10408) );
  SDFFRXL BF2I_a01_r_reg_8_ ( .D(n4865), .SI(n11083), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11082), .QN(n10407) );
  SDFFRXL BF2I_a07_r_reg_9_ ( .D(n4863), .SI(n6208), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(n6209), .QN(n10406) );
  SDFFRXL BF2I_a06_r_reg_9_ ( .D(n4862), .SI(n11002), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(n11001), .QN(n10405) );
  SDFFRXL BF2I_a05_r_reg_9_ ( .D(n4861), .SI(n11018), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(n11017), .QN(n10404) );
  SDFFRXL BF2I_a04_r_reg_9_ ( .D(n4860), .SI(n11034), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(n11033), .QN(n10403) );
  SDFFRXL BF2I_a03_r_reg_9_ ( .D(n4859), .SI(n11050), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11049), .QN(n10402) );
  SDFFRXL BF2I_a02_r_reg_9_ ( .D(n4858), .SI(n11066), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11065), .QN(n10401) );
  SDFFRXL BF2I_a01_r_reg_9_ ( .D(n4857), .SI(n11082), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11081), .QN(n10400) );
  SDFFRXL BF2I_a07_r_reg_10_ ( .D(n4855), .SI(n6209), .SE(test_se), .CK(clk), 
        .RN(n9032), .Q(n6210), .QN(n10399) );
  SDFFRXL BF2I_a06_r_reg_10_ ( .D(n4854), .SI(n11001), .SE(test_se), .CK(clk), 
        .RN(n9032), .Q(n11000), .QN(n10398) );
  SDFFRXL BF2I_a05_r_reg_10_ ( .D(n4853), .SI(n11017), .SE(test_se), .CK(clk), 
        .RN(n9032), .Q(n11016), .QN(n10397) );
  SDFFRXL BF2I_a04_r_reg_10_ ( .D(n4852), .SI(n11033), .SE(test_se), .CK(clk), 
        .RN(n9032), .Q(n11032), .QN(n10396) );
  SDFFRXL BF2I_a03_r_reg_10_ ( .D(n4851), .SI(n11049), .SE(test_se), .CK(clk), 
        .RN(n9032), .Q(n11048), .QN(n10395) );
  SDFFRXL BF2I_a02_r_reg_10_ ( .D(n4850), .SI(n11065), .SE(test_se), .CK(clk), 
        .RN(n9032), .Q(n11064), .QN(n10394) );
  SDFFRXL BF2I_a01_r_reg_10_ ( .D(n4849), .SI(n11081), .SE(test_se), .CK(clk), 
        .RN(n9032), .Q(n11080), .QN(n10393) );
  SDFFRXL BF2I_a07_r_reg_11_ ( .D(n4847), .SI(n6210), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n6211), .QN(n10392) );
  SDFFRXL BF2I_a06_r_reg_11_ ( .D(n4846), .SI(n11000), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n10999), .QN(n10391) );
  SDFFRXL BF2I_a05_r_reg_11_ ( .D(n4845), .SI(n11016), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n11015), .QN(n10390) );
  SDFFRXL BF2I_a04_r_reg_11_ ( .D(n4844), .SI(n11032), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n11031), .QN(n10389) );
  SDFFRXL BF2I_a03_r_reg_11_ ( .D(n4843), .SI(n11048), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n11047), .QN(n10388) );
  SDFFRXL BF2I_a02_r_reg_11_ ( .D(n4842), .SI(n11064), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n11063), .QN(n10387) );
  SDFFRXL BF2I_a01_r_reg_11_ ( .D(n4841), .SI(n11080), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n11079), .QN(n10386) );
  SDFFRXL BF2I_a07_r_reg_12_ ( .D(n4839), .SI(n6211), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(n6212), .QN(n10385) );
  SDFFRXL BF2I_a06_r_reg_12_ ( .D(n4838), .SI(n10999), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(n10998), .QN(n10384) );
  SDFFRXL BF2I_a05_r_reg_12_ ( .D(n4837), .SI(n11015), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(n11014), .QN(n10383) );
  SDFFRXL BF2I_a04_r_reg_12_ ( .D(n4836), .SI(n11031), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11030), .QN(n10382) );
  SDFFRXL BF2I_a03_r_reg_12_ ( .D(n4835), .SI(n11047), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11046), .QN(n10381) );
  SDFFRXL BF2I_a02_r_reg_12_ ( .D(n4834), .SI(n11063), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11062), .QN(n10380) );
  SDFFRXL BF2I_a01_r_reg_12_ ( .D(n4833), .SI(n11079), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11078), .QN(n10379) );
  SDFFRXL BF2I_a07_r_reg_13_ ( .D(n4831), .SI(n6212), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n6213), .QN(n10378) );
  SDFFRXL BF2I_a06_r_reg_13_ ( .D(n4830), .SI(n10998), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n10997), .QN(n10377) );
  SDFFRXL BF2I_a05_r_reg_13_ ( .D(n4829), .SI(n11014), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n11013), .QN(n10376) );
  SDFFRXL BF2I_a04_r_reg_13_ ( .D(n4828), .SI(n11030), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n11029), .QN(n10375) );
  SDFFRXL BF2I_a03_r_reg_13_ ( .D(n4827), .SI(n11046), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n11045), .QN(n10374) );
  SDFFRXL BF2I_a02_r_reg_13_ ( .D(n4826), .SI(n11062), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n11061), .QN(n10373) );
  SDFFRXL BF2I_a01_r_reg_13_ ( .D(n4825), .SI(n11078), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n11077), .QN(n10372) );
  SDFFRXL BF2I_a07_r_reg_14_ ( .D(n4823), .SI(n6213), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n6214), .QN(n10371) );
  SDFFRXL BF2I_a06_r_reg_14_ ( .D(n4822), .SI(n10997), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n10996), .QN(n10370) );
  SDFFRXL BF2I_a05_r_reg_14_ ( .D(n4821), .SI(n11013), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n11012), .QN(n10369) );
  SDFFRXL BF2I_a04_r_reg_14_ ( .D(n4820), .SI(n11029), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n11028), .QN(n10368) );
  SDFFRXL BF2I_a03_r_reg_14_ ( .D(n4819), .SI(n11045), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n11044), .QN(n10367) );
  SDFFRXL BF2I_a02_r_reg_14_ ( .D(n4818), .SI(n11061), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n11060), .QN(n10366) );
  SDFFRXL BF2I_a01_r_reg_14_ ( .D(n4817), .SI(n11077), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n11076), .QN(n10365) );
  SDFFRXL BF2I_a07_r_reg_15_ ( .D(n4815), .SI(n6214), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(n6215), .QN(n10364) );
  SDFFRXL BF2I_a06_r_reg_15_ ( .D(n4814), .SI(n10996), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(n10995), .QN(n10363) );
  SDFFRXL BF2I_a05_r_reg_15_ ( .D(n4813), .SI(n11012), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11011), .QN(n10362) );
  SDFFRXL BF2I_a04_r_reg_15_ ( .D(n4812), .SI(n11028), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11027), .QN(n10361) );
  SDFFRXL BF2I_a03_r_reg_15_ ( .D(n4811), .SI(n11044), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11043), .QN(n10360) );
  SDFFRXL BF2I_a02_r_reg_15_ ( .D(n4810), .SI(n11060), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11059), .QN(n10359) );
  SDFFRXL BF2I_a01_r_reg_15_ ( .D(n4809), .SI(n11076), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11075), .QN(n10358) );
  SDFFRXL BF2II_a_s_reg ( .D(counter[2]), .SI(n11093), .SE(test_se), .CK(clk), 
        .RN(n9128), .Q(n11092), .QN(n10474) );
  SDFFRXL BF2II_a03_i_reg_0_ ( .D(n4807), .SI(n11125), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(n11124), .QN(n10357) );
  SDFFRXL BF2II_a02_i_reg_0_ ( .D(n4806), .SI(n11157), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(n11156), .QN(n10356) );
  SDFFRXL BF2II_a01_i_reg_0_ ( .D(n4805), .SI(N145), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(n11188), .QN(n10355) );
  SDFFRXL BF2II_a03_r_reg_0_ ( .D(n4803), .SI(n11109), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(n11108), .QN(n10354) );
  SDFFRXL BF2II_a02_r_reg_0_ ( .D(n4802), .SI(n11141), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(n11140), .QN(n10353) );
  SDFFRXL BF2II_a01_r_reg_0_ ( .D(n4801), .SI(n11173), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(n11172), .QN(n10352) );
  SDFFRXL BF2II_a03_r_reg_1_ ( .D(n4799), .SI(n11108), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11107), .QN(n10351) );
  SDFFRXL BF2II_a02_r_reg_1_ ( .D(n4798), .SI(n11140), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11139), .QN(n10350) );
  SDFFRXL BF2II_a01_r_reg_1_ ( .D(n4797), .SI(n11172), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(n11171), .QN(n10349) );
  SDFFRXL BF2II_a03_i_reg_1_ ( .D(n4795), .SI(n11124), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(n11123), .QN(n10348) );
  SDFFRXL BF2II_a02_i_reg_1_ ( .D(n4794), .SI(n11156), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(n11155), .QN(n10347) );
  SDFFRXL BF2II_a01_i_reg_1_ ( .D(n4793), .SI(n11188), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(n11187), .QN(n10346) );
  SDFFRXL BF2II_a03_r_reg_2_ ( .D(n4791), .SI(n11107), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11106), .QN(n10345) );
  SDFFRXL BF2II_a02_r_reg_2_ ( .D(n4790), .SI(n11139), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11138), .QN(n10344) );
  SDFFRXL BF2II_a01_r_reg_2_ ( .D(n4789), .SI(n11171), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11170), .QN(n10343) );
  SDFFRXL BF2II_a03_i_reg_2_ ( .D(n4787), .SI(n11123), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11122), .QN(n10342) );
  SDFFRXL BF2II_a02_i_reg_2_ ( .D(n4786), .SI(n11155), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11154), .QN(n10341) );
  SDFFRXL BF2II_a01_i_reg_2_ ( .D(n4785), .SI(n11187), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(n11186), .QN(n10340) );
  SDFFRXL BF2II_a03_r_reg_3_ ( .D(n4783), .SI(n11106), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n11105), .QN(n10339) );
  SDFFRXL BF2II_a02_r_reg_3_ ( .D(n4782), .SI(n11138), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n11137), .QN(n10338) );
  SDFFRXL BF2II_a01_r_reg_3_ ( .D(n4781), .SI(n11170), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n11169), .QN(n10337) );
  SDFFRXL BF2II_a03_i_reg_3_ ( .D(n4779), .SI(n11122), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n11121), .QN(n10336) );
  SDFFRXL BF2II_a02_i_reg_3_ ( .D(n4778), .SI(n11154), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n11153), .QN(n10335) );
  SDFFRXL BF2II_a01_i_reg_3_ ( .D(n4777), .SI(n11186), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n11185), .QN(n10334) );
  SDFFRXL BF2II_a03_r_reg_4_ ( .D(n4775), .SI(n11105), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n11104), .QN(n10333) );
  SDFFRXL BF2II_a02_r_reg_4_ ( .D(n4774), .SI(n11137), .SE(test_se), .CK(clk), 
        .RN(n9042), .Q(n11136), .QN(n10332) );
  SDFFRXL BF2II_a01_r_reg_4_ ( .D(n4773), .SI(n11169), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(n11168), .QN(n10331) );
  SDFFRXL BF2II_a03_i_reg_4_ ( .D(n4771), .SI(n11121), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(n11120), .QN(n10330) );
  SDFFRXL BF2II_a02_i_reg_4_ ( .D(n4770), .SI(n11153), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(n11152), .QN(n10329) );
  SDFFRXL BF2II_a01_i_reg_4_ ( .D(n4769), .SI(n11185), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(n11184), .QN(n10328) );
  SDFFRXL BF2II_a03_r_reg_5_ ( .D(n4767), .SI(n11104), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11103), .QN(n10327) );
  SDFFRXL BF2II_a02_r_reg_5_ ( .D(n4766), .SI(n11136), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11135), .QN(n10326) );
  SDFFRXL BF2II_a01_r_reg_5_ ( .D(n4765), .SI(n11168), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11167), .QN(n10325) );
  SDFFRXL BF2II_a03_i_reg_5_ ( .D(n4763), .SI(n11120), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11119), .QN(n10324) );
  SDFFRXL BF2II_a02_i_reg_5_ ( .D(n4762), .SI(n11152), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(n11151), .QN(n10323) );
  SDFFRXL BF2II_a01_i_reg_5_ ( .D(n4761), .SI(n11184), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(n11183), .QN(n10322) );
  SDFFRXL BF2II_a03_r_reg_6_ ( .D(n4759), .SI(n11103), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n11102), .QN(n10321) );
  SDFFRXL BF2II_a02_r_reg_6_ ( .D(n4758), .SI(n11135), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n11134), .QN(n10320) );
  SDFFRXL BF2II_a01_r_reg_6_ ( .D(n4757), .SI(n11167), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n11166), .QN(n10319) );
  SDFFRXL BF2II_a03_i_reg_6_ ( .D(n4755), .SI(n11119), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n11118), .QN(n10318) );
  SDFFRXL BF2II_a02_i_reg_6_ ( .D(n4754), .SI(n11151), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n11150), .QN(n10317) );
  SDFFRXL BF2II_a01_i_reg_6_ ( .D(n4753), .SI(n11183), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n11182), .QN(n10316) );
  SDFFRXL BF2II_a03_r_reg_7_ ( .D(n4751), .SI(n11102), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n11101), .QN(n10315) );
  SDFFRXL BF2II_a02_r_reg_7_ ( .D(n4750), .SI(n11134), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(n11133), .QN(n10314) );
  SDFFRXL BF2II_a01_r_reg_7_ ( .D(n4749), .SI(n11166), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(n11165), .QN(n10313) );
  SDFFRXL BF2II_a03_i_reg_7_ ( .D(n4747), .SI(n11118), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(n11117), .QN(n10312) );
  SDFFRXL BF2II_a02_i_reg_7_ ( .D(n4746), .SI(n11150), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(n11149), .QN(n10311) );
  SDFFRXL BF2II_a01_i_reg_7_ ( .D(n4745), .SI(n11182), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(n11181), .QN(n10310) );
  SDFFRXL BF2II_a03_r_reg_8_ ( .D(n4743), .SI(n11101), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11100), .QN(n10309) );
  SDFFRXL BF2II_a02_r_reg_8_ ( .D(n4742), .SI(n11133), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11132), .QN(n10308) );
  SDFFRXL BF2II_a01_r_reg_8_ ( .D(n4741), .SI(n11165), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11164), .QN(n10307) );
  SDFFRXL BF2II_a03_i_reg_8_ ( .D(n4739), .SI(n11117), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(n11116), .QN(n10306) );
  SDFFRXL BF2II_a02_i_reg_8_ ( .D(n4738), .SI(n11149), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(n11148), .QN(n10305) );
  SDFFRXL BF2II_a01_i_reg_8_ ( .D(n4737), .SI(n11181), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(n11180), .QN(n10304) );
  SDFFRXL BF2II_a03_r_reg_9_ ( .D(n4735), .SI(n11100), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11099), .QN(n10303) );
  SDFFRXL BF2II_a02_r_reg_9_ ( .D(n4734), .SI(n11132), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11131), .QN(n10302) );
  SDFFRXL BF2II_a01_r_reg_9_ ( .D(n4733), .SI(n11164), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11163), .QN(n10301) );
  SDFFRXL BF2II_a03_i_reg_9_ ( .D(n4731), .SI(n11116), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11115), .QN(n10300) );
  SDFFRXL BF2II_a02_i_reg_9_ ( .D(n4730), .SI(n11148), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11147), .QN(n10299) );
  SDFFRXL BF2II_a01_i_reg_9_ ( .D(n4729), .SI(n11180), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n11179), .QN(n10298) );
  SDFFRXL BF2II_a03_r_reg_10_ ( .D(n4727), .SI(n11099), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(n11098), .QN(n10297) );
  SDFFRXL BF2II_a02_r_reg_10_ ( .D(n4726), .SI(n11131), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(n11130), .QN(n10296) );
  SDFFRXL BF2II_a01_r_reg_10_ ( .D(n4725), .SI(n11163), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(n11162), .QN(n10295) );
  SDFFRXL BF2II_a03_i_reg_10_ ( .D(n4723), .SI(n11115), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(n11114), .QN(n10294) );
  SDFFRXL BF2II_a02_i_reg_10_ ( .D(n4722), .SI(n11147), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(n11146), .QN(n10293) );
  SDFFRXL BF2II_a01_i_reg_10_ ( .D(n4721), .SI(n11179), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(n11178), .QN(n10292) );
  SDFFRXL BF2II_a03_r_reg_11_ ( .D(n4719), .SI(n11098), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n11097), .QN(n10291) );
  SDFFRXL BF2II_a02_r_reg_11_ ( .D(n4718), .SI(n11130), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n11129), .QN(n10290) );
  SDFFRXL BF2II_a01_r_reg_11_ ( .D(n4717), .SI(n11162), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(n11161), .QN(n10289) );
  SDFFRXL BF2II_a03_i_reg_11_ ( .D(n4715), .SI(n11114), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(n11113), .QN(n10288) );
  SDFFRXL BF2II_a02_i_reg_11_ ( .D(n4714), .SI(n11146), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(n11145), .QN(n10287) );
  SDFFRXL BF2II_a01_i_reg_11_ ( .D(n4713), .SI(n11178), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(n11177), .QN(n10286) );
  SDFFRXL BF2II_a03_r_reg_12_ ( .D(n4711), .SI(n11097), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11096), .QN(n10285) );
  SDFFRXL BF2II_a02_r_reg_12_ ( .D(n4710), .SI(n11129), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11128), .QN(n10284) );
  SDFFRXL BF2II_a01_r_reg_12_ ( .D(n4709), .SI(n11161), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11160), .QN(n10283) );
  SDFFRXL BF2II_a03_i_reg_12_ ( .D(n4707), .SI(n11113), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11112), .QN(n10282) );
  SDFFRXL BF2II_a02_i_reg_12_ ( .D(n4706), .SI(n11145), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11144), .QN(n10281) );
  SDFFRXL BF2II_a01_i_reg_12_ ( .D(n4705), .SI(n11177), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(n11176), .QN(n10280) );
  SDFFRXL BF2II_a03_r_reg_13_ ( .D(n4703), .SI(n11096), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(n11095), .QN(n10279) );
  SDFFRXL BF2II_a02_r_reg_13_ ( .D(n4702), .SI(n11128), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(n11127), .QN(n10278) );
  SDFFRXL BF2II_a01_r_reg_13_ ( .D(n4701), .SI(n11160), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(n11159), .QN(n10277) );
  SDFFRXL BF2II_a03_i_reg_13_ ( .D(n4699), .SI(n11112), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(n11111), .QN(n10276) );
  SDFFRXL BF2II_a02_i_reg_13_ ( .D(n4698), .SI(n11144), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(n11143), .QN(n10275) );
  SDFFRXL BF2II_a01_i_reg_13_ ( .D(n4697), .SI(n11176), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(n11175), .QN(n10274) );
  SDFFRXL BF2II_a03_r_reg_14_ ( .D(n4695), .SI(n11095), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n11094), .QN(n10273) );
  SDFFRXL BF2II_a02_r_reg_14_ ( .D(n4694), .SI(n11127), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n11126), .QN(n10272) );
  SDFFRXL BF2II_a01_r_reg_14_ ( .D(n4693), .SI(n11159), .SE(test_se), .CK(clk), 
        .RN(n9025), .Q(n11158), .QN(n10271) );
  SDFFRXL BF2II_a03_i_reg_14_ ( .D(n4691), .SI(n11111), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(n11110), .QN(n10270) );
  SDFFRXL BF2II_a02_i_reg_14_ ( .D(n4690), .SI(n11143), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(n11142), .QN(n10269) );
  SDFFRXL BF2II_a01_i_reg_14_ ( .D(n4689), .SI(n11175), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(n11174), .QN(n10268) );
  SDFFRXL BF2II_a03_r_reg_15_ ( .D(n4687), .SI(n11094), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11093), .QN(n10267) );
  SDFFRXL BF2II_a02_r_reg_15_ ( .D(n4686), .SI(n11126), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11125), .QN(n10266) );
  SDFFRXL BF2II_a01_r_reg_15_ ( .D(n4685), .SI(n11158), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11157), .QN(n10265) );
  SDFFRXL BF2II_a03_i_reg_15_ ( .D(n4683), .SI(n11110), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11109), .QN(n10264) );
  SDFFRXL BF2II_a02_i_reg_15_ ( .D(n4682), .SI(n11142), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11141), .QN(n10263) );
  SDFFRXL BF2II_a01_i_reg_15_ ( .D(n4681), .SI(n11174), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(n11173), .QN(n10262) );
  SDFFRXL BF2I_b01_r_reg_0_ ( .D(n4679), .SI(n6279), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(n6216), .QN(n10261) );
  SDFFRXL BF2I_b01_r_reg_1_ ( .D(n4677), .SI(n6216), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(n6217), .QN(n10260) );
  SDFFRXL BF2I_b01_r_reg_2_ ( .D(n4675), .SI(n6217), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(n6218), .QN(n10259) );
  SDFFRXL BF2I_b01_r_reg_3_ ( .D(n4673), .SI(n6218), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n6219), .QN(n10258) );
  SDFFRXL BF2I_b01_r_reg_4_ ( .D(n4671), .SI(n6219), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(n6220), .QN(n10257) );
  SDFFRXL BF2I_b01_r_reg_5_ ( .D(n4669), .SI(n6220), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(n6221), .QN(n10256) );
  SDFFRXL BF2I_b01_r_reg_6_ ( .D(n4667), .SI(n6221), .SE(test_se), .CK(clk), 
        .RN(n9037), .Q(n6222), .QN(n10255) );
  SDFFRXL BF2I_b01_r_reg_7_ ( .D(n4665), .SI(n6222), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(n6223), .QN(n10254) );
  SDFFRXL BF2I_b01_r_reg_8_ ( .D(n4663), .SI(n6223), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(n6224), .QN(n10253) );
  SDFFRXL BF2I_b01_r_reg_9_ ( .D(n4661), .SI(n6224), .SE(test_se), .CK(clk), 
        .RN(n9032), .Q(n6225), .QN(n10252) );
  SDFFRXL BF2I_b01_r_reg_10_ ( .D(n4659), .SI(n6225), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(n6226), .QN(n10251) );
  SDFFRXL BF2I_b01_r_reg_11_ ( .D(n4657), .SI(n6226), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(n6227), .QN(n10250) );
  SDFFRXL BF2I_b01_r_reg_12_ ( .D(n4655), .SI(n6227), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n6228), .QN(n10249) );
  SDFFRXL BF2I_b01_r_reg_13_ ( .D(n4653), .SI(n6228), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(n6229), .QN(n10248) );
  SDFFRXL BF2I_b01_r_reg_14_ ( .D(n4651), .SI(n6229), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(n6230), .QN(n10247) );
  SDFFRXL BF2I_b01_r_reg_15_ ( .D(n4649), .SI(n6230), .SE(test_se), .CK(clk), 
        .RN(n9020), .Q(n6231), .QN(n10246) );
  SDFFRXL BF2I_b01_r_reg_16_ ( .D(n4647), .SI(n6231), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n6232), .QN(n10245) );
  SDFFRXL BF2I_b01_r_reg_17_ ( .D(n4645), .SI(n6232), .SE(test_se), .CK(clk), 
        .RN(n9014), .Q(n6233), .QN(n10244) );
  SDFFRXL BF2I_b01_r_reg_18_ ( .D(n4643), .SI(n6233), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(n6234), .QN(n10243) );
  SDFFRXL BF2I_b01_r_reg_19_ ( .D(n4641), .SI(n6234), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(n6235), .QN(n10242) );
  SDFFRXL BF2I_b01_r_reg_20_ ( .D(n4639), .SI(n6235), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(n6236), .QN(n10241) );
  SDFFRXL BF2I_b01_r_reg_21_ ( .D(n4637), .SI(n6236), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(n6237), .QN(n10240) );
  SDFFRXL BF2I_b01_r_reg_22_ ( .D(n4635), .SI(n6237), .SE(test_se), .CK(clk), 
        .RN(n8987), .Q(n6238), .QN(n10239) );
  SDFFRXL BF2I_b01_r_reg_23_ ( .D(n4633), .SI(n6238), .SE(test_se), .CK(clk), 
        .RN(n8987), .Q(n6239), .QN(n10238) );
  SDFFRXL BF2I_b01_r_reg_24_ ( .D(n4631), .SI(n6239), .SE(test_se), .CK(clk), 
        .RN(n8987), .Q(n6240), .QN(n10237) );
  SDFFRXL BF2I_b01_r_reg_25_ ( .D(n4629), .SI(n6240), .SE(test_se), .CK(clk), 
        .RN(n8987), .Q(n6241), .QN(n10236) );
  SDFFRXL BF2I_b01_r_reg_26_ ( .D(n4627), .SI(n6241), .SE(test_se), .CK(clk), 
        .RN(n8987), .Q(n6242), .QN(n10235) );
  SDFFRXL BF2I_b01_r_reg_27_ ( .D(n4625), .SI(n6242), .SE(test_se), .CK(clk), 
        .RN(n8987), .Q(n6243), .QN(n10234) );
  SDFFRXL BF2I_b01_r_reg_28_ ( .D(n4623), .SI(n6243), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(n6244), .QN(n10233) );
  SDFFRXL BF2I_b01_r_reg_29_ ( .D(n4621), .SI(n6244), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(n6245), .QN(n10232) );
  SDFFRXL BF2I_b01_r_reg_30_ ( .D(n4619), .SI(n6245), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(n6246), .QN(n10231) );
  SDFFRXL BF2I_b01_r_reg_31_ ( .D(n4617), .SI(n6246), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(n6247), .QN(n10230) );
  SDFFRXL BF2I_b01_i_reg_0_ ( .D(n4615), .SI(BF2I_b_xr_n[31]), .SE(test_se), 
        .CK(clk), .RN(n9048), .Q(n6248), .QN(n10229) );
  SDFFRXL BF2I_b01_i_reg_1_ ( .D(n4613), .SI(n6248), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(n6249), .QN(n10228) );
  SDFFRXL BF2I_b01_i_reg_2_ ( .D(n4611), .SI(n6249), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(n6250), .QN(n10227) );
  SDFFRXL BF2I_b01_i_reg_3_ ( .D(n4609), .SI(n6250), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(n6251), .QN(n10226) );
  SDFFRXL BF2I_b01_i_reg_4_ ( .D(n4607), .SI(n6251), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(n6252), .QN(n10225) );
  SDFFRXL BF2I_b01_i_reg_5_ ( .D(n4605), .SI(n6252), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(n6253), .QN(n10224) );
  SDFFRXL BF2I_b01_i_reg_6_ ( .D(n4603), .SI(n6253), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(n6254), .QN(n10223) );
  SDFFRXL BF2I_b01_i_reg_7_ ( .D(n4601), .SI(n6254), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(n6255), .QN(n10222) );
  SDFFRXL BF2I_b01_i_reg_8_ ( .D(n4599), .SI(n6255), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(n6256), .QN(n10221) );
  SDFFRXL BF2I_b01_i_reg_9_ ( .D(n4597), .SI(n6256), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(n6257), .QN(n10220) );
  SDFFRXL BF2I_b01_i_reg_10_ ( .D(n4595), .SI(n6257), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(n6258), .QN(n10219) );
  SDFFRXL BF2I_b01_i_reg_11_ ( .D(n4593), .SI(n6258), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(n6259), .QN(n10218) );
  SDFFRXL BF2I_b01_i_reg_12_ ( .D(n4591), .SI(n6259), .SE(test_se), .CK(clk), 
        .RN(n9027), .Q(n6260), .QN(n10217) );
  SDFFRXL BF2I_b01_i_reg_13_ ( .D(n4589), .SI(n6260), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(n6261), .QN(n10216) );
  SDFFRXL BF2I_b01_i_reg_14_ ( .D(n4587), .SI(n6261), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(n6262), .QN(n10215) );
  SDFFRXL BF2I_b01_i_reg_15_ ( .D(n4585), .SI(n6262), .SE(test_se), .CK(clk), 
        .RN(n9022), .Q(n6263), .QN(n10214) );
  SDFFRXL BF2I_b01_i_reg_16_ ( .D(n4583), .SI(n6263), .SE(test_se), .CK(clk), 
        .RN(n9022), .Q(n6264), .QN(n10213) );
  SDFFRXL BF2I_b01_i_reg_17_ ( .D(n4581), .SI(n6264), .SE(test_se), .CK(clk), 
        .RN(n9022), .Q(n6265), .QN(n10212) );
  SDFFRXL BF2I_b01_i_reg_18_ ( .D(n4579), .SI(n6265), .SE(test_se), .CK(clk), 
        .RN(n9022), .Q(n6266), .QN(n10211) );
  SDFFRXL BF2I_b01_i_reg_19_ ( .D(n4577), .SI(n6266), .SE(test_se), .CK(clk), 
        .RN(n9022), .Q(n6267), .QN(n10210) );
  SDFFRXL BF2I_b01_i_reg_20_ ( .D(n4575), .SI(n6267), .SE(test_se), .CK(clk), 
        .RN(n9022), .Q(n6268), .QN(n10209) );
  SDFFRXL BF2I_b01_i_reg_21_ ( .D(n4573), .SI(n6268), .SE(test_se), .CK(clk), 
        .RN(n9021), .Q(n6269), .QN(n10208) );
  SDFFRXL BF2I_b01_i_reg_22_ ( .D(n4571), .SI(n6269), .SE(test_se), .CK(clk), 
        .RN(n9021), .Q(n6270), .QN(n10207) );
  SDFFRXL BF2I_b01_i_reg_23_ ( .D(n4569), .SI(n6270), .SE(test_se), .CK(clk), 
        .RN(n9020), .Q(n6271), .QN(n10206) );
  SDFFRXL BF2I_b01_i_reg_24_ ( .D(n4567), .SI(n6271), .SE(test_se), .CK(clk), 
        .RN(n9020), .Q(n6272), .QN(n10205) );
  SDFFRXL BF2I_b01_i_reg_25_ ( .D(n4565), .SI(n6272), .SE(test_se), .CK(clk), 
        .RN(n9020), .Q(n6273), .QN(n10204) );
  SDFFRXL BF2I_b01_i_reg_26_ ( .D(n4563), .SI(n6273), .SE(test_se), .CK(clk), 
        .RN(n9020), .Q(n6274), .QN(n10203) );
  SDFFRXL BF2I_b01_i_reg_27_ ( .D(n4561), .SI(n6274), .SE(test_se), .CK(clk), 
        .RN(n9021), .Q(n6275), .QN(n10202) );
  SDFFRXL BF2I_b01_i_reg_28_ ( .D(n4559), .SI(n6275), .SE(test_se), .CK(clk), 
        .RN(n9021), .Q(n6276), .QN(n10201) );
  SDFFRXL BF2I_b01_i_reg_29_ ( .D(n4557), .SI(n6276), .SE(test_se), .CK(clk), 
        .RN(n9021), .Q(n6277), .QN(n10200) );
  SDFFRXL BF2I_b01_i_reg_30_ ( .D(n4555), .SI(n6277), .SE(test_se), .CK(clk), 
        .RN(n9021), .Q(n6278), .QN(n10199) );
  SDFFRXL BF2I_b01_i_reg_31_ ( .D(n4553), .SI(n6278), .SE(test_se), .CK(clk), 
        .RN(n9021), .Q(n6279), .QN(n10198) );
  SDFFRXL BF2II_b_s_reg ( .D(counter[0]), .SI(BF2II_b_xr_n[31]), .SE(test_se), 
        .CK(clk), .RN(n9128), .Q(n11091), .QN(n10473) );
  SDFFRXL fft_d7_q_reg_31_ ( .D(n4455), .SI(n10739), .SE(test_se), .CK(clk), 
        .RN(n8985), .Q(n10738), .QN(n10165) );
  SDFFRXL fft_d7_q_reg_30_ ( .D(n4454), .SI(n10740), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(n10739), .QN(n10164) );
  SDFFRXL fft_d7_q_reg_29_ ( .D(n4453), .SI(n10741), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(n10740), .QN(n10163) );
  SDFFRXL fft_d7_q_reg_28_ ( .D(n4452), .SI(n10742), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10741), .QN(n10162) );
  SDFFRXL fft_d7_q_reg_27_ ( .D(n4451), .SI(n10743), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10742), .QN(n10161) );
  SDFFRXL fft_d7_q_reg_26_ ( .D(n4450), .SI(n10744), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10743), .QN(n10160) );
  SDFFRXL fft_d7_q_reg_25_ ( .D(n4449), .SI(n10745), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10744), .QN(n10159) );
  SDFFRXL fft_d7_q_reg_24_ ( .D(n4448), .SI(n10746), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10745), .QN(n10158) );
  SDFFRXL fft_d7_q_reg_23_ ( .D(n4447), .SI(n10747), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(n10746), .QN(n10157) );
  SDFFRXL fft_d7_q_reg_22_ ( .D(n4446), .SI(n10748), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(n10747), .QN(n10156) );
  SDFFRXL fft_d7_q_reg_21_ ( .D(n4445), .SI(n10749), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(n10748), .QN(n10155) );
  SDFFRXL fft_d7_q_reg_20_ ( .D(n4444), .SI(n10750), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10749), .QN(n10154) );
  SDFFRXL fft_d7_q_reg_19_ ( .D(n4443), .SI(n10751), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10750), .QN(n10153) );
  SDFFRXL fft_d7_q_reg_18_ ( .D(n4442), .SI(n10752), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(n10751), .QN(n10152) );
  SDFFRXL fft_d7_q_reg_17_ ( .D(n4441), .SI(n10753), .SE(test_se), .CK(clk), 
        .RN(n9014), .Q(n10752), .QN(n10151) );
  SDFFRXL fft_d7_q_reg_16_ ( .D(n4440), .SI(n10754), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n10753), .QN(n10150) );
  SDFFRXL fft_d7_q_reg_15_ ( .D(n4439), .SI(n10755), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10754), .QN(n10149) );
  SDFFRXL fft_d7_q_reg_14_ ( .D(n4438), .SI(n10756), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(n10755), .QN(n10148) );
  SDFFRXL fft_d7_q_reg_13_ ( .D(n4437), .SI(n10757), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(n10756), .QN(n10147) );
  SDFFRXL fft_d7_q_reg_12_ ( .D(n4436), .SI(n10758), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(n10757), .QN(n10146) );
  SDFFRXL fft_d7_q_reg_11_ ( .D(n4435), .SI(n10759), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(n10758), .QN(n10145) );
  SDFFRXL fft_d7_q_reg_10_ ( .D(n4434), .SI(n10760), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(n10759), .QN(n10144) );
  SDFFRXL fft_d7_q_reg_9_ ( .D(n4433), .SI(n10761), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(n10760), .QN(n10143) );
  SDFFRXL fft_d7_q_reg_8_ ( .D(n4432), .SI(n10762), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(n10761), .QN(n10142) );
  SDFFRXL fft_d7_q_reg_7_ ( .D(n4431), .SI(n10763), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(n10762), .QN(n10141) );
  SDFFRXL fft_d7_q_reg_6_ ( .D(n4430), .SI(n10764), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10763), .QN(n10140) );
  SDFFRXL fft_d7_q_reg_5_ ( .D(n4429), .SI(n10765), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10764), .QN(n10139) );
  SDFFRXL fft_d7_q_reg_4_ ( .D(n4428), .SI(n10766), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(n10765), .QN(n10138) );
  SDFFRXL fft_d7_q_reg_3_ ( .D(n4427), .SI(n10767), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(n10766), .QN(n10137) );
  SDFFRXL fft_d7_q_reg_2_ ( .D(n4426), .SI(n10768), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10767), .QN(n10136) );
  SDFFRXL fft_d7_q_reg_1_ ( .D(n4425), .SI(n10769), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10768), .QN(n10135) );
  SDFFRXL fft_d7_q_reg_0_ ( .D(n4424), .SI(fft_d6[31]), .SE(test_se), .CK(clk), 
        .RN(n9017), .Q(n10769), .QN(n10134) );
  SDFFRXL fft_d11_q_reg_31_ ( .D(n4423), .SI(n10611), .SE(test_se), .CK(clk), 
        .RN(n8985), .Q(n10610), .QN(n10133) );
  SDFFRXL fft_d11_q_reg_30_ ( .D(n4422), .SI(n10612), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(n10611), .QN(n10132) );
  SDFFRXL fft_d11_q_reg_29_ ( .D(n4421), .SI(n10613), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(n10612), .QN(n10131) );
  SDFFRXL fft_d11_q_reg_28_ ( .D(n4420), .SI(n10614), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10613), .QN(n10130) );
  SDFFRXL fft_d11_q_reg_27_ ( .D(n4419), .SI(n10615), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10614), .QN(n10129) );
  SDFFRXL fft_d11_q_reg_26_ ( .D(n4418), .SI(n10616), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10615), .QN(n10128) );
  SDFFRXL fft_d11_q_reg_25_ ( .D(n4417), .SI(n10617), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10616), .QN(n10127) );
  SDFFRXL fft_d11_q_reg_24_ ( .D(n4416), .SI(n10618), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10617), .QN(n10126) );
  SDFFRXL fft_d11_q_reg_23_ ( .D(n4415), .SI(n10619), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10618), .QN(n10125) );
  SDFFRXL fft_d11_q_reg_22_ ( .D(n4414), .SI(n10620), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(n10619), .QN(n10124) );
  SDFFRXL fft_d11_q_reg_21_ ( .D(n4413), .SI(n10621), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(n10620), .QN(n10123) );
  SDFFRXL fft_d11_q_reg_20_ ( .D(n4412), .SI(n10622), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10621), .QN(n10122) );
  SDFFRXL fft_d11_q_reg_19_ ( .D(n4411), .SI(n10623), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10622), .QN(n10121) );
  SDFFRXL fft_d11_q_reg_18_ ( .D(n4410), .SI(n10624), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(n10623), .QN(n10120) );
  SDFFRXL fft_d11_q_reg_17_ ( .D(n4409), .SI(n10625), .SE(test_se), .CK(clk), 
        .RN(n9014), .Q(n10624), .QN(n10119) );
  SDFFRXL fft_d11_q_reg_16_ ( .D(n4408), .SI(n10626), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n10625), .QN(n10118) );
  SDFFRXL fft_d11_q_reg_15_ ( .D(n4407), .SI(n10627), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10626), .QN(n10117) );
  SDFFRXL fft_d11_q_reg_14_ ( .D(n4406), .SI(n10628), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10627), .QN(n10116) );
  SDFFRXL fft_d11_q_reg_13_ ( .D(n4405), .SI(n10629), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(n10628), .QN(n10115) );
  SDFFRXL fft_d11_q_reg_12_ ( .D(n4404), .SI(n10630), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(n10629), .QN(n10114) );
  SDFFRXL fft_d11_q_reg_11_ ( .D(n4403), .SI(n10631), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(n10630), .QN(n10113) );
  SDFFRXL fft_d11_q_reg_10_ ( .D(n4402), .SI(n10632), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(n10631), .QN(n10112) );
  SDFFRXL fft_d11_q_reg_9_ ( .D(n4401), .SI(n10633), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(n10632), .QN(n10111) );
  SDFFRXL fft_d11_q_reg_8_ ( .D(n4400), .SI(n10634), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(n10633), .QN(n101101) );
  SDFFRXL fft_d11_q_reg_7_ ( .D(n4399), .SI(n10635), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(n10634), .QN(n10109) );
  SDFFRXL fft_d11_q_reg_6_ ( .D(n4398), .SI(n10636), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10635), .QN(n10108) );
  SDFFRXL fft_d11_q_reg_5_ ( .D(n4397), .SI(n10637), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10636), .QN(n10107) );
  SDFFRXL fft_d11_q_reg_4_ ( .D(n4396), .SI(n10638), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(n10637), .QN(n10106) );
  SDFFRXL fft_d11_q_reg_3_ ( .D(n4395), .SI(n10639), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(n10638), .QN(n10105) );
  SDFFRXL fft_d11_q_reg_2_ ( .D(n4394), .SI(n10640), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10639), .QN(n10104) );
  SDFFRXL fft_d11_q_reg_1_ ( .D(n4393), .SI(n10641), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10640), .QN(n10103) );
  SDFFRXL fft_d11_q_reg_0_ ( .D(n4392), .SI(fft_d10[31]), .SE(test_se), .CK(
        clk), .RN(n9017), .Q(n10641), .QN(n10102) );
  SDFFRXL fft_d3_q_reg_31_ ( .D(n4391), .SI(n10867), .SE(test_se), .CK(clk), 
        .RN(n8985), .Q(n10866), .QN(n10101) );
  SDFFRXL fft_d3_q_reg_30_ ( .D(n4390), .SI(n10868), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(n10867), .QN(n10100) );
  SDFFRXL fft_d3_q_reg_29_ ( .D(n4389), .SI(n10869), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(n10868), .QN(n10099) );
  SDFFRXL fft_d3_q_reg_28_ ( .D(n4388), .SI(n10870), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10869), .QN(n10098) );
  SDFFRXL fft_d3_q_reg_27_ ( .D(n4387), .SI(n10871), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10870), .QN(n10097) );
  SDFFRXL fft_d3_q_reg_26_ ( .D(n4386), .SI(n10872), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10871), .QN(n10096) );
  SDFFRXL fft_d3_q_reg_25_ ( .D(n4385), .SI(n10873), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10872), .QN(n10095) );
  SDFFRXL fft_d3_q_reg_24_ ( .D(n4384), .SI(n10874), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10873), .QN(n10094) );
  SDFFRXL fft_d3_q_reg_23_ ( .D(n4383), .SI(n10875), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10874), .QN(n10093) );
  SDFFRXL fft_d3_q_reg_22_ ( .D(n4382), .SI(n10876), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10875), .QN(n10092) );
  SDFFRXL fft_d3_q_reg_21_ ( .D(n4381), .SI(n10877), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(n10876), .QN(n10091) );
  SDFFRXL fft_d3_q_reg_20_ ( .D(n4380), .SI(n10878), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10877), .QN(n10090) );
  SDFFRXL fft_d3_q_reg_19_ ( .D(n4379), .SI(n10879), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10878), .QN(n10089) );
  SDFFRXL fft_d3_q_reg_18_ ( .D(n4378), .SI(n10880), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10879), .QN(n10088) );
  SDFFRXL fft_d3_q_reg_17_ ( .D(n4377), .SI(n10881), .SE(test_se), .CK(clk), 
        .RN(n9014), .Q(n10880), .QN(n10087) );
  SDFFRXL fft_d3_q_reg_16_ ( .D(n4376), .SI(n10882), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n10881), .QN(n10086) );
  SDFFRXL fft_d3_q_reg_15_ ( .D(n4375), .SI(n10883), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10882), .QN(n10085) );
  SDFFRXL fft_d3_q_reg_14_ ( .D(n4374), .SI(n10884), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10883), .QN(n10084) );
  SDFFRXL fft_d3_q_reg_13_ ( .D(n4373), .SI(n10885), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10884), .QN(n10083) );
  SDFFRXL fft_d3_q_reg_12_ ( .D(n4372), .SI(n10886), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(n10885), .QN(n10082) );
  SDFFRXL fft_d3_q_reg_11_ ( .D(n4371), .SI(n10887), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(n10886), .QN(n10081) );
  SDFFRXL fft_d3_q_reg_10_ ( .D(n4370), .SI(n10888), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(n10887), .QN(n10080) );
  SDFFRXL fft_d3_q_reg_9_ ( .D(n4369), .SI(n10889), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(n10888), .QN(n10079) );
  SDFFRXL fft_d3_q_reg_8_ ( .D(n4368), .SI(n10890), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(n10889), .QN(n10078) );
  SDFFRXL fft_d3_q_reg_7_ ( .D(n4367), .SI(n10891), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(n10890), .QN(n10077) );
  SDFFRXL fft_d3_q_reg_6_ ( .D(n4366), .SI(n10892), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10891), .QN(n10076) );
  SDFFRXL fft_d3_q_reg_5_ ( .D(n4365), .SI(n10893), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10892), .QN(n10075) );
  SDFFRXL fft_d3_q_reg_4_ ( .D(n4364), .SI(n10894), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(n10893), .QN(n10074) );
  SDFFRXL fft_d3_q_reg_3_ ( .D(n4363), .SI(n10895), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(n10894), .QN(n10073) );
  SDFFRXL fft_d3_q_reg_2_ ( .D(n4362), .SI(n10896), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10895), .QN(n10072) );
  SDFFRXL fft_d3_q_reg_1_ ( .D(n4361), .SI(n10897), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10896), .QN(n10071) );
  SDFFRXL fft_d3_q_reg_0_ ( .D(n4360), .SI(fft_d2[31]), .SE(test_se), .CK(clk), 
        .RN(n9016), .Q(n10897), .QN(n10070) );
  SDFFRXL fft_d13_q_reg_31_ ( .D(n4359), .SI(n10547), .SE(test_se), .CK(clk), 
        .RN(n8985), .Q(n10546), .QN(n10069) );
  SDFFRXL fft_d13_q_reg_30_ ( .D(n4358), .SI(n10548), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(n10547), .QN(n10068) );
  SDFFRXL fft_d13_q_reg_29_ ( .D(n4357), .SI(n10549), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(n10548), .QN(n10067) );
  SDFFRXL fft_d13_q_reg_28_ ( .D(n4356), .SI(n10550), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10549), .QN(n10066) );
  SDFFRXL fft_d13_q_reg_27_ ( .D(n4355), .SI(n10551), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10550), .QN(n10065) );
  SDFFRXL fft_d13_q_reg_26_ ( .D(n4354), .SI(n10552), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10551), .QN(n10064) );
  SDFFRXL fft_d13_q_reg_25_ ( .D(n4353), .SI(n10553), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10552), .QN(n10063) );
  SDFFRXL fft_d13_q_reg_24_ ( .D(n4352), .SI(n10554), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10553), .QN(n10062) );
  SDFFRXL fft_d13_q_reg_23_ ( .D(n4351), .SI(n10555), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10554), .QN(n10061) );
  SDFFRXL fft_d13_q_reg_22_ ( .D(n4350), .SI(n10556), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10555), .QN(n10060) );
  SDFFRXL fft_d13_q_reg_21_ ( .D(n4349), .SI(n10557), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(n10556), .QN(n10059) );
  SDFFRXL fft_d13_q_reg_20_ ( .D(n4348), .SI(n10558), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10557), .QN(n10058) );
  SDFFRXL fft_d13_q_reg_19_ ( .D(n4347), .SI(n10559), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10558), .QN(n10057) );
  SDFFRXL fft_d13_q_reg_18_ ( .D(n4346), .SI(n10560), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10559), .QN(n10056) );
  SDFFRXL fft_d13_q_reg_17_ ( .D(n4345), .SI(n10561), .SE(test_se), .CK(clk), 
        .RN(n9014), .Q(n10560), .QN(n10055) );
  SDFFRXL fft_d13_q_reg_16_ ( .D(n4344), .SI(n10562), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n10561), .QN(n10054) );
  SDFFRXL fft_d13_q_reg_15_ ( .D(n4343), .SI(n10563), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10562), .QN(n10053) );
  SDFFRXL fft_d13_q_reg_14_ ( .D(n4342), .SI(n10564), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10563), .QN(n10052) );
  SDFFRXL fft_d13_q_reg_13_ ( .D(n4341), .SI(n10565), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10564), .QN(n10051) );
  SDFFRXL fft_d13_q_reg_12_ ( .D(n4340), .SI(n10566), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10565), .QN(n10050) );
  SDFFRXL fft_d13_q_reg_11_ ( .D(n4339), .SI(n10567), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(n10566), .QN(n10049) );
  SDFFRXL fft_d13_q_reg_10_ ( .D(n4338), .SI(n10568), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(n10567), .QN(n10048) );
  SDFFRXL fft_d13_q_reg_9_ ( .D(n4337), .SI(n10569), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(n10568), .QN(n10047) );
  SDFFRXL fft_d13_q_reg_8_ ( .D(n4336), .SI(n10570), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(n10569), .QN(n10046) );
  SDFFRXL fft_d13_q_reg_7_ ( .D(n4335), .SI(n10571), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(n10570), .QN(n10045) );
  SDFFRXL fft_d13_q_reg_6_ ( .D(n4334), .SI(n10572), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10571), .QN(n10044) );
  SDFFRXL fft_d13_q_reg_5_ ( .D(n4333), .SI(n10573), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10572), .QN(n10043) );
  SDFFRXL fft_d13_q_reg_4_ ( .D(n4332), .SI(n10574), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10573), .QN(n10042) );
  SDFFRXL fft_d13_q_reg_3_ ( .D(n4331), .SI(n10575), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(n10574), .QN(n10041) );
  SDFFRXL fft_d13_q_reg_2_ ( .D(n4330), .SI(n10576), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10575), .QN(n10040) );
  SDFFRXL fft_d13_q_reg_1_ ( .D(n4329), .SI(n10577), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10576), .QN(n10039) );
  SDFFRXL fft_d13_q_reg_0_ ( .D(n4328), .SI(fft_d12[31]), .SE(test_se), .CK(
        clk), .RN(n9016), .Q(n10577), .QN(n10038) );
  SDFFRXL fft_d5_q_reg_31_ ( .D(n4327), .SI(n10803), .SE(test_se), .CK(clk), 
        .RN(n8985), .Q(n10802), .QN(n10037) );
  SDFFRXL fft_d5_q_reg_30_ ( .D(n4326), .SI(n10804), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(n10803), .QN(n10036) );
  SDFFRXL fft_d5_q_reg_29_ ( .D(n4325), .SI(n10805), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(n10804), .QN(n10035) );
  SDFFRXL fft_d5_q_reg_28_ ( .D(n4324), .SI(n10806), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10805), .QN(n10034) );
  SDFFRXL fft_d5_q_reg_27_ ( .D(n4323), .SI(n10807), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10806), .QN(n10033) );
  SDFFRXL fft_d5_q_reg_26_ ( .D(n4322), .SI(n10808), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10807), .QN(n10032) );
  SDFFRXL fft_d5_q_reg_25_ ( .D(n4321), .SI(n10809), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10808), .QN(n10031) );
  SDFFRXL fft_d5_q_reg_24_ ( .D(n4320), .SI(n10810), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10809), .QN(n10030) );
  SDFFRXL fft_d5_q_reg_23_ ( .D(n4319), .SI(n10811), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10810), .QN(n10029) );
  SDFFRXL fft_d5_q_reg_22_ ( .D(n4318), .SI(n10812), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10811), .QN(n10028) );
  SDFFRXL fft_d5_q_reg_21_ ( .D(n4317), .SI(n10813), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(n10812), .QN(n10027) );
  SDFFRXL fft_d5_q_reg_20_ ( .D(n4316), .SI(n10814), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10813), .QN(n10026) );
  SDFFRXL fft_d5_q_reg_19_ ( .D(n4315), .SI(n10815), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10814), .QN(n10025) );
  SDFFRXL fft_d5_q_reg_18_ ( .D(n4314), .SI(n10816), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10815), .QN(n10024) );
  SDFFRXL fft_d5_q_reg_17_ ( .D(n4313), .SI(n10817), .SE(test_se), .CK(clk), 
        .RN(n9014), .Q(n10816), .QN(n10023) );
  SDFFRXL fft_d5_q_reg_16_ ( .D(n4312), .SI(n10818), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n10817), .QN(n10022) );
  SDFFRXL fft_d5_q_reg_15_ ( .D(n4311), .SI(n10819), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10818), .QN(n10021) );
  SDFFRXL fft_d5_q_reg_14_ ( .D(n4310), .SI(n10820), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10819), .QN(n10020) );
  SDFFRXL fft_d5_q_reg_13_ ( .D(n4309), .SI(n10821), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10820), .QN(n10019) );
  SDFFRXL fft_d5_q_reg_12_ ( .D(n4308), .SI(n10822), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10821), .QN(n10018) );
  SDFFRXL fft_d5_q_reg_11_ ( .D(n4307), .SI(n10823), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10822), .QN(n10017) );
  SDFFRXL fft_d5_q_reg_10_ ( .D(n4306), .SI(n10824), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(n10823), .QN(n10016) );
  SDFFRXL fft_d5_q_reg_9_ ( .D(n4305), .SI(n10825), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(n10824), .QN(n10015) );
  SDFFRXL fft_d5_q_reg_8_ ( .D(n4304), .SI(n10826), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(n10825), .QN(n10014) );
  SDFFRXL fft_d5_q_reg_7_ ( .D(n4303), .SI(n10827), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(n10826), .QN(n10013) );
  SDFFRXL fft_d5_q_reg_6_ ( .D(n4302), .SI(n10828), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10827), .QN(n10012) );
  SDFFRXL fft_d5_q_reg_5_ ( .D(n4301), .SI(n10829), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10828), .QN(n10011) );
  SDFFRXL fft_d5_q_reg_4_ ( .D(n4300), .SI(n10830), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10829), .QN(n10010) );
  SDFFRXL fft_d5_q_reg_3_ ( .D(n4299), .SI(n10831), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(n10830), .QN(n10009) );
  SDFFRXL fft_d5_q_reg_2_ ( .D(n4298), .SI(n10832), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10831), .QN(n10008) );
  SDFFRXL fft_d5_q_reg_1_ ( .D(n4297), .SI(n10833), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10832), .QN(n10007) );
  SDFFRXL fft_d5_q_reg_0_ ( .D(n4296), .SI(fft_d4[31]), .SE(test_se), .CK(clk), 
        .RN(n9016), .Q(n10833), .QN(n10006) );
  SDFFRXL fft_d9_q_reg_31_ ( .D(n4295), .SI(n10675), .SE(test_se), .CK(clk), 
        .RN(n8985), .Q(n10674), .QN(n10005) );
  SDFFRXL fft_d9_q_reg_30_ ( .D(n4294), .SI(n10676), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(n10675), .QN(n10004) );
  SDFFRXL fft_d9_q_reg_29_ ( .D(n4293), .SI(n10677), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(n10676), .QN(n10003) );
  SDFFRXL fft_d9_q_reg_28_ ( .D(n4292), .SI(n10678), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10677), .QN(n10002) );
  SDFFRXL fft_d9_q_reg_27_ ( .D(n4291), .SI(n10679), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10678), .QN(n10001) );
  SDFFRXL fft_d9_q_reg_26_ ( .D(n4290), .SI(n10680), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10679), .QN(n10000) );
  SDFFRXL fft_d9_q_reg_25_ ( .D(n4289), .SI(n10681), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10680), .QN(n9999) );
  SDFFRXL fft_d9_q_reg_24_ ( .D(n4288), .SI(n10682), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10681), .QN(n9998) );
  SDFFRXL fft_d9_q_reg_23_ ( .D(n4287), .SI(n10683), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10682), .QN(n9997) );
  SDFFRXL fft_d9_q_reg_22_ ( .D(n4286), .SI(n10684), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10683), .QN(n9996) );
  SDFFRXL fft_d9_q_reg_21_ ( .D(n4285), .SI(n10685), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(n10684), .QN(n9995) );
  SDFFRXL fft_d9_q_reg_20_ ( .D(n4284), .SI(n10686), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10685), .QN(n9994) );
  SDFFRXL fft_d9_q_reg_19_ ( .D(n4283), .SI(n10687), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10686), .QN(n9993) );
  SDFFRXL fft_d9_q_reg_18_ ( .D(n4282), .SI(n10688), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10687), .QN(n9992) );
  SDFFRXL fft_d9_q_reg_17_ ( .D(n4281), .SI(n10689), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10688), .QN(n9991) );
  SDFFRXL fft_d9_q_reg_16_ ( .D(n4280), .SI(n10690), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n10689), .QN(n9990) );
  SDFFRXL fft_d9_q_reg_15_ ( .D(n4279), .SI(n10691), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10690), .QN(n9989) );
  SDFFRXL fft_d9_q_reg_14_ ( .D(n4278), .SI(n10692), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10691), .QN(n9988) );
  SDFFRXL fft_d9_q_reg_13_ ( .D(n4277), .SI(n10693), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10692), .QN(n9987) );
  SDFFRXL fft_d9_q_reg_12_ ( .D(n4276), .SI(n10694), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10693), .QN(n9986) );
  SDFFRXL fft_d9_q_reg_11_ ( .D(n4275), .SI(n10695), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10694), .QN(n9985) );
  SDFFRXL fft_d9_q_reg_10_ ( .D(n4274), .SI(n10696), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10695), .QN(n9984) );
  SDFFRXL fft_d9_q_reg_9_ ( .D(n4273), .SI(n10697), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(n10696), .QN(n9983) );
  SDFFRXL fft_d9_q_reg_8_ ( .D(n4272), .SI(n10698), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(n10697), .QN(n9982) );
  SDFFRXL fft_d9_q_reg_7_ ( .D(n4271), .SI(n10699), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(n10698), .QN(n9981) );
  SDFFRXL fft_d9_q_reg_6_ ( .D(n4270), .SI(n10700), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10699), .QN(n9980) );
  SDFFRXL fft_d9_q_reg_5_ ( .D(n4269), .SI(n10701), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10700), .QN(n9979) );
  SDFFRXL fft_d9_q_reg_4_ ( .D(n4268), .SI(n10702), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10701), .QN(n9978) );
  SDFFRXL fft_d9_q_reg_3_ ( .D(n4267), .SI(n10703), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(n10702), .QN(n9977) );
  SDFFRXL fft_d9_q_reg_2_ ( .D(n4266), .SI(n10704), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10703), .QN(n9976) );
  SDFFRXL fft_d9_q_reg_1_ ( .D(n4265), .SI(n10705), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10704), .QN(n9975) );
  SDFFRXL fft_d9_q_reg_0_ ( .D(n4264), .SI(fft_d8[31]), .SE(test_se), .CK(clk), 
        .RN(n9016), .Q(n10705), .QN(n9974) );
  SDFFRXL fft_d1_q_reg_31_ ( .D(n4263), .SI(n10931), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10930), .QN(n9973) );
  SDFFRXL fft_d1_q_reg_30_ ( .D(n4262), .SI(n10932), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(n10931), .QN(n9972) );
  SDFFRXL fft_d1_q_reg_29_ ( .D(n4261), .SI(n10933), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(n10932), .QN(n9971) );
  SDFFRXL fft_d1_q_reg_28_ ( .D(n4260), .SI(n10934), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10933), .QN(n9970) );
  SDFFRXL fft_d1_q_reg_27_ ( .D(n4259), .SI(n10935), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10934), .QN(n9969) );
  SDFFRXL fft_d1_q_reg_26_ ( .D(n4258), .SI(n10936), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10935), .QN(n9968) );
  SDFFRXL fft_d1_q_reg_25_ ( .D(n4257), .SI(n10937), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10936), .QN(n9967) );
  SDFFRXL fft_d1_q_reg_24_ ( .D(n4256), .SI(n10938), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10937), .QN(n9966) );
  SDFFRXL fft_d1_q_reg_23_ ( .D(n4255), .SI(n10939), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10938), .QN(n9965) );
  SDFFRXL fft_d1_q_reg_22_ ( .D(n4254), .SI(n10940), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10939), .QN(n9964) );
  SDFFRXL fft_d1_q_reg_21_ ( .D(n4253), .SI(n10941), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10940), .QN(n9963) );
  SDFFRXL fft_d1_q_reg_20_ ( .D(n4252), .SI(n10942), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10941), .QN(n9962) );
  SDFFRXL fft_d1_q_reg_19_ ( .D(n4251), .SI(n10943), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10942), .QN(n9961) );
  SDFFRXL fft_d1_q_reg_18_ ( .D(n4250), .SI(n10944), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10943), .QN(n9960) );
  SDFFRXL fft_d1_q_reg_17_ ( .D(n4249), .SI(n10945), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10944), .QN(n9959) );
  SDFFRXL fft_d1_q_reg_16_ ( .D(n4248), .SI(n10946), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n10945), .QN(n9958) );
  SDFFRXL fft_d1_q_reg_15_ ( .D(n4247), .SI(n10947), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10946), .QN(n9957) );
  SDFFRXL fft_d1_q_reg_14_ ( .D(n4246), .SI(n10948), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10947), .QN(n9956) );
  SDFFRXL fft_d1_q_reg_13_ ( .D(n4245), .SI(n10949), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10948), .QN(n9955) );
  SDFFRXL fft_d1_q_reg_12_ ( .D(n4244), .SI(n10950), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10949), .QN(n9954) );
  SDFFRXL fft_d1_q_reg_11_ ( .D(n4243), .SI(n10951), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10950), .QN(n9953) );
  SDFFRXL fft_d1_q_reg_10_ ( .D(n4242), .SI(n10952), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10951), .QN(n9952) );
  SDFFRXL fft_d1_q_reg_9_ ( .D(n4241), .SI(n10953), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10952), .QN(n9951) );
  SDFFRXL fft_d1_q_reg_8_ ( .D(n4240), .SI(n10954), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(n10953), .QN(n9950) );
  SDFFRXL fft_d1_q_reg_7_ ( .D(n4239), .SI(n10955), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(n10954), .QN(n9949) );
  SDFFRXL fft_d1_q_reg_6_ ( .D(n4238), .SI(n10956), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10955), .QN(n9948) );
  SDFFRXL fft_d1_q_reg_5_ ( .D(n4237), .SI(n10957), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10956), .QN(n9947) );
  SDFFRXL fft_d1_q_reg_4_ ( .D(n4236), .SI(n10958), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10957), .QN(n9946) );
  SDFFRXL fft_d1_q_reg_3_ ( .D(n4235), .SI(n10959), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10958), .QN(n9945) );
  SDFFRXL fft_d1_q_reg_2_ ( .D(n4234), .SI(n10960), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10959), .QN(n9944) );
  SDFFRXL fft_d1_q_reg_1_ ( .D(n4233), .SI(n10961), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10960), .QN(n9943) );
  SDFFRXL fft_d1_q_reg_0_ ( .D(n4232), .SI(fft_d0[31]), .SE(test_se), .CK(clk), 
        .RN(n9016), .Q(n10961), .QN(n9942) );
  SDFFRXL fft_d14_q_reg_31_ ( .D(n4231), .SI(n10515), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10514), .QN(n9941) );
  SDFFRXL fft_d14_q_reg_30_ ( .D(n4230), .SI(n10516), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(n10515), .QN(n9940) );
  SDFFRXL fft_d14_q_reg_29_ ( .D(n4229), .SI(n10517), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(n10516), .QN(n9939) );
  SDFFRXL fft_d14_q_reg_28_ ( .D(n4228), .SI(n10518), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10517), .QN(n9938) );
  SDFFRXL fft_d14_q_reg_27_ ( .D(n4227), .SI(n10519), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10518), .QN(n9937) );
  SDFFRXL fft_d14_q_reg_26_ ( .D(n4226), .SI(n10520), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10519), .QN(n9936) );
  SDFFRXL fft_d14_q_reg_25_ ( .D(n4225), .SI(n10521), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10520), .QN(n9935) );
  SDFFRXL fft_d14_q_reg_24_ ( .D(n4224), .SI(n10522), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10521), .QN(n9934) );
  SDFFRXL fft_d14_q_reg_23_ ( .D(n4223), .SI(n10523), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10522), .QN(n9933) );
  SDFFRXL fft_d14_q_reg_22_ ( .D(n4222), .SI(n10524), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10523), .QN(n9932) );
  SDFFRXL fft_d14_q_reg_21_ ( .D(n4221), .SI(n10525), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10524), .QN(n9931) );
  SDFFRXL fft_d14_q_reg_20_ ( .D(n4220), .SI(n10526), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10525), .QN(n9930) );
  SDFFRXL fft_d14_q_reg_19_ ( .D(n4219), .SI(n10527), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10526), .QN(n9929) );
  SDFFRXL fft_d14_q_reg_18_ ( .D(n4218), .SI(n10528), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10527), .QN(n9928) );
  SDFFRXL fft_d14_q_reg_17_ ( .D(n4217), .SI(n10529), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10528), .QN(n9927) );
  SDFFRXL fft_d14_q_reg_16_ ( .D(n4216), .SI(n10530), .SE(test_se), .CK(clk), 
        .RN(n9019), .Q(n10529), .QN(n9926) );
  SDFFRXL fft_d14_q_reg_15_ ( .D(n4215), .SI(n10531), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10530), .QN(n9925) );
  SDFFRXL fft_d14_q_reg_14_ ( .D(n4214), .SI(n10532), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10531), .QN(n9924) );
  SDFFRXL fft_d14_q_reg_13_ ( .D(n4213), .SI(n10533), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10532), .QN(n9923) );
  SDFFRXL fft_d14_q_reg_12_ ( .D(n4212), .SI(n10534), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10533), .QN(n9922) );
  SDFFRXL fft_d14_q_reg_11_ ( .D(n4211), .SI(n10535), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10534), .QN(n9921) );
  SDFFRXL fft_d14_q_reg_10_ ( .D(n4210), .SI(n10536), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10535), .QN(n9920) );
  SDFFRXL fft_d14_q_reg_9_ ( .D(n4209), .SI(n10537), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10536), .QN(n9919) );
  SDFFRXL fft_d14_q_reg_8_ ( .D(n4208), .SI(n10538), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(n10537), .QN(n9918) );
  SDFFRXL fft_d14_q_reg_7_ ( .D(n4207), .SI(n10539), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(n10538), .QN(n9917) );
  SDFFRXL fft_d14_q_reg_6_ ( .D(n4206), .SI(n10540), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10539), .QN(n9916) );
  SDFFRXL fft_d14_q_reg_5_ ( .D(n4205), .SI(n10541), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10540), .QN(n9915) );
  SDFFRXL fft_d14_q_reg_4_ ( .D(n4204), .SI(n10542), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10541), .QN(n9914) );
  SDFFRXL fft_d14_q_reg_3_ ( .D(n4203), .SI(n10543), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10542), .QN(n9913) );
  SDFFRXL fft_d14_q_reg_2_ ( .D(n4202), .SI(n10544), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10543), .QN(n9912) );
  SDFFRXL fft_d14_q_reg_1_ ( .D(n4201), .SI(n10545), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10544), .QN(n9911) );
  SDFFRXL fft_d14_q_reg_0_ ( .D(n4200), .SI(fft_d13[31]), .SE(test_se), .CK(
        clk), .RN(n9016), .Q(n10545), .QN(n9910) );
  SDFFRXL fft_d6_q_reg_31_ ( .D(n4199), .SI(n10771), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10770), .QN(n9909) );
  SDFFRXL fft_d6_q_reg_30_ ( .D(n4198), .SI(n10772), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(n10771), .QN(n9908) );
  SDFFRXL fft_d6_q_reg_29_ ( .D(n4197), .SI(n10773), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(n10772), .QN(n9907) );
  SDFFRXL fft_d6_q_reg_28_ ( .D(n4196), .SI(n10774), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(n10773), .QN(n9906) );
  SDFFRXL fft_d6_q_reg_27_ ( .D(n4195), .SI(n10775), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10774), .QN(n9905) );
  SDFFRXL fft_d6_q_reg_26_ ( .D(n4194), .SI(n10776), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10775), .QN(n9904) );
  SDFFRXL fft_d6_q_reg_25_ ( .D(n4193), .SI(n10777), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10776), .QN(n9903) );
  SDFFRXL fft_d6_q_reg_24_ ( .D(n4192), .SI(n10778), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10777), .QN(n9902) );
  SDFFRXL fft_d6_q_reg_23_ ( .D(n4191), .SI(n10779), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10778), .QN(n9901) );
  SDFFRXL fft_d6_q_reg_22_ ( .D(n4190), .SI(n10780), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10779), .QN(n9900) );
  SDFFRXL fft_d6_q_reg_21_ ( .D(n4189), .SI(n10781), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10780), .QN(n9899) );
  SDFFRXL fft_d6_q_reg_20_ ( .D(n4188), .SI(n10782), .SE(test_se), .CK(clk), 
        .RN(n8998), .Q(n10781), .QN(n9898) );
  SDFFRXL fft_d6_q_reg_19_ ( .D(n4187), .SI(n10783), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10782), .QN(n9897) );
  SDFFRXL fft_d6_q_reg_18_ ( .D(n4186), .SI(n10784), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10783), .QN(n9896) );
  SDFFRXL fft_d6_q_reg_17_ ( .D(n4185), .SI(n10785), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10784), .QN(n9895) );
  SDFFRXL fft_d6_q_reg_16_ ( .D(n4184), .SI(n10786), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(n10785), .QN(n9894) );
  SDFFRXL fft_d6_q_reg_15_ ( .D(n4183), .SI(n10787), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10786), .QN(n9893) );
  SDFFRXL fft_d6_q_reg_14_ ( .D(n4182), .SI(n10788), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10787), .QN(n9892) );
  SDFFRXL fft_d6_q_reg_13_ ( .D(n4181), .SI(n10789), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10788), .QN(n9891) );
  SDFFRXL fft_d6_q_reg_12_ ( .D(n4180), .SI(n10790), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10789), .QN(n9890) );
  SDFFRXL fft_d6_q_reg_11_ ( .D(n4179), .SI(n10791), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10790), .QN(n9889) );
  SDFFRXL fft_d6_q_reg_10_ ( .D(n4178), .SI(n10792), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10791), .QN(n9888) );
  SDFFRXL fft_d6_q_reg_9_ ( .D(n4177), .SI(n10793), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10792), .QN(n9887) );
  SDFFRXL fft_d6_q_reg_8_ ( .D(n4176), .SI(n10794), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(n10793), .QN(n9886) );
  SDFFRXL fft_d6_q_reg_7_ ( .D(n4175), .SI(n10795), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(n10794), .QN(n9885) );
  SDFFRXL fft_d6_q_reg_6_ ( .D(n4174), .SI(n10796), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(n10795), .QN(n9884) );
  SDFFRXL fft_d6_q_reg_5_ ( .D(n4173), .SI(n10797), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10796), .QN(n9883) );
  SDFFRXL fft_d6_q_reg_4_ ( .D(n4172), .SI(n10798), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10797), .QN(n9882) );
  SDFFRXL fft_d6_q_reg_3_ ( .D(n4171), .SI(n10799), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10798), .QN(n9881) );
  SDFFRXL fft_d6_q_reg_2_ ( .D(n4170), .SI(n10800), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(n10799), .QN(n9880) );
  SDFFRXL fft_d6_q_reg_1_ ( .D(n4169), .SI(n10801), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10800), .QN(n9879) );
  SDFFRXL fft_d6_q_reg_0_ ( .D(n4168), .SI(fft_d5[31]), .SE(test_se), .CK(clk), 
        .RN(n9016), .Q(n10801), .QN(n9878) );
  SDFFRXL fft_d10_q_reg_31_ ( .D(n4167), .SI(n10643), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10642), .QN(n9877) );
  SDFFRXL fft_d10_q_reg_30_ ( .D(n4166), .SI(n10644), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(n10643), .QN(n9876) );
  SDFFRXL fft_d10_q_reg_29_ ( .D(n4165), .SI(n10645), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(n10644), .QN(n9875) );
  SDFFRXL fft_d10_q_reg_28_ ( .D(n4164), .SI(n10646), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(n10645), .QN(n9874) );
  SDFFRXL fft_d10_q_reg_27_ ( .D(n4163), .SI(n10647), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(n10646), .QN(n9873) );
  SDFFRXL fft_d10_q_reg_26_ ( .D(n4162), .SI(n10648), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10647), .QN(n9872) );
  SDFFRXL fft_d10_q_reg_25_ ( .D(n4161), .SI(n10649), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10648), .QN(n9871) );
  SDFFRXL fft_d10_q_reg_24_ ( .D(n4160), .SI(n10650), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10649), .QN(n9870) );
  SDFFRXL fft_d10_q_reg_23_ ( .D(n4159), .SI(n10651), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10650), .QN(n9869) );
  SDFFRXL fft_d10_q_reg_22_ ( .D(n4158), .SI(n10652), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10651), .QN(n9868) );
  SDFFRXL fft_d10_q_reg_21_ ( .D(n4157), .SI(n10653), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10652), .QN(n9867) );
  SDFFRXL fft_d10_q_reg_20_ ( .D(n4156), .SI(n10654), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(n10653), .QN(n9866) );
  SDFFRXL fft_d10_q_reg_19_ ( .D(n4155), .SI(n10655), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10654), .QN(n9865) );
  SDFFRXL fft_d10_q_reg_18_ ( .D(n4154), .SI(n10656), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10655), .QN(n9864) );
  SDFFRXL fft_d10_q_reg_17_ ( .D(n4153), .SI(n10657), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10656), .QN(n9863) );
  SDFFRXL fft_d10_q_reg_16_ ( .D(n4152), .SI(n10658), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(n10657), .QN(n9862) );
  SDFFRXL fft_d10_q_reg_15_ ( .D(n4151), .SI(n10659), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10658), .QN(n9861) );
  SDFFRXL fft_d10_q_reg_14_ ( .D(n4150), .SI(n10660), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10659), .QN(n9860) );
  SDFFRXL fft_d10_q_reg_13_ ( .D(n4149), .SI(n10661), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10660), .QN(n9859) );
  SDFFRXL fft_d10_q_reg_12_ ( .D(n4148), .SI(n10662), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10661), .QN(n9858) );
  SDFFRXL fft_d10_q_reg_11_ ( .D(n4147), .SI(n10663), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10662), .QN(n9857) );
  SDFFRXL fft_d10_q_reg_10_ ( .D(n4146), .SI(n10664), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10663), .QN(n9856) );
  SDFFRXL fft_d10_q_reg_9_ ( .D(n4145), .SI(n10665), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10664), .QN(n9855) );
  SDFFRXL fft_d10_q_reg_8_ ( .D(n4144), .SI(n10666), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(n10665), .QN(n9854) );
  SDFFRXL fft_d10_q_reg_7_ ( .D(n4143), .SI(n10667), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(n10666), .QN(n9853) );
  SDFFRXL fft_d10_q_reg_6_ ( .D(n4142), .SI(n10668), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(n10667), .QN(n9852) );
  SDFFRXL fft_d10_q_reg_5_ ( .D(n4141), .SI(n10669), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10668), .QN(n9851) );
  SDFFRXL fft_d10_q_reg_4_ ( .D(n4140), .SI(n10670), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10669), .QN(n9850) );
  SDFFRXL fft_d10_q_reg_3_ ( .D(n4139), .SI(n10671), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10670), .QN(n9849) );
  SDFFRXL fft_d10_q_reg_2_ ( .D(n4138), .SI(n10672), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(n10671), .QN(n9848) );
  SDFFRXL fft_d10_q_reg_1_ ( .D(n4137), .SI(n10673), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10672), .QN(n9847) );
  SDFFRXL fft_d10_q_reg_0_ ( .D(n4136), .SI(fft_d9[31]), .SE(test_se), .CK(clk), .RN(n9016), .Q(n10673), .QN(n9846) );
  SDFFRXL fft_d2_q_reg_31_ ( .D(n4135), .SI(n10899), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10898), .QN(n9845) );
  SDFFRXL fft_d2_q_reg_30_ ( .D(n4134), .SI(n10900), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(n10899), .QN(n9844) );
  SDFFRXL fft_d2_q_reg_29_ ( .D(n4133), .SI(n10901), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(n10900), .QN(n9843) );
  SDFFRXL fft_d2_q_reg_28_ ( .D(n4132), .SI(n10902), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(n10901), .QN(n9842) );
  SDFFRXL fft_d2_q_reg_27_ ( .D(n4131), .SI(n10903), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(n10902), .QN(n9841) );
  SDFFRXL fft_d2_q_reg_26_ ( .D(n4130), .SI(n10904), .SE(test_se), .CK(clk), 
        .RN(n8960), .Q(n10903), .QN(n9840) );
  SDFFRXL fft_d2_q_reg_25_ ( .D(n4129), .SI(n10905), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10904), .QN(n9839) );
  SDFFRXL fft_d2_q_reg_24_ ( .D(n4128), .SI(n10906), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10905), .QN(n9838) );
  SDFFRXL fft_d2_q_reg_23_ ( .D(n4127), .SI(n10907), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10906), .QN(n9837) );
  SDFFRXL fft_d2_q_reg_22_ ( .D(n4126), .SI(n10908), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10907), .QN(n9836) );
  SDFFRXL fft_d2_q_reg_21_ ( .D(n4125), .SI(n10909), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10908), .QN(n9835) );
  SDFFRXL fft_d2_q_reg_20_ ( .D(n4124), .SI(n10910), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(n10909), .QN(n9834) );
  SDFFRXL fft_d2_q_reg_19_ ( .D(n4123), .SI(n10911), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10910), .QN(n9833) );
  SDFFRXL fft_d2_q_reg_18_ ( .D(n4122), .SI(n10912), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10911), .QN(n9832) );
  SDFFRXL fft_d2_q_reg_17_ ( .D(n4121), .SI(n10913), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10912), .QN(n9831) );
  SDFFRXL fft_d2_q_reg_16_ ( .D(n4120), .SI(n10914), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(n10913), .QN(n9830) );
  SDFFRXL fft_d2_q_reg_15_ ( .D(n4119), .SI(n10915), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10914), .QN(n9829) );
  SDFFRXL fft_d2_q_reg_14_ ( .D(n4118), .SI(n10916), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10915), .QN(n9828) );
  SDFFRXL fft_d2_q_reg_13_ ( .D(n4117), .SI(n10917), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10916), .QN(n9827) );
  SDFFRXL fft_d2_q_reg_12_ ( .D(n4116), .SI(n10918), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10917), .QN(n9826) );
  SDFFRXL fft_d2_q_reg_11_ ( .D(n4115), .SI(n10919), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10918), .QN(n9825) );
  SDFFRXL fft_d2_q_reg_10_ ( .D(n4114), .SI(n10920), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10919), .QN(n9824) );
  SDFFRXL fft_d2_q_reg_9_ ( .D(n4113), .SI(n10921), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10920), .QN(n9823) );
  SDFFRXL fft_d2_q_reg_8_ ( .D(n4112), .SI(n10922), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(n10921), .QN(n9822) );
  SDFFRXL fft_d2_q_reg_7_ ( .D(n4111), .SI(n10923), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(n10922), .QN(n9821) );
  SDFFRXL fft_d2_q_reg_6_ ( .D(n4110), .SI(n10924), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(n10923), .QN(n9820) );
  SDFFRXL fft_d2_q_reg_5_ ( .D(n4109), .SI(n10925), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10924), .QN(n9819) );
  SDFFRXL fft_d2_q_reg_4_ ( .D(n4108), .SI(n10926), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10925), .QN(n9818) );
  SDFFRXL fft_d2_q_reg_3_ ( .D(n4107), .SI(n10927), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10926), .QN(n9817) );
  SDFFRXL fft_d2_q_reg_2_ ( .D(n4106), .SI(n10928), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(n10927), .QN(n9816) );
  SDFFRXL fft_d2_q_reg_1_ ( .D(n4105), .SI(n10929), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10928), .QN(n9815) );
  SDFFRXL fft_d2_q_reg_0_ ( .D(n4104), .SI(fft_d1[31]), .SE(test_se), .CK(clk), 
        .RN(n9016), .Q(n10929), .QN(n9814) );
  SDFFRXL fft_d12_q_reg_31_ ( .D(n4103), .SI(n10579), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10578), .QN(n9813) );
  SDFFRXL fft_d12_q_reg_30_ ( .D(n4102), .SI(n10580), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(n10579), .QN(n9812) );
  SDFFRXL fft_d12_q_reg_29_ ( .D(n4101), .SI(n10581), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(n10580), .QN(n9811) );
  SDFFRXL fft_d12_q_reg_28_ ( .D(n4100), .SI(n10582), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(n10581), .QN(n9810) );
  SDFFRXL fft_d12_q_reg_27_ ( .D(n4099), .SI(n10583), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(n10582), .QN(n9809) );
  SDFFRXL fft_d12_q_reg_26_ ( .D(n4098), .SI(n10584), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(n10583), .QN(n9808) );
  SDFFRXL fft_d12_q_reg_25_ ( .D(n4097), .SI(n10585), .SE(test_se), .CK(clk), 
        .RN(n8955), .Q(n10584), .QN(n9807) );
  SDFFRXL fft_d12_q_reg_24_ ( .D(n4096), .SI(n10586), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10585), .QN(n9806) );
  SDFFRXL fft_d12_q_reg_23_ ( .D(n4095), .SI(n10587), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10586), .QN(n9805) );
  SDFFRXL fft_d12_q_reg_22_ ( .D(n4094), .SI(n10588), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10587), .QN(n9804) );
  SDFFRXL fft_d12_q_reg_21_ ( .D(n4093), .SI(n10589), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10588), .QN(n9803) );
  SDFFRXL fft_d12_q_reg_20_ ( .D(n4092), .SI(n10590), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(n10589), .QN(n9802) );
  SDFFRXL fft_d12_q_reg_19_ ( .D(n4091), .SI(n10591), .SE(test_se), .CK(clk), 
        .RN(n9003), .Q(n10590), .QN(n9801) );
  SDFFRXL fft_d12_q_reg_18_ ( .D(n4090), .SI(n10592), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10591), .QN(n9800) );
  SDFFRXL fft_d12_q_reg_17_ ( .D(n4089), .SI(n10593), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10592), .QN(n9799) );
  SDFFRXL fft_d12_q_reg_16_ ( .D(n4088), .SI(n10594), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(n10593), .QN(n9798) );
  SDFFRXL fft_d12_q_reg_15_ ( .D(n4087), .SI(n10595), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10594), .QN(n9797) );
  SDFFRXL fft_d12_q_reg_14_ ( .D(n4086), .SI(n10596), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10595), .QN(n9796) );
  SDFFRXL fft_d12_q_reg_13_ ( .D(n4085), .SI(n10597), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10596), .QN(n9795) );
  SDFFRXL fft_d12_q_reg_12_ ( .D(n4084), .SI(n10598), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10597), .QN(n9794) );
  SDFFRXL fft_d12_q_reg_11_ ( .D(n4083), .SI(n10599), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10598), .QN(n9793) );
  SDFFRXL fft_d12_q_reg_10_ ( .D(n4082), .SI(n10600), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10599), .QN(n9792) );
  SDFFRXL fft_d12_q_reg_9_ ( .D(n4081), .SI(n10601), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10600), .QN(n9791) );
  SDFFRXL fft_d12_q_reg_8_ ( .D(n4080), .SI(n10602), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(n10601), .QN(n9790) );
  SDFFRXL fft_d12_q_reg_7_ ( .D(n4079), .SI(n10603), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(n10602), .QN(n9789) );
  SDFFRXL fft_d12_q_reg_6_ ( .D(n4078), .SI(n10604), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(n10603), .QN(n9788) );
  SDFFRXL fft_d12_q_reg_5_ ( .D(n4077), .SI(n10605), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10604), .QN(n9787) );
  SDFFRXL fft_d12_q_reg_4_ ( .D(n4076), .SI(n10606), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10605), .QN(n9786) );
  SDFFRXL fft_d12_q_reg_3_ ( .D(n4075), .SI(n10607), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10606), .QN(n9785) );
  SDFFRXL fft_d12_q_reg_2_ ( .D(n4074), .SI(n10608), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(n10607), .QN(n9784) );
  SDFFRXL fft_d12_q_reg_1_ ( .D(n4073), .SI(n10609), .SE(test_se), .CK(clk), 
        .RN(n9011), .Q(n10608), .QN(n9783) );
  SDFFRXL fft_d12_q_reg_0_ ( .D(n4072), .SI(fft_d11[31]), .SE(test_se), .CK(
        clk), .RN(n9016), .Q(n10609), .QN(n9782) );
  SDFFRXL fft_d4_q_reg_31_ ( .D(n4071), .SI(n10835), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10834), .QN(n9781) );
  SDFFRXL fft_d4_q_reg_30_ ( .D(n4070), .SI(n10836), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(n10835), .QN(n9780) );
  SDFFRXL fft_d4_q_reg_29_ ( .D(n4069), .SI(n10837), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(n10836), .QN(n9779) );
  SDFFRXL fft_d4_q_reg_28_ ( .D(n4068), .SI(n10838), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(n10837), .QN(n9778) );
  SDFFRXL fft_d4_q_reg_27_ ( .D(n4067), .SI(n10839), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(n10838), .QN(n9777) );
  SDFFRXL fft_d4_q_reg_26_ ( .D(n4066), .SI(n10840), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(n10839), .QN(n9776) );
  SDFFRXL fft_d4_q_reg_25_ ( .D(n4065), .SI(n10841), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(n10840), .QN(n9775) );
  SDFFRXL fft_d4_q_reg_24_ ( .D(n4064), .SI(n10842), .SE(test_se), .CK(clk), 
        .RN(n8950), .Q(n10841), .QN(n9774) );
  SDFFRXL fft_d4_q_reg_23_ ( .D(n4063), .SI(n10843), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10842), .QN(n9773) );
  SDFFRXL fft_d4_q_reg_22_ ( .D(n4062), .SI(n10844), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10843), .QN(n9772) );
  SDFFRXL fft_d4_q_reg_21_ ( .D(n4061), .SI(n10845), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10844), .QN(n9771) );
  SDFFRXL fft_d4_q_reg_20_ ( .D(n4060), .SI(n10846), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(n10845), .QN(n9770) );
  SDFFRXL fft_d4_q_reg_19_ ( .D(n4059), .SI(n10847), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(n10846), .QN(n9769) );
  SDFFRXL fft_d4_q_reg_18_ ( .D(n4058), .SI(n10848), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10847), .QN(n9768) );
  SDFFRXL fft_d4_q_reg_17_ ( .D(n4057), .SI(n10849), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10848), .QN(n9767) );
  SDFFRXL fft_d4_q_reg_16_ ( .D(n4056), .SI(n10850), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(n10849), .QN(n9766) );
  SDFFRXL fft_d4_q_reg_15_ ( .D(n4055), .SI(n10851), .SE(test_se), .CK(clk), 
        .RN(n8982), .Q(n10850), .QN(n9765) );
  SDFFRXL fft_d4_q_reg_14_ ( .D(n4054), .SI(n10852), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10851), .QN(n9764) );
  SDFFRXL fft_d4_q_reg_13_ ( .D(n4053), .SI(n10853), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10852), .QN(n9763) );
  SDFFRXL fft_d4_q_reg_12_ ( .D(n4052), .SI(n10854), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10853), .QN(n9762) );
  SDFFRXL fft_d4_q_reg_11_ ( .D(n4051), .SI(n10855), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10854), .QN(n9761) );
  SDFFRXL fft_d4_q_reg_10_ ( .D(n4050), .SI(n10856), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10855), .QN(n9760) );
  SDFFRXL fft_d4_q_reg_9_ ( .D(n4049), .SI(n10857), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10856), .QN(n9759) );
  SDFFRXL fft_d4_q_reg_8_ ( .D(n4048), .SI(n10858), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(n10857), .QN(n9758) );
  SDFFRXL fft_d4_q_reg_7_ ( .D(n4047), .SI(n10859), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(n10858), .QN(n9757) );
  SDFFRXL fft_d4_q_reg_6_ ( .D(n4046), .SI(n10860), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(n10859), .QN(n9756) );
  SDFFRXL fft_d4_q_reg_5_ ( .D(n4045), .SI(n10861), .SE(test_se), .CK(clk), 
        .RN(n8990), .Q(n10860), .QN(n9755) );
  SDFFRXL fft_d4_q_reg_4_ ( .D(n4044), .SI(n10862), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10861), .QN(n9754) );
  SDFFRXL fft_d4_q_reg_3_ ( .D(n4043), .SI(n10863), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10862), .QN(n9753) );
  SDFFRXL fft_d4_q_reg_2_ ( .D(n4042), .SI(n10864), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(n10863), .QN(n9752) );
  SDFFRXL fft_d4_q_reg_1_ ( .D(n4041), .SI(n10865), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(n10864), .QN(n9751) );
  SDFFRXL fft_d4_q_reg_0_ ( .D(n4040), .SI(fft_d3[31]), .SE(test_se), .CK(clk), 
        .RN(n9016), .Q(n10865), .QN(n9750) );
  SDFFRXL fft_d8_q_reg_31_ ( .D(n4039), .SI(n10707), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10706), .QN(n9749) );
  SDFFRXL fft_d8_q_reg_30_ ( .D(n4038), .SI(n10708), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(n10707), .QN(n9748) );
  SDFFRXL fft_d8_q_reg_29_ ( .D(n4037), .SI(n10709), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(n10708), .QN(n9747) );
  SDFFRXL fft_d8_q_reg_28_ ( .D(n4036), .SI(n10710), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(n10709), .QN(n9746) );
  SDFFRXL fft_d8_q_reg_27_ ( .D(n4035), .SI(n10711), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(n10710), .QN(n9745) );
  SDFFRXL fft_d8_q_reg_26_ ( .D(n4034), .SI(n10712), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(n10711), .QN(n9744) );
  SDFFRXL fft_d8_q_reg_25_ ( .D(n4033), .SI(n10713), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(n10712), .QN(n9743) );
  SDFFRXL fft_d8_q_reg_24_ ( .D(n4032), .SI(n10714), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(n10713), .QN(n9742) );
  SDFFRXL fft_d8_q_reg_23_ ( .D(n4031), .SI(n10715), .SE(test_se), .CK(clk), 
        .RN(n8945), .Q(n10714), .QN(n9741) );
  SDFFRXL fft_d8_q_reg_22_ ( .D(n4030), .SI(n10716), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10715), .QN(n9740) );
  SDFFRXL fft_d8_q_reg_21_ ( .D(n4029), .SI(n10717), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10716), .QN(n9739) );
  SDFFRXL fft_d8_q_reg_20_ ( .D(n4028), .SI(n10718), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(n10717), .QN(n9738) );
  SDFFRXL fft_d8_q_reg_19_ ( .D(n4027), .SI(n10719), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(n10718), .QN(n9737) );
  SDFFRXL fft_d8_q_reg_18_ ( .D(n4026), .SI(n10720), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10719), .QN(n9736) );
  SDFFRXL fft_d8_q_reg_17_ ( .D(n4025), .SI(n10721), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10720), .QN(n9735) );
  SDFFRXL fft_d8_q_reg_16_ ( .D(n4024), .SI(n10722), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(n10721), .QN(n9734) );
  SDFFRXL fft_d8_q_reg_15_ ( .D(n4023), .SI(n10723), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(n10722), .QN(n9733) );
  SDFFRXL fft_d8_q_reg_14_ ( .D(n4022), .SI(n10724), .SE(test_se), .CK(clk), 
        .RN(n8977), .Q(n10723), .QN(n9732) );
  SDFFRXL fft_d8_q_reg_13_ ( .D(n4021), .SI(n10725), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10724), .QN(n9731) );
  SDFFRXL fft_d8_q_reg_12_ ( .D(n4020), .SI(n10726), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10725), .QN(n9730) );
  SDFFRXL fft_d8_q_reg_11_ ( .D(n4019), .SI(n10727), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10726), .QN(n9729) );
  SDFFRXL fft_d8_q_reg_10_ ( .D(n4018), .SI(n10728), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10727), .QN(n9728) );
  SDFFRXL fft_d8_q_reg_9_ ( .D(n4017), .SI(n10729), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10728), .QN(n9727) );
  SDFFRXL fft_d8_q_reg_8_ ( .D(n4016), .SI(n10730), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(n10729), .QN(n9726) );
  SDFFRXL fft_d8_q_reg_7_ ( .D(n4015), .SI(n10731), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(n10730), .QN(n9725) );
  SDFFRXL fft_d8_q_reg_6_ ( .D(n4014), .SI(n10732), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(n10731), .QN(n9724) );
  SDFFRXL fft_d8_q_reg_5_ ( .D(n4013), .SI(n10733), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(n10732), .QN(n9723) );
  SDFFRXL fft_d8_q_reg_4_ ( .D(n4012), .SI(n10734), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10733), .QN(n9722) );
  SDFFRXL fft_d8_q_reg_3_ ( .D(n4011), .SI(n10735), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10734), .QN(n9721) );
  SDFFRXL fft_d8_q_reg_2_ ( .D(n40101), .SI(n10736), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(n10735), .QN(n9720) );
  SDFFRXL fft_d8_q_reg_1_ ( .D(n4009), .SI(n10737), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(n10736), .QN(n9719) );
  SDFFRXL fft_d8_q_reg_0_ ( .D(n4008), .SI(fft_d7[31]), .SE(test_se), .CK(clk), 
        .RN(n9016), .Q(n10737), .QN(n9718) );
  SDFFRXL fft_d0_q_reg_31_ ( .D(n4007), .SI(n10963), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(n10962), .QN(n9717) );
  SDFFRXL fft_d0_q_reg_30_ ( .D(n4006), .SI(n10964), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(n10963), .QN(n9716) );
  SDFFRXL fft_d0_q_reg_29_ ( .D(n4005), .SI(n10965), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(n10964), .QN(n9715) );
  SDFFRXL fft_d0_q_reg_28_ ( .D(n4004), .SI(n10966), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(n10965), .QN(n9714) );
  SDFFRXL fft_d0_q_reg_27_ ( .D(n4003), .SI(n10967), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(n10966), .QN(n9713) );
  SDFFRXL fft_d0_q_reg_26_ ( .D(n4002), .SI(n10968), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(n10967), .QN(n9712) );
  SDFFRXL fft_d0_q_reg_25_ ( .D(n4001), .SI(n10969), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(n10968), .QN(n9711) );
  SDFFRXL fft_d0_q_reg_24_ ( .D(n4000), .SI(n10970), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(n10969), .QN(n9710) );
  SDFFRXL fft_d0_q_reg_23_ ( .D(n3999), .SI(n10971), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(n10970), .QN(n9709) );
  SDFFRXL fft_d0_q_reg_22_ ( .D(n3998), .SI(n10972), .SE(test_se), .CK(clk), 
        .RN(n8940), .Q(n10971), .QN(n9708) );
  SDFFRXL fft_d0_q_reg_21_ ( .D(n3997), .SI(n10973), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(n10972), .QN(n9707) );
  SDFFRXL fft_d0_q_reg_20_ ( .D(n3996), .SI(n10974), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(n10973), .QN(n9706) );
  SDFFRXL fft_d0_q_reg_19_ ( .D(n3995), .SI(n10975), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(n10974), .QN(n9705) );
  SDFFRXL fft_d0_q_reg_18_ ( .D(n3994), .SI(n10976), .SE(test_se), .CK(clk), 
        .RN(n9008), .Q(n10975), .QN(n9704) );
  SDFFRXL fft_d0_q_reg_17_ ( .D(n3993), .SI(n10977), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(n10976), .QN(n9703) );
  SDFFRXL fft_d0_q_reg_16_ ( .D(n3992), .SI(n10978), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(n10977), .QN(n9702) );
  SDFFRXL fft_d0_q_reg_15_ ( .D(n3991), .SI(n10979), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(n10978), .QN(n9701) );
  SDFFRXL fft_d0_q_reg_14_ ( .D(n3990), .SI(n10980), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(n10979), .QN(n9700) );
  SDFFRXL fft_d0_q_reg_13_ ( .D(n3989), .SI(n10981), .SE(test_se), .CK(clk), 
        .RN(n8972), .Q(n10980), .QN(n9699) );
  SDFFRXL fft_d0_q_reg_12_ ( .D(n3988), .SI(n10982), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(n10981), .QN(n9698) );
  SDFFRXL fft_d0_q_reg_11_ ( .D(n3987), .SI(n10983), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(n10982), .QN(n9697) );
  SDFFRXL fft_d0_q_reg_10_ ( .D(n3986), .SI(n10984), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(n10983), .QN(n9696) );
  SDFFRXL fft_d0_q_reg_9_ ( .D(n3985), .SI(n10985), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(n10984), .QN(n9695) );
  SDFFRXL fft_d0_q_reg_8_ ( .D(n3984), .SI(n10986), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(n10985), .QN(n9694) );
  SDFFRXL fft_d0_q_reg_7_ ( .D(n3983), .SI(n10987), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(n10986), .QN(n9693) );
  SDFFRXL fft_d0_q_reg_6_ ( .D(n3982), .SI(n10988), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(n10987), .QN(n9692) );
  SDFFRXL fft_d0_q_reg_5_ ( .D(n3981), .SI(n10989), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(n10988), .QN(n9691) );
  SDFFRXL fft_d0_q_reg_4_ ( .D(n3980), .SI(n10990), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(n10989), .QN(n9690) );
  SDFFRXL fft_d0_q_reg_3_ ( .D(n3979), .SI(n10991), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(n10990), .QN(n9689) );
  SDFFRXL fft_d0_q_reg_2_ ( .D(n3978), .SI(n10992), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(n10991), .QN(n9688) );
  SDFFRXL fft_d0_q_reg_1_ ( .D(n3977), .SI(n10993), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(n10992), .QN(n9687) );
  SDFFRXL fft_d0_q_reg_0_ ( .D(n3976), .SI(done), .SE(test_se), .CK(clk), .RN(
        n9016), .Q(n10993), .QN(n9686) );
  SDFFRXL Analysis_STATE_reg ( .D(n3462), .SI(n11189), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(n6193), .QN(n10475) );
  SDFFRXL AnalysisOutput_STATE_reg ( .D(n3461), .SI(test_si), .SE(test_se), 
        .CK(clk), .RN(n9127), .Q(n11189), .QN(n9685) );
  SDFFRXL fft_dmax_reg_0_ ( .D(N1193), .SI(fft_d15[31]), .SE(test_se), .CK(clk), .RN(n8938), .Q(n10513), .QN(n2850) );
  SDFFRXL fft_dmax_reg_31_ ( .D(N1224), .SI(n10483), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10482), .QN(n2860) );
  SDFFRXL fft_dmax_reg_30_ ( .D(N1223), .SI(n10484), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10483), .QN(n2870) );
  SDFFRXL fft_dmax_reg_29_ ( .D(N1222), .SI(n10485), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10484), .QN(n2880) );
  SDFFRXL fft_dmax_reg_28_ ( .D(N1221), .SI(n10486), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10485), .QN(n2890) );
  SDFFRXL fft_dmax_reg_27_ ( .D(N1220), .SI(n10487), .SE(test_se), .CK(clk), 
        .RN(n8935), .Q(n10486), .QN(n290) );
  SDFFRXL fft_dmax_reg_26_ ( .D(N1219), .SI(n10488), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10487), .QN(n291) );
  SDFFRXL fft_dmax_reg_25_ ( .D(N1218), .SI(n10489), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10488), .QN(n292) );
  SDFFRXL fft_dmax_reg_24_ ( .D(N1217), .SI(n10490), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10489), .QN(n293) );
  SDFFRXL fft_dmax_reg_23_ ( .D(N1216), .SI(n10491), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10490), .QN(n294) );
  SDFFRXL fft_dmax_reg_22_ ( .D(N1215), .SI(n10492), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10491), .QN(n295) );
  SDFFRXL fft_dmax_reg_21_ ( .D(N1214), .SI(n10493), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10492), .QN(n296) );
  SDFFRXL fft_dmax_reg_20_ ( .D(N1213), .SI(n10494), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10493), .QN(n297) );
  SDFFRXL fft_dmax_reg_19_ ( .D(N1212), .SI(n10495), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10494), .QN(n298) );
  SDFFRXL fft_dmax_reg_18_ ( .D(N1211), .SI(n10496), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10495), .QN(n299) );
  SDFFRXL fft_dmax_reg_17_ ( .D(N1210), .SI(n10497), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10496), .QN(n3000) );
  SDFFRXL fft_dmax_reg_16_ ( .D(N1209), .SI(n10498), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10497), .QN(n3010) );
  SDFFRXL fft_dmax_reg_15_ ( .D(N1208), .SI(n10499), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10498), .QN(n3020) );
  SDFFRXL fft_dmax_reg_14_ ( .D(N1207), .SI(n10500), .SE(test_se), .CK(clk), 
        .RN(n8936), .Q(n10499), .QN(n3030) );
  SDFFRXL fft_dmax_reg_13_ ( .D(N1206), .SI(n10501), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10500), .QN(n3040) );
  SDFFRXL fft_dmax_reg_12_ ( .D(N1205), .SI(n10502), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10501), .QN(n3050) );
  SDFFRXL fft_dmax_reg_11_ ( .D(N1204), .SI(n10503), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10502), .QN(n3060) );
  SDFFRXL fft_dmax_reg_10_ ( .D(N1203), .SI(n10504), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10503), .QN(n30700) );
  SDFFRXL fft_dmax_reg_9_ ( .D(N1202), .SI(n10505), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10504), .QN(n3080) );
  SDFFRXL fft_dmax_reg_8_ ( .D(N1201), .SI(n10506), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10505), .QN(n3090) );
  SDFFRXL fft_dmax_reg_7_ ( .D(N1200), .SI(n10507), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10506), .QN(n3100) );
  SDFFRXL fft_dmax_reg_6_ ( .D(N1199), .SI(n10508), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10507), .QN(n3110) );
  SDFFRXL fft_dmax_reg_5_ ( .D(N1198), .SI(n10509), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10508), .QN(n3120) );
  SDFFRXL fft_dmax_reg_4_ ( .D(N1197), .SI(n10510), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10509), .QN(n3130) );
  SDFFRXL fft_dmax_reg_3_ ( .D(N1196), .SI(n10511), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10510), .QN(n3140) );
  SDFFRXL fft_dmax_reg_2_ ( .D(N1195), .SI(n10512), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10511), .QN(n3150) );
  SDFFRXL fft_dmax_reg_1_ ( .D(N1194), .SI(n10513), .SE(test_se), .CK(clk), 
        .RN(n8937), .Q(n10512), .QN(n3160) );
  SDFFRXL freq_max_reg_3_ ( .D(N1192), .SI(n11209), .SE(test_se), .CK(clk), 
        .RN(n8938), .Q(n11210), .QN(n6196) );
  SDFFRXL freq_max_reg_2_ ( .D(N1191), .SI(n11208), .SE(test_se), .CK(clk), 
        .RN(n8938), .Q(n11209), .QN(n6197) );
  SDFFRXL freq_max_reg_1_ ( .D(N1190), .SI(n11207), .SE(test_se), .CK(clk), 
        .RN(n8938), .Q(n11208), .QN(n6198) );
  SDFFRXL freq_max_reg_0_ ( .D(N1189), .SI(fir_valid), .SE(test_se), .CK(clk), 
        .RN(n8938), .Q(n11207), .QN(n6199) );
  SDFFRXL counter_reg_0_ ( .D(n6187), .SI(n10994), .SE(test_se), .CK(clk), 
        .RN(n9128), .Q(counter[0]), .QN(n6075) );
  SDFFRXL counter_reg_1_ ( .D(n6184), .SI(counter[0]), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(counter[1]), .QN(n6074) );
  SDFFRXL counter_reg_2_ ( .D(n6183), .SI(counter[1]), .SE(test_se), .CK(clk), 
        .RN(n9128), .Q(counter[2]), .QN(n6073) );
  SDFFRXL counter_reg_3_ ( .D(n6182), .SI(counter[2]), .SE(test_se), .CK(clk), 
        .RN(n9128), .Q(counter[3]), .QN(n6072) );
  SDFFRXL d32_reg_31_ ( .D(n4936), .SI(d32[30]), .SE(test_se), .CK(clk), .RN(
        n9049), .Q(d32[31]) );
  SDFFRXL d30_reg_32_ ( .D(n4987), .SI(d30[31]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d30[32]) );
  SDFFRXL d30_reg_33_ ( .D(n4986), .SI(d30[32]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d30[33]) );
  SDFFRXL d30_reg_34_ ( .D(n4985), .SI(d30[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d30[34]) );
  SDFFRXL d30_reg_35_ ( .D(n4984), .SI(d30[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d30[35]) );
  SDFFRXL d31_reg_0_ ( .D(n4983), .SI(d30[35]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d31[0]) );
  SDFFRXL d31_reg_2_ ( .D(n4981), .SI(d31[1]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d31[2]) );
  SDFFRXL d31_reg_3_ ( .D(n4980), .SI(d31[2]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d31[3]) );
  SDFFRXL d31_reg_4_ ( .D(n4979), .SI(d31[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d31[4]) );
  SDFFRXL d31_reg_5_ ( .D(n4978), .SI(d31[4]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d31[5]) );
  SDFFRXL d31_reg_6_ ( .D(n4977), .SI(d31[5]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d31[6]) );
  SDFFRXL d31_reg_7_ ( .D(n4976), .SI(d31[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d31[7]) );
  SDFFRXL d31_reg_8_ ( .D(n4975), .SI(d31[7]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d31[8]) );
  SDFFRXL d31_reg_9_ ( .D(n4974), .SI(d31[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d31[9]) );
  SDFFRXL d31_reg_10_ ( .D(n4973), .SI(d31[9]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d31[10]) );
  SDFFRXL d31_reg_11_ ( .D(n4972), .SI(d31[10]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d31[11]) );
  SDFFRXL d31_reg_12_ ( .D(n4971), .SI(d31[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d31[12]) );
  SDFFRXL d31_reg_13_ ( .D(n4970), .SI(d31[12]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d31[13]) );
  SDFFRXL d31_reg_14_ ( .D(n4969), .SI(d31[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d31[14]) );
  SDFFRXL d31_reg_15_ ( .D(n4968), .SI(d31[14]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d31[15]) );
  SDFFRXL d05_reg_0_ ( .D(n5884), .SI(d04[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d05[0]) );
  SDFFRXL d06_reg_0_ ( .D(n5848), .SI(d05[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d06[0]) );
  SDFFRXL d07_reg_1_ ( .D(n5813), .SI(d07[0]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d07[1]) );
  SDFFRXL d07_reg_0_ ( .D(n5812), .SI(d06[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d07[0]) );
  SDFFRXL d09_reg_0_ ( .D(n5740), .SI(d08[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d09[0]) );
  SDFFRXL d10_reg_0_ ( .D(n5704), .SI(d09[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d10[0]) );
  SDFFRXL d11_reg_1_ ( .D(n5669), .SI(d11[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d11[1]) );
  SDFFRXL d11_reg_0_ ( .D(n5668), .SI(d10[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d11[0]) );
  SDFFRXL d12_reg_0_ ( .D(n5632), .SI(d11[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d12[0]) );
  SDFFRXL d13_reg_1_ ( .D(n5597), .SI(d13[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d13[1]) );
  SDFFRXL d13_reg_0_ ( .D(n5596), .SI(d12[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d13[0]) );
  SDFFRXL d14_reg_0_ ( .D(n5560), .SI(d13[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d14[0]) );
  SDFFRXL d17_reg_0_ ( .D(n5452), .SI(d16[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d17[0]) );
  SDFFRXL d18_reg_1_ ( .D(n5417), .SI(d18[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d18[1]) );
  SDFFRXL d18_reg_0_ ( .D(n5416), .SI(d17[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d18[0]) );
  SDFFRXL d19_reg_0_ ( .D(n5380), .SI(d18[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d19[0]) );
  SDFFRXL d20_reg_1_ ( .D(n5345), .SI(d20[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d20[1]) );
  SDFFRXL d20_reg_0_ ( .D(n5344), .SI(d19[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d20[0]) );
  SDFFRXL d21_reg_0_ ( .D(n5308), .SI(d20[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d21[0]) );
  SDFFRXL d22_reg_0_ ( .D(n5272), .SI(d21[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d22[0]) );
  SDFFRXL d24_reg_1_ ( .D(n5201), .SI(d24[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d24[1]) );
  SDFFRXL d24_reg_0_ ( .D(n5200), .SI(d23[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d24[0]) );
  SDFFRXL d25_reg_0_ ( .D(n5164), .SI(d24[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d25[0]) );
  SDFFRXL d26_reg_0_ ( .D(n5128), .SI(d25[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d26[0]) );
  SDFFRXL d30_reg_0_ ( .D(n5019), .SI(d29[35]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d30[0]) );
  SDFFRXL FFT_STATE_reg_1_ ( .D(n6178), .SI(n10476), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(n10472), .QN(n6190) );
  SDFFRXL FFT_STATE_reg_0_ ( .D(n6179), .SI(BF2I_b_s), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(n10476), .QN(n6194) );
  SDFFRXL BF2II_a00_r_reg_1_ ( .D(n4796), .SI(N130), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(N131), .QN(n6109) );
  SDFFRXL BF2II_a00_i_reg_1_ ( .D(n4792), .SI(N113), .SE(test_se), .CK(clk), 
        .RN(n9046), .Q(N114), .QN(n6093) );
  SDFFRXL BF2II_a00_r_reg_2_ ( .D(n4788), .SI(N131), .SE(test_se), .CK(clk), 
        .RN(n9045), .Q(N132), .QN(n6108) );
  SDFFRXL BF2II_a00_i_reg_2_ ( .D(n4784), .SI(N114), .SE(test_se), .CK(clk), 
        .RN(n9044), .Q(N115), .QN(n6092) );
  SDFFRXL BF2II_a00_r_reg_3_ ( .D(n4780), .SI(N132), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(N133), .QN(n6107) );
  SDFFRXL BF2II_a00_i_reg_3_ ( .D(n4776), .SI(N115), .SE(test_se), .CK(clk), 
        .RN(n9043), .Q(N116), .QN(n6091) );
  SDFFRXL BF2II_a00_r_reg_4_ ( .D(n4772), .SI(N133), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(N134), .QN(n6106) );
  SDFFRXL BF2II_a00_i_reg_4_ ( .D(n4768), .SI(N116), .SE(test_se), .CK(clk), 
        .RN(n9041), .Q(N117), .QN(n6090) );
  SDFFRXL BF2II_a00_r_reg_5_ ( .D(n4764), .SI(N134), .SE(test_se), .CK(clk), 
        .RN(n9040), .Q(N135), .QN(n6105) );
  SDFFRXL BF2II_a00_i_reg_5_ ( .D(n4760), .SI(N117), .SE(test_se), .CK(clk), 
        .RN(n9039), .Q(N118), .QN(n6089) );
  SDFFRXL BF2II_a00_r_reg_6_ ( .D(n4756), .SI(N135), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(N136), .QN(n6104) );
  SDFFRXL BF2II_a00_i_reg_6_ ( .D(n4752), .SI(N118), .SE(test_se), .CK(clk), 
        .RN(n9038), .Q(N119), .QN(n6088) );
  SDFFRXL BF2II_a00_r_reg_7_ ( .D(n4748), .SI(N136), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(N137), .QN(n6103) );
  SDFFRXL BF2II_a00_i_reg_7_ ( .D(n4744), .SI(N119), .SE(test_se), .CK(clk), 
        .RN(n9036), .Q(N120), .QN(n6087) );
  SDFFRXL BF2II_a00_r_reg_8_ ( .D(n4740), .SI(N137), .SE(test_se), .CK(clk), 
        .RN(n9035), .Q(N138), .QN(n6102) );
  SDFFRXL BF2II_a00_i_reg_8_ ( .D(n4736), .SI(N120), .SE(test_se), .CK(clk), 
        .RN(n9034), .Q(N121), .QN(n6086) );
  SDFFRXL BF2II_a00_r_reg_9_ ( .D(n4732), .SI(N138), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(N139), .QN(n6101) );
  SDFFRXL BF2II_a00_i_reg_9_ ( .D(n4728), .SI(N121), .SE(test_se), .CK(clk), 
        .RN(n9033), .Q(N122), .QN(n6085) );
  SDFFRXL BF2II_a00_r_reg_10_ ( .D(n4724), .SI(N139), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(N140), .QN(n6100) );
  SDFFRXL BF2II_a00_i_reg_10_ ( .D(n4720), .SI(N122), .SE(test_se), .CK(clk), 
        .RN(n9031), .Q(N123), .QN(n6084) );
  SDFFRXL BF2II_a00_r_reg_11_ ( .D(n4716), .SI(N140), .SE(test_se), .CK(clk), 
        .RN(n9030), .Q(N141), .QN(n6099) );
  SDFFRXL BF2II_a00_i_reg_11_ ( .D(n4712), .SI(N123), .SE(test_se), .CK(clk), 
        .RN(n9029), .Q(N124), .QN(n6083) );
  SDFFRXL BF2II_a00_r_reg_12_ ( .D(n4708), .SI(N141), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(N142), .QN(n6098) );
  SDFFRXL BF2II_a00_i_reg_12_ ( .D(n4704), .SI(N124), .SE(test_se), .CK(clk), 
        .RN(n9028), .Q(N125), .QN(n6082) );
  SDFFRXL BF2II_a00_r_reg_13_ ( .D(n4700), .SI(N142), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(N143), .QN(n6097) );
  SDFFRXL BF2II_a00_i_reg_13_ ( .D(n4696), .SI(N125), .SE(test_se), .CK(clk), 
        .RN(n9026), .Q(N126), .QN(n6081) );
  SDFFRXL BF2II_a00_r_reg_14_ ( .D(n4692), .SI(N143), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(N144), .QN(n6096) );
  SDFFRXL BF2II_a00_i_reg_14_ ( .D(n4688), .SI(N126), .SE(test_se), .CK(clk), 
        .RN(n9024), .Q(N127), .QN(n6080) );
  SDFFRXL BF2II_a00_r_reg_15_ ( .D(n4684), .SI(N144), .SE(test_se), .CK(clk), 
        .RN(n9023), .Q(N145), .QN(n6095) );
  SDFFRXL BF2II_a00_i_reg_15_ ( .D(n4680), .SI(N127), .SE(test_se), .CK(clk), 
        .RN(n9022), .Q(N128), .QN(n6079) );
  SDFFRXL BF2II_b00_r_reg_1_ ( .D(n4550), .SI(BF2II_b_xr_n[0]), .SE(test_se), 
        .CK(clk), .RN(n9046), .Q(BF2II_b_xr_n[1]), .QN(n6174) );
  SDFFRXL BF2II_b00_r_reg_2_ ( .D(n4549), .SI(BF2II_b_xr_n[1]), .SE(test_se), 
        .CK(clk), .RN(n9044), .Q(BF2II_b_xr_n[2]), .QN(n6173) );
  SDFFRXL BF2II_b00_r_reg_3_ ( .D(n4548), .SI(BF2II_b_xr_n[2]), .SE(test_se), 
        .CK(clk), .RN(n9042), .Q(BF2II_b_xr_n[3]), .QN(n6172) );
  SDFFRXL BF2II_b00_r_reg_4_ ( .D(n4547), .SI(BF2II_b_xr_n[3]), .SE(test_se), 
        .CK(clk), .RN(n9041), .Q(BF2II_b_xr_n[4]), .QN(n6171) );
  SDFFRXL BF2II_b00_r_reg_5_ ( .D(n4546), .SI(BF2II_b_xr_n[4]), .SE(test_se), 
        .CK(clk), .RN(n9039), .Q(BF2II_b_xr_n[5]), .QN(n6170) );
  SDFFRXL BF2II_b00_r_reg_6_ ( .D(n4545), .SI(BF2II_b_xr_n[5]), .SE(test_se), 
        .CK(clk), .RN(n9037), .Q(BF2II_b_xr_n[6]), .QN(n6169) );
  SDFFRXL BF2II_b00_r_reg_7_ ( .D(n4544), .SI(BF2II_b_xr_n[6]), .SE(test_se), 
        .CK(clk), .RN(n9036), .Q(BF2II_b_xr_n[7]), .QN(n6168) );
  SDFFRXL BF2II_b00_r_reg_8_ ( .D(n4543), .SI(BF2II_b_xr_n[7]), .SE(test_se), 
        .CK(clk), .RN(n9034), .Q(BF2II_b_xr_n[8]), .QN(n6167) );
  SDFFRXL BF2II_b00_r_reg_9_ ( .D(n4542), .SI(BF2II_b_xr_n[8]), .SE(test_se), 
        .CK(clk), .RN(n9032), .Q(BF2II_b_xr_n[9]), .QN(n6166) );
  SDFFRXL BF2II_b00_r_reg_10_ ( .D(n4541), .SI(BF2II_b_xr_n[9]), .SE(test_se), 
        .CK(clk), .RN(n9031), .Q(BF2II_b_xr_n[10]), .QN(n6165) );
  SDFFRXL BF2II_b00_r_reg_11_ ( .D(n4540), .SI(BF2II_b_xr_n[10]), .SE(test_se), 
        .CK(clk), .RN(n9029), .Q(BF2II_b_xr_n[11]), .QN(n6164) );
  SDFFRXL BF2II_b00_r_reg_12_ ( .D(n4539), .SI(BF2II_b_xr_n[11]), .SE(test_se), 
        .CK(clk), .RN(n9027), .Q(BF2II_b_xr_n[12]), .QN(n6163) );
  SDFFRXL BF2II_b00_r_reg_13_ ( .D(n4538), .SI(BF2II_b_xr_n[12]), .SE(test_se), 
        .CK(clk), .RN(n9025), .Q(BF2II_b_xr_n[13]), .QN(n6162) );
  SDFFRXL BF2II_b00_r_reg_14_ ( .D(n4537), .SI(BF2II_b_xr_n[13]), .SE(test_se), 
        .CK(clk), .RN(n9024), .Q(BF2II_b_xr_n[14]), .QN(n6161) );
  SDFFRXL BF2II_b00_r_reg_15_ ( .D(n4536), .SI(BF2II_b_xr_n[14]), .SE(test_se), 
        .CK(clk), .RN(n9020), .Q(BF2II_b_xr_n[15]), .QN(n6160) );
  SDFFRXL BF2II_b00_r_reg_16_ ( .D(n4535), .SI(BF2II_b_xr_n[15]), .SE(test_se), 
        .CK(clk), .RN(n9019), .Q(BF2II_b_xr_n[16]), .QN(n6159) );
  SDFFRXL BF2II_b00_r_reg_17_ ( .D(n4534), .SI(BF2II_b_xr_n[16]), .SE(test_se), 
        .CK(clk), .RN(n9014), .Q(BF2II_b_xr_n[17]), .QN(n6158) );
  SDFFRXL BF2II_b00_r_reg_18_ ( .D(n4533), .SI(BF2II_b_xr_n[17]), .SE(test_se), 
        .CK(clk), .RN(n9009), .Q(BF2II_b_xr_n[18]), .QN(n6157) );
  SDFFRXL BF2II_b00_r_reg_19_ ( .D(n4532), .SI(BF2II_b_xr_n[18]), .SE(test_se), 
        .CK(clk), .RN(n9004), .Q(BF2II_b_xr_n[19]), .QN(n6156) );
  SDFFRXL BF2II_b00_r_reg_20_ ( .D(n4531), .SI(BF2II_b_xr_n[19]), .SE(test_se), 
        .CK(clk), .RN(n8998), .Q(BF2II_b_xr_n[20]), .QN(n6155) );
  SDFFRXL BF2II_b00_r_reg_21_ ( .D(n4530), .SI(BF2II_b_xr_n[20]), .SE(test_se), 
        .CK(clk), .RN(n8993), .Q(BF2II_b_xr_n[21]), .QN(n6154) );
  SDFFRXL BF2II_b00_r_reg_22_ ( .D(n4529), .SI(BF2II_b_xr_n[21]), .SE(test_se), 
        .CK(clk), .RN(n8987), .Q(BF2II_b_xr_n[22]), .QN(n6153) );
  SDFFRXL BF2II_b00_r_reg_23_ ( .D(n4528), .SI(BF2II_b_xr_n[22]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[23]), .QN(n6152) );
  SDFFRXL BF2II_b00_r_reg_24_ ( .D(n4527), .SI(BF2II_b_xr_n[23]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[24]), .QN(n6151) );
  SDFFRXL BF2II_b00_r_reg_25_ ( .D(n4526), .SI(BF2II_b_xr_n[24]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[25]), .QN(n6150) );
  SDFFRXL BF2II_b00_r_reg_26_ ( .D(n4525), .SI(BF2II_b_xr_n[25]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[26]), .QN(n6149) );
  SDFFRXL BF2II_b00_r_reg_27_ ( .D(n4524), .SI(BF2II_b_xr_n[26]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[27]), .QN(n6148) );
  SDFFRXL BF2II_b00_r_reg_28_ ( .D(n4523), .SI(BF2II_b_xr_n[27]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[28]), .QN(n6147) );
  SDFFRXL BF2II_b00_r_reg_29_ ( .D(n4522), .SI(BF2II_b_xr_n[28]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[29]), .QN(n6146) );
  SDFFRXL BF2II_b00_r_reg_30_ ( .D(n4521), .SI(BF2II_b_xr_n[29]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[30]), .QN(n6145) );
  SDFFRXL BF2II_b00_r_reg_31_ ( .D(n4520), .SI(BF2II_b_xr_n[30]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xr_n[31]), .QN(n6144) );
  SDFFRXL BF2II_b00_i_reg_16_ ( .D(n4519), .SI(BF2II_b_xi_n[15]), .SE(test_se), 
        .CK(clk), .RN(n9019), .Q(BF2II_b_xi_n[16]), .QN(n6127) );
  SDFFRXL BF2II_b00_i_reg_31_ ( .D(n4518), .SI(BF2II_b_xi_n[30]), .SE(test_se), 
        .CK(clk), .RN(n8985), .Q(BF2II_b_xi_n[31]), .QN(n6112) );
  SDFFRXL BF2II_b00_i_reg_1_ ( .D(n4516), .SI(BF2II_b_xi_n[0]), .SE(test_se), 
        .CK(clk), .RN(n9046), .Q(BF2II_b_xi_n[1]), .QN(n6142) );
  SDFFRXL BF2II_b00_i_reg_2_ ( .D(n4515), .SI(BF2II_b_xi_n[1]), .SE(test_se), 
        .CK(clk), .RN(n9044), .Q(BF2II_b_xi_n[2]), .QN(n6141) );
  SDFFRXL BF2II_b00_i_reg_3_ ( .D(n4514), .SI(BF2II_b_xi_n[2]), .SE(test_se), 
        .CK(clk), .RN(n9042), .Q(BF2II_b_xi_n[3]), .QN(n6140) );
  SDFFRXL BF2II_b00_i_reg_4_ ( .D(n4513), .SI(BF2II_b_xi_n[3]), .SE(test_se), 
        .CK(clk), .RN(n9041), .Q(BF2II_b_xi_n[4]), .QN(n6139) );
  SDFFRXL BF2II_b00_i_reg_5_ ( .D(n4512), .SI(BF2II_b_xi_n[4]), .SE(test_se), 
        .CK(clk), .RN(n9039), .Q(BF2II_b_xi_n[5]), .QN(n6138) );
  SDFFRXL BF2II_b00_i_reg_6_ ( .D(n4511), .SI(BF2II_b_xi_n[5]), .SE(test_se), 
        .CK(clk), .RN(n9037), .Q(BF2II_b_xi_n[6]), .QN(n6137) );
  SDFFRXL BF2II_b00_i_reg_7_ ( .D(n4510), .SI(BF2II_b_xi_n[6]), .SE(test_se), 
        .CK(clk), .RN(n9036), .Q(BF2II_b_xi_n[7]), .QN(n6136) );
  SDFFRXL BF2II_b00_i_reg_8_ ( .D(n4509), .SI(BF2II_b_xi_n[7]), .SE(test_se), 
        .CK(clk), .RN(n9034), .Q(BF2II_b_xi_n[8]), .QN(n6135) );
  SDFFRXL BF2II_b00_i_reg_9_ ( .D(n4508), .SI(BF2II_b_xi_n[8]), .SE(test_se), 
        .CK(clk), .RN(n9032), .Q(BF2II_b_xi_n[9]), .QN(n6134) );
  SDFFRXL BF2II_b00_i_reg_10_ ( .D(n4507), .SI(BF2II_b_xi_n[9]), .SE(test_se), 
        .CK(clk), .RN(n9030), .Q(BF2II_b_xi_n[10]), .QN(n6133) );
  SDFFRXL BF2II_b00_i_reg_11_ ( .D(n4506), .SI(BF2II_b_xi_n[10]), .SE(test_se), 
        .CK(clk), .RN(n9029), .Q(BF2II_b_xi_n[11]), .QN(n6132) );
  SDFFRXL BF2II_b00_i_reg_12_ ( .D(n4505), .SI(BF2II_b_xi_n[11]), .SE(test_se), 
        .CK(clk), .RN(n9027), .Q(BF2II_b_xi_n[12]), .QN(n6131) );
  SDFFRXL BF2II_b00_i_reg_13_ ( .D(n4504), .SI(BF2II_b_xi_n[12]), .SE(test_se), 
        .CK(clk), .RN(n9025), .Q(BF2II_b_xi_n[13]), .QN(n6130) );
  SDFFRXL BF2II_b00_i_reg_14_ ( .D(n4503), .SI(BF2II_b_xi_n[13]), .SE(test_se), 
        .CK(clk), .RN(n9024), .Q(BF2II_b_xi_n[14]), .QN(n6129) );
  SDFFRXL BF2II_b00_i_reg_15_ ( .D(n4502), .SI(BF2II_b_xi_n[14]), .SE(test_se), 
        .CK(clk), .RN(n9020), .Q(BF2II_b_xi_n[15]), .QN(n6128) );
  SDFFRXL BF2II_b00_i_reg_17_ ( .D(n4501), .SI(BF2II_b_xi_n[16]), .SE(test_se), 
        .CK(clk), .RN(n9014), .Q(BF2II_b_xi_n[17]), .QN(n6126) );
  SDFFRXL BF2II_b00_i_reg_18_ ( .D(n4500), .SI(BF2II_b_xi_n[17]), .SE(test_se), 
        .CK(clk), .RN(n9009), .Q(BF2II_b_xi_n[18]), .QN(n6125) );
  SDFFRXL BF2II_b00_i_reg_19_ ( .D(n4499), .SI(BF2II_b_xi_n[18]), .SE(test_se), 
        .CK(clk), .RN(n9004), .Q(BF2II_b_xi_n[19]), .QN(n6124) );
  SDFFRXL BF2II_b00_i_reg_20_ ( .D(n4498), .SI(BF2II_b_xi_n[19]), .SE(test_se), 
        .CK(clk), .RN(n8998), .Q(BF2II_b_xi_n[20]), .QN(n6123) );
  SDFFRXL BF2II_b00_i_reg_21_ ( .D(n4497), .SI(BF2II_b_xi_n[20]), .SE(test_se), 
        .CK(clk), .RN(n8993), .Q(BF2II_b_xi_n[21]), .QN(n6122) );
  SDFFRXL BF2II_b00_i_reg_22_ ( .D(n4496), .SI(BF2II_b_xi_n[21]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xi_n[22]), .QN(n6121) );
  SDFFRXL BF2II_b00_i_reg_23_ ( .D(n4495), .SI(BF2II_b_xi_n[22]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xi_n[23]), .QN(n6120) );
  SDFFRXL BF2II_b00_i_reg_24_ ( .D(n4494), .SI(BF2II_b_xi_n[23]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xi_n[24]), .QN(n6119) );
  SDFFRXL BF2II_b00_i_reg_25_ ( .D(n4493), .SI(BF2II_b_xi_n[24]), .SE(test_se), 
        .CK(clk), .RN(n8986), .Q(BF2II_b_xi_n[25]), .QN(n6118) );
  SDFFRXL BF2II_b00_i_reg_26_ ( .D(n4492), .SI(BF2II_b_xi_n[25]), .SE(test_se), 
        .CK(clk), .RN(n8985), .Q(BF2II_b_xi_n[26]), .QN(n6117) );
  SDFFRXL BF2II_b00_i_reg_27_ ( .D(n4491), .SI(BF2II_b_xi_n[26]), .SE(test_se), 
        .CK(clk), .RN(n8985), .Q(BF2II_b_xi_n[27]), .QN(n6116) );
  SDFFRXL BF2II_b00_i_reg_28_ ( .D(n4490), .SI(BF2II_b_xi_n[27]), .SE(test_se), 
        .CK(clk), .RN(n8985), .Q(BF2II_b_xi_n[28]), .QN(n6115) );
  SDFFRXL BF2II_b00_i_reg_29_ ( .D(n4489), .SI(BF2II_b_xi_n[28]), .SE(test_se), 
        .CK(clk), .RN(n8985), .Q(BF2II_b_xi_n[29]), .QN(n6114) );
  SDFFRXL BF2II_b00_i_reg_30_ ( .D(n4488), .SI(BF2II_b_xi_n[29]), .SE(test_se), 
        .CK(clk), .RN(n8985), .Q(BF2II_b_xi_n[30]), .QN(n6113) );
  SDFFRXL d32_reg_16_ ( .D(n4951), .SI(d31[31]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d32[16]) );
  SDFFRXL fft_d15_q_reg_31_ ( .D(n4487), .SI(fft_d15_q[30]), .SE(test_se), 
        .CK(clk), .RN(n8985), .Q(fft_d15_q[31]), .QN(n10197) );
  SDFFRXL fft_d15_q_reg_30_ ( .D(n4486), .SI(fft_d15_q[29]), .SE(test_se), 
        .CK(clk), .RN(n8980), .Q(fft_d15_q[30]), .QN(n10196) );
  SDFFRXL fft_d15_q_reg_28_ ( .D(n4484), .SI(fft_d15_q[27]), .SE(test_se), 
        .CK(clk), .RN(n8970), .Q(fft_d15_q[28]), .QN(n10194) );
  SDFFRXL fft_d15_q_reg_26_ ( .D(n4482), .SI(fft_d15_q[25]), .SE(test_se), 
        .CK(clk), .RN(n8960), .Q(fft_d15_q[26]), .QN(n10192) );
  SDFFRXL fft_d15_q_reg_15_ ( .D(n4471), .SI(fft_d15_q[14]), .SE(test_se), 
        .CK(clk), .RN(n8983), .Q(fft_d15_q[15]), .QN(n10181) );
  SDFFRXL fft_d15_q_reg_14_ ( .D(n4470), .SI(fft_d15_q[13]), .SE(test_se), 
        .CK(clk), .RN(n8978), .Q(fft_d15_q[14]), .QN(n10180) );
  SDFFRXL fft_d15_q_reg_12_ ( .D(n4468), .SI(fft_d15_q[11]), .SE(test_se), 
        .CK(clk), .RN(n8968), .Q(fft_d15_q[12]), .QN(n10178) );
  SDFFRXL fft_d15_q_reg_10_ ( .D(n4466), .SI(fft_d15_q[9]), .SE(test_se), .CK(
        clk), .RN(n8958), .Q(fft_d15_q[10]), .QN(n10176) );
  SDFFRXL fft_d15_q_reg_23_ ( .D(n4479), .SI(fft_d15_q[22]), .SE(test_se), 
        .CK(clk), .RN(n8946), .Q(fft_d15_q[23]), .QN(n10189) );
  SDFFRXL fft_d15_q_reg_22_ ( .D(n4478), .SI(fft_d15_q[21]), .SE(test_se), 
        .CK(clk), .RN(n8941), .Q(fft_d15_q[22]), .QN(n10188) );
  SDFFRXL fft_d15_q_reg_21_ ( .D(n4477), .SI(fft_d15_q[20]), .SE(test_se), 
        .CK(clk), .RN(n8993), .Q(fft_d15_q[21]), .QN(n10187) );
  SDFFRXL fft_d15_q_reg_20_ ( .D(n4476), .SI(fft_d15_q[19]), .SE(test_se), 
        .CK(clk), .RN(n8998), .Q(fft_d15_q[20]), .QN(n10186) );
  SDFFRXL fft_d15_q_reg_19_ ( .D(n4475), .SI(fft_d15_q[18]), .SE(test_se), 
        .CK(clk), .RN(n9003), .Q(fft_d15_q[19]), .QN(n10185) );
  SDFFRXL fft_d15_q_reg_18_ ( .D(n4474), .SI(fft_d15_q[17]), .SE(test_se), 
        .CK(clk), .RN(n9009), .Q(fft_d15_q[18]), .QN(n10184) );
  SDFFRXL fft_d15_q_reg_17_ ( .D(n4473), .SI(fft_d15_q[16]), .SE(test_se), 
        .CK(clk), .RN(n9014), .Q(fft_d15_q[17]), .QN(n10183) );
  SDFFRXL fft_d15_q_reg_7_ ( .D(n4463), .SI(fft_d15_q[6]), .SE(test_se), .CK(
        clk), .RN(n8943), .Q(fft_d15_q[7]), .QN(n10173) );
  SDFFRXL fft_d15_q_reg_6_ ( .D(n4462), .SI(fft_d15_q[5]), .SE(test_se), .CK(
        clk), .RN(n8938), .Q(fft_d15_q[6]), .QN(n10172) );
  SDFFRXL fft_d15_q_reg_5_ ( .D(n4461), .SI(fft_d15_q[4]), .SE(test_se), .CK(
        clk), .RN(n8991), .Q(fft_d15_q[5]), .QN(n10171) );
  SDFFRXL fft_d15_q_reg_4_ ( .D(n4460), .SI(fft_d15_q[3]), .SE(test_se), .CK(
        clk), .RN(n8996), .Q(fft_d15_q[4]), .QN(n10170) );
  SDFFRXL fft_d15_q_reg_3_ ( .D(n4459), .SI(fft_d15_q[2]), .SE(test_se), .CK(
        clk), .RN(n9001), .Q(fft_d15_q[3]), .QN(n10169) );
  SDFFRXL fft_d15_q_reg_2_ ( .D(n4458), .SI(fft_d15_q[1]), .SE(test_se), .CK(
        clk), .RN(n9006), .Q(fft_d15_q[2]), .QN(n10168) );
  SDFFRXL fft_d15_q_reg_1_ ( .D(n4457), .SI(fft_d15_q[0]), .SE(test_se), .CK(
        clk), .RN(n9011), .Q(fft_d15_q[1]), .QN(n10167) );
  SDFFRXL fft_d15_q_reg_24_ ( .D(n4480), .SI(fft_d15_q[23]), .SE(test_se), 
        .CK(clk), .RN(n8951), .Q(fft_d15_q[24]), .QN(n10190) );
  SDFFRXL fft_d15_q_reg_8_ ( .D(n4464), .SI(fft_d15_q[7]), .SE(test_se), .CK(
        clk), .RN(n8948), .Q(fft_d15_q[8]), .QN(n10174) );
  SDFFRXL d31_reg_1_ ( .D(n4982), .SI(d31[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d31[1]) );
  SDFFRXL fft_d15_q_reg_29_ ( .D(n4485), .SI(fft_d15_q[28]), .SE(test_se), 
        .CK(clk), .RN(n8975), .Q(fft_d15_q[29]), .QN(n10195) );
  SDFFRXL fft_d15_q_reg_27_ ( .D(n4483), .SI(fft_d15_q[26]), .SE(test_se), 
        .CK(clk), .RN(n8965), .Q(fft_d15_q[27]), .QN(n10193) );
  SDFFRXL fft_d15_q_reg_25_ ( .D(n4481), .SI(fft_d15_q[24]), .SE(test_se), 
        .CK(clk), .RN(n8955), .Q(fft_d15_q[25]), .QN(n10191) );
  SDFFRXL fft_d15_q_reg_13_ ( .D(n4469), .SI(fft_d15_q[12]), .SE(test_se), 
        .CK(clk), .RN(n8973), .Q(fft_d15_q[13]), .QN(n10179) );
  SDFFRXL fft_d15_q_reg_11_ ( .D(n4467), .SI(fft_d15_q[10]), .SE(test_se), 
        .CK(clk), .RN(n8963), .Q(fft_d15_q[11]), .QN(n10177) );
  SDFFRXL fft_d15_q_reg_9_ ( .D(n4465), .SI(fft_d15_q[8]), .SE(test_se), .CK(
        clk), .RN(n8953), .Q(fft_d15_q[9]), .QN(n10175) );
  SDFFRXL fft_d15_q_reg_16_ ( .D(n4472), .SI(fft_d15_q[15]), .SE(test_se), 
        .CK(clk), .RN(n9019), .Q(fft_d15_q[16]), .QN(n10182) );
  SDFFRXL fft_d15_q_reg_0_ ( .D(n4456), .SI(fft_d14[31]), .SE(test_se), .CK(
        clk), .RN(n9017), .Q(fft_d15_q[0]), .QN(n10166) );
  SDFFRXL BF2II_a00_i_reg_0_ ( .D(n4804), .SI(n6193), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(N113), .QN(n6094) );
  SDFFRXL BF2II_b00_r_reg_0_ ( .D(n4551), .SI(BF2II_b_xi_n[31]), .SE(test_se), 
        .CK(clk), .RN(n9047), .Q(BF2II_b_xr_n[0]), .QN(n6175) );
  SDFFRXL BF2II_b00_i_reg_0_ ( .D(n4517), .SI(n11092), .SE(test_se), .CK(clk), 
        .RN(n9047), .Q(BF2II_b_xi_n[0]), .QN(n6143) );
  SDFFRXL BF2I_a00_r_reg_1_ ( .D(n4920), .SI(BF2I_a_xr_n[0]), .SE(test_se), 
        .CK(clk), .RN(n9047), .Q(BF2I_a_xr_n[1]), .QN(n1936) );
  SDFFRXL BF2I_a00_r_reg_2_ ( .D(n4912), .SI(BF2I_a_xr_n[1]), .SE(test_se), 
        .CK(clk), .RN(n9045), .Q(BF2I_a_xr_n[2]), .QN(n1928) );
  SDFFRXL BF2I_a00_r_reg_3_ ( .D(n4904), .SI(BF2I_a_xr_n[2]), .SE(test_se), 
        .CK(clk), .RN(n9043), .Q(BF2I_a_xr_n[3]), .QN(n1920) );
  SDFFRXL BF2I_a00_r_reg_4_ ( .D(n4896), .SI(BF2I_a_xr_n[3]), .SE(test_se), 
        .CK(clk), .RN(n9042), .Q(BF2I_a_xr_n[4]), .QN(n1912) );
  SDFFRXL BF2I_a00_r_reg_5_ ( .D(n4888), .SI(BF2I_a_xr_n[4]), .SE(test_se), 
        .CK(clk), .RN(n9040), .Q(BF2I_a_xr_n[5]), .QN(n1904) );
  SDFFRXL BF2I_a00_r_reg_6_ ( .D(n4880), .SI(BF2I_a_xr_n[5]), .SE(test_se), 
        .CK(clk), .RN(n9038), .Q(BF2I_a_xr_n[6]), .QN(n1896) );
  SDFFRXL BF2I_a00_r_reg_7_ ( .D(n4872), .SI(BF2I_a_xr_n[6]), .SE(test_se), 
        .CK(clk), .RN(n9037), .Q(BF2I_a_xr_n[7]), .QN(n1888) );
  SDFFRXL BF2I_a00_r_reg_8_ ( .D(n4864), .SI(BF2I_a_xr_n[7]), .SE(test_se), 
        .CK(clk), .RN(n9035), .Q(BF2I_a_xr_n[8]), .QN(n1880) );
  SDFFRXL BF2I_a00_r_reg_9_ ( .D(n4856), .SI(BF2I_a_xr_n[8]), .SE(test_se), 
        .CK(clk), .RN(n9033), .Q(BF2I_a_xr_n[9]), .QN(n1872) );
  SDFFRXL BF2I_a00_r_reg_10_ ( .D(n4848), .SI(BF2I_a_xr_n[9]), .SE(test_se), 
        .CK(clk), .RN(n9032), .Q(BF2I_a_xr_n[10]), .QN(n1864) );
  SDFFRXL BF2I_a00_r_reg_11_ ( .D(n4840), .SI(BF2I_a_xr_n[10]), .SE(test_se), 
        .CK(clk), .RN(n9030), .Q(BF2I_a_xr_n[11]), .QN(n1856) );
  SDFFRXL BF2I_a00_r_reg_12_ ( .D(n4832), .SI(BF2I_a_xr_n[11]), .SE(test_se), 
        .CK(clk), .RN(n9028), .Q(BF2I_a_xr_n[12]), .QN(n1848) );
  SDFFRXL BF2I_a00_r_reg_13_ ( .D(n4824), .SI(BF2I_a_xr_n[12]), .SE(test_se), 
        .CK(clk), .RN(n9026), .Q(BF2I_a_xr_n[13]), .QN(n1840) );
  SDFFRXL BF2I_a00_r_reg_14_ ( .D(n4816), .SI(BF2I_a_xr_n[13]), .SE(test_se), 
        .CK(clk), .RN(n9025), .Q(BF2I_a_xr_n[14]), .QN(n1832) );
  SDFFRXL BF2I_a00_r_reg_15_ ( .D(n4808), .SI(BF2I_a_xr_n[14]), .SE(test_se), 
        .CK(clk), .RN(n9023), .Q(BF2I_a_xr_n[15]), .QN(n1824) );
  SDFFRXL BF2I_b00_r_reg_1_ ( .D(n4676), .SI(BF2I_b_xr_n[0]), .SE(test_se), 
        .CK(clk), .RN(n9046), .Q(BF2I_b_xr_n[1]), .QN(n1723) );
  SDFFRXL BF2I_b00_r_reg_2_ ( .D(n4674), .SI(BF2I_b_xr_n[1]), .SE(test_se), 
        .CK(clk), .RN(n9044), .Q(BF2I_b_xr_n[2]), .QN(n1721) );
  SDFFRXL BF2I_b00_r_reg_3_ ( .D(n4672), .SI(BF2I_b_xr_n[2]), .SE(test_se), 
        .CK(clk), .RN(n9042), .Q(BF2I_b_xr_n[3]), .QN(n1719) );
  SDFFRXL BF2I_b00_r_reg_4_ ( .D(n4670), .SI(BF2I_b_xr_n[3]), .SE(test_se), 
        .CK(clk), .RN(n9041), .Q(BF2I_b_xr_n[4]), .QN(n1717) );
  SDFFRXL BF2I_b00_r_reg_5_ ( .D(n4668), .SI(BF2I_b_xr_n[4]), .SE(test_se), 
        .CK(clk), .RN(n9039), .Q(BF2I_b_xr_n[5]), .QN(n1715) );
  SDFFRXL BF2I_b00_r_reg_6_ ( .D(n4666), .SI(BF2I_b_xr_n[5]), .SE(test_se), 
        .CK(clk), .RN(n9037), .Q(BF2I_b_xr_n[6]), .QN(n1713) );
  SDFFRXL BF2I_b00_r_reg_7_ ( .D(n4664), .SI(BF2I_b_xr_n[6]), .SE(test_se), 
        .CK(clk), .RN(n9036), .Q(BF2I_b_xr_n[7]), .QN(n1711) );
  SDFFRXL BF2I_b00_r_reg_8_ ( .D(n4662), .SI(BF2I_b_xr_n[7]), .SE(test_se), 
        .CK(clk), .RN(n9034), .Q(BF2I_b_xr_n[8]), .QN(n1709) );
  SDFFRXL BF2I_b00_r_reg_9_ ( .D(n4660), .SI(BF2I_b_xr_n[8]), .SE(test_se), 
        .CK(clk), .RN(n9032), .Q(BF2I_b_xr_n[9]), .QN(n1707) );
  SDFFRXL BF2I_b00_r_reg_10_ ( .D(n4658), .SI(BF2I_b_xr_n[9]), .SE(test_se), 
        .CK(clk), .RN(n9031), .Q(BF2I_b_xr_n[10]), .QN(n1705) );
  SDFFRXL BF2I_b00_r_reg_11_ ( .D(n4656), .SI(BF2I_b_xr_n[10]), .SE(test_se), 
        .CK(clk), .RN(n9029), .Q(BF2I_b_xr_n[11]), .QN(n1703) );
  SDFFRXL BF2I_b00_r_reg_12_ ( .D(n4654), .SI(BF2I_b_xr_n[11]), .SE(test_se), 
        .CK(clk), .RN(n9027), .Q(BF2I_b_xr_n[12]), .QN(n1701) );
  SDFFRXL BF2I_b00_r_reg_13_ ( .D(n4652), .SI(BF2I_b_xr_n[12]), .SE(test_se), 
        .CK(clk), .RN(n9026), .Q(BF2I_b_xr_n[13]), .QN(n1699) );
  SDFFRXL BF2I_b00_r_reg_14_ ( .D(n4650), .SI(BF2I_b_xr_n[13]), .SE(test_se), 
        .CK(clk), .RN(n9024), .Q(BF2I_b_xr_n[14]), .QN(n1697) );
  SDFFRXL BF2I_b00_r_reg_15_ ( .D(n4648), .SI(BF2I_b_xr_n[14]), .SE(test_se), 
        .CK(clk), .RN(n9020), .Q(BF2I_b_xr_n[15]), .QN(n1695) );
  SDFFRXL BF2I_b00_r_reg_16_ ( .D(n4646), .SI(BF2I_b_xr_n[15]), .SE(test_se), 
        .CK(clk), .RN(n9019), .Q(BF2I_b_xr_n[16]), .QN(n1693) );
  SDFFRXL BF2I_b00_r_reg_17_ ( .D(n4644), .SI(BF2I_b_xr_n[16]), .SE(test_se), 
        .CK(clk), .RN(n9014), .Q(BF2I_b_xr_n[17]), .QN(n1691) );
  SDFFRXL BF2I_b00_r_reg_18_ ( .D(n4642), .SI(BF2I_b_xr_n[17]), .SE(test_se), 
        .CK(clk), .RN(n9009), .Q(BF2I_b_xr_n[18]), .QN(n1689) );
  SDFFRXL BF2I_b00_r_reg_19_ ( .D(n4640), .SI(BF2I_b_xr_n[18]), .SE(test_se), 
        .CK(clk), .RN(n9004), .Q(BF2I_b_xr_n[19]), .QN(n1687) );
  SDFFRXL BF2I_b00_r_reg_20_ ( .D(n4638), .SI(BF2I_b_xr_n[19]), .SE(test_se), 
        .CK(clk), .RN(n8998), .Q(BF2I_b_xr_n[20]), .QN(n1685) );
  SDFFRXL BF2I_b00_r_reg_21_ ( .D(n4636), .SI(BF2I_b_xr_n[20]), .SE(test_se), 
        .CK(clk), .RN(n8993), .Q(BF2I_b_xr_n[21]), .QN(n1683) );
  SDFFRXL BF2I_b00_r_reg_22_ ( .D(n4634), .SI(BF2I_b_xr_n[21]), .SE(test_se), 
        .CK(clk), .RN(n8987), .Q(BF2I_b_xr_n[22]), .QN(n1681) );
  SDFFRXL BF2I_b00_r_reg_23_ ( .D(n4632), .SI(BF2I_b_xr_n[22]), .SE(test_se), 
        .CK(clk), .RN(n8987), .Q(BF2I_b_xr_n[23]), .QN(n1679) );
  SDFFRXL BF2I_b00_r_reg_24_ ( .D(n4630), .SI(BF2I_b_xr_n[23]), .SE(test_se), 
        .CK(clk), .RN(n8987), .Q(BF2I_b_xr_n[24]), .QN(n1677) );
  SDFFRXL BF2I_b00_r_reg_25_ ( .D(n4628), .SI(BF2I_b_xr_n[24]), .SE(test_se), 
        .CK(clk), .RN(n8987), .Q(BF2I_b_xr_n[25]), .QN(n1675) );
  SDFFRXL BF2I_b00_r_reg_26_ ( .D(n4626), .SI(BF2I_b_xr_n[25]), .SE(test_se), 
        .CK(clk), .RN(n8987), .Q(BF2I_b_xr_n[26]), .QN(n1673) );
  SDFFRXL BF2I_b00_r_reg_27_ ( .D(n4624), .SI(BF2I_b_xr_n[26]), .SE(test_se), 
        .CK(clk), .RN(n8987), .Q(BF2I_b_xr_n[27]), .QN(n1671) );
  SDFFRXL BF2I_b00_r_reg_28_ ( .D(n4622), .SI(BF2I_b_xr_n[27]), .SE(test_se), 
        .CK(clk), .RN(n8988), .Q(BF2I_b_xr_n[28]), .QN(n1669) );
  SDFFRXL BF2I_b00_r_reg_29_ ( .D(n4620), .SI(BF2I_b_xr_n[28]), .SE(test_se), 
        .CK(clk), .RN(n8988), .Q(BF2I_b_xr_n[29]), .QN(n1667) );
  SDFFRXL BF2I_b00_r_reg_30_ ( .D(n4618), .SI(BF2I_b_xr_n[29]), .SE(test_se), 
        .CK(clk), .RN(n8988), .Q(BF2I_b_xr_n[30]), .QN(n1665) );
  SDFFRXL BF2I_b00_r_reg_31_ ( .D(n4616), .SI(BF2I_b_xr_n[30]), .SE(test_se), 
        .CK(clk), .RN(n8988), .Q(BF2I_b_xr_n[31]), .QN(n1663) );
  SDFFRXL BF2I_b00_i_reg_1_ ( .D(n4612), .SI(BF2I_b_xi_n[0]), .SE(test_se), 
        .CK(clk), .RN(n9046), .Q(BF2I_b_xi_n[1]), .QN(n1659) );
  SDFFRXL BF2I_b00_i_reg_2_ ( .D(n4610), .SI(BF2I_b_xi_n[1]), .SE(test_se), 
        .CK(clk), .RN(n9044), .Q(BF2I_b_xi_n[2]), .QN(n1657) );
  SDFFRXL BF2I_b00_i_reg_3_ ( .D(n4608), .SI(BF2I_b_xi_n[2]), .SE(test_se), 
        .CK(clk), .RN(n9043), .Q(BF2I_b_xi_n[3]), .QN(n1655) );
  SDFFRXL BF2I_b00_i_reg_4_ ( .D(n4606), .SI(BF2I_b_xi_n[3]), .SE(test_se), 
        .CK(clk), .RN(n9041), .Q(BF2I_b_xi_n[4]), .QN(n1653) );
  SDFFRXL BF2I_b00_i_reg_5_ ( .D(n4604), .SI(BF2I_b_xi_n[4]), .SE(test_se), 
        .CK(clk), .RN(n9039), .Q(BF2I_b_xi_n[5]), .QN(n1651) );
  SDFFRXL BF2I_b00_i_reg_6_ ( .D(n4602), .SI(BF2I_b_xi_n[5]), .SE(test_se), 
        .CK(clk), .RN(n9038), .Q(BF2I_b_xi_n[6]), .QN(n1649) );
  SDFFRXL BF2I_b00_i_reg_7_ ( .D(n4600), .SI(BF2I_b_xi_n[6]), .SE(test_se), 
        .CK(clk), .RN(n9036), .Q(BF2I_b_xi_n[7]), .QN(n1647) );
  SDFFRXL BF2I_b00_i_reg_8_ ( .D(n4598), .SI(BF2I_b_xi_n[7]), .SE(test_se), 
        .CK(clk), .RN(n9034), .Q(BF2I_b_xi_n[8]), .QN(n1645) );
  SDFFRXL BF2I_b00_i_reg_9_ ( .D(n4596), .SI(BF2I_b_xi_n[8]), .SE(test_se), 
        .CK(clk), .RN(n9032), .Q(BF2I_b_xi_n[9]), .QN(n1643) );
  SDFFRXL BF2I_b00_i_reg_10_ ( .D(n4594), .SI(BF2I_b_xi_n[9]), .SE(test_se), 
        .CK(clk), .RN(n9031), .Q(BF2I_b_xi_n[10]), .QN(n1641) );
  SDFFRXL BF2I_b00_i_reg_11_ ( .D(n4592), .SI(BF2I_b_xi_n[10]), .SE(test_se), 
        .CK(clk), .RN(n9029), .Q(BF2I_b_xi_n[11]), .QN(n1639) );
  SDFFRXL BF2I_b00_i_reg_12_ ( .D(n4590), .SI(BF2I_b_xi_n[11]), .SE(test_se), 
        .CK(clk), .RN(n9027), .Q(BF2I_b_xi_n[12]), .QN(n1637) );
  SDFFRXL BF2I_b00_i_reg_13_ ( .D(n4588), .SI(BF2I_b_xi_n[12]), .SE(test_se), 
        .CK(clk), .RN(n9026), .Q(BF2I_b_xi_n[13]), .QN(n1635) );
  SDFFRXL BF2I_b00_i_reg_14_ ( .D(n4586), .SI(BF2I_b_xi_n[13]), .SE(test_se), 
        .CK(clk), .RN(n9024), .Q(BF2I_b_xi_n[14]), .QN(n1633) );
  SDFFRXL BF2I_b00_i_reg_15_ ( .D(n4584), .SI(BF2I_b_xi_n[14]), .SE(test_se), 
        .CK(clk), .RN(n9022), .Q(BF2I_b_xi_n[15]), .QN(n1631) );
  SDFFRXL BF2I_b00_i_reg_16_ ( .D(n4582), .SI(BF2I_b_xi_n[15]), .SE(test_se), 
        .CK(clk), .RN(n9022), .Q(BF2I_b_xi_n[16]), .QN(n1629) );
  SDFFRXL BF2I_b00_i_reg_17_ ( .D(n4580), .SI(BF2I_b_xi_n[16]), .SE(test_se), 
        .CK(clk), .RN(n9022), .Q(BF2I_b_xi_n[17]), .QN(n1627) );
  SDFFRXL BF2I_b00_i_reg_18_ ( .D(n4578), .SI(BF2I_b_xi_n[17]), .SE(test_se), 
        .CK(clk), .RN(n9022), .Q(BF2I_b_xi_n[18]), .QN(n1625) );
  SDFFRXL BF2I_b00_i_reg_19_ ( .D(n4576), .SI(BF2I_b_xi_n[18]), .SE(test_se), 
        .CK(clk), .RN(n9022), .Q(BF2I_b_xi_n[19]), .QN(n1623) );
  SDFFRXL BF2I_b00_i_reg_20_ ( .D(n4574), .SI(BF2I_b_xi_n[19]), .SE(test_se), 
        .CK(clk), .RN(n9022), .Q(BF2I_b_xi_n[20]), .QN(n1621) );
  SDFFRXL BF2I_b00_i_reg_21_ ( .D(n4572), .SI(BF2I_b_xi_n[20]), .SE(test_se), 
        .CK(clk), .RN(n9021), .Q(BF2I_b_xi_n[21]), .QN(n1619) );
  SDFFRXL BF2I_b00_i_reg_22_ ( .D(n4570), .SI(BF2I_b_xi_n[21]), .SE(test_se), 
        .CK(clk), .RN(n9021), .Q(BF2I_b_xi_n[22]), .QN(n1617) );
  SDFFRXL BF2I_b00_i_reg_23_ ( .D(n4568), .SI(BF2I_b_xi_n[22]), .SE(test_se), 
        .CK(clk), .RN(n9020), .Q(BF2I_b_xi_n[23]), .QN(n1615) );
  SDFFRXL BF2I_b00_i_reg_24_ ( .D(n4566), .SI(BF2I_b_xi_n[23]), .SE(test_se), 
        .CK(clk), .RN(n9020), .Q(BF2I_b_xi_n[24]), .QN(n1613) );
  SDFFRXL BF2I_b00_i_reg_25_ ( .D(n4564), .SI(BF2I_b_xi_n[24]), .SE(test_se), 
        .CK(clk), .RN(n9020), .Q(BF2I_b_xi_n[25]), .QN(n1611) );
  SDFFRXL BF2I_b00_i_reg_26_ ( .D(n4562), .SI(BF2I_b_xi_n[25]), .SE(test_se), 
        .CK(clk), .RN(n9020), .Q(BF2I_b_xi_n[26]), .QN(n1609) );
  SDFFRXL BF2I_b00_i_reg_27_ ( .D(n4560), .SI(BF2I_b_xi_n[26]), .SE(test_se), 
        .CK(clk), .RN(n9020), .Q(BF2I_b_xi_n[27]), .QN(n1607) );
  SDFFRXL BF2I_b00_i_reg_28_ ( .D(n4558), .SI(BF2I_b_xi_n[27]), .SE(test_se), 
        .CK(clk), .RN(n9021), .Q(BF2I_b_xi_n[28]), .QN(n1605) );
  SDFFRXL BF2I_b00_i_reg_29_ ( .D(n4556), .SI(BF2I_b_xi_n[28]), .SE(test_se), 
        .CK(clk), .RN(n9021), .Q(BF2I_b_xi_n[29]), .QN(n1603) );
  SDFFRXL BF2I_b00_i_reg_30_ ( .D(n4554), .SI(BF2I_b_xi_n[29]), .SE(test_se), 
        .CK(clk), .RN(n9021), .Q(BF2I_b_xi_n[30]), .QN(n1601) );
  SDFFRXL BF2I_b00_i_reg_31_ ( .D(n4552), .SI(BF2I_b_xi_n[30]), .SE(test_se), 
        .CK(clk), .RN(n9021), .Q(BF2I_b_xi_n[31]), .QN(n1599) );
  SDFFRXL d32_reg_17_ ( .D(n4950), .SI(d32[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d32[17]) );
  SDFFRXL d32_reg_18_ ( .D(n4949), .SI(d32[17]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d32[18]) );
  SDFFRXL d32_reg_19_ ( .D(n4948), .SI(d32[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d32[19]) );
  SDFFRXL d32_reg_20_ ( .D(n4947), .SI(d32[19]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d32[20]) );
  SDFFRXL d32_reg_21_ ( .D(n4946), .SI(d32[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d32[21]) );
  SDFFRXL d32_reg_22_ ( .D(n4945), .SI(d32[21]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d32[22]) );
  SDFFRXL d32_reg_23_ ( .D(n4944), .SI(d32[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d32[23]) );
  SDFFRXL d32_reg_24_ ( .D(n4943), .SI(d32[23]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d32[24]) );
  SDFFRXL d32_reg_25_ ( .D(n4942), .SI(d32[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d32[25]) );
  SDFFRXL d32_reg_26_ ( .D(n4941), .SI(d32[25]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d32[26]) );
  SDFFRXL d32_reg_27_ ( .D(n4940), .SI(d32[26]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d32[27]) );
  SDFFRXL d32_reg_28_ ( .D(n4939), .SI(d32[27]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d32[28]) );
  SDFFRXL d32_reg_29_ ( .D(n4938), .SI(d32[28]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d32[29]) );
  SDFFRXL d32_reg_30_ ( .D(n4937), .SI(d32[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d32[30]) );
  SDFFRXL d01_reg_35_ ( .D(n6064), .SI(d01[34]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d01[35]), .QN(n3079) );
  SDFFRXL d01_reg_34_ ( .D(n6062), .SI(d01[33]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d01[34]), .QN(n3078) );
  SDFFRXL d01_reg_33_ ( .D(n6061), .SI(d01[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d01[33]), .QN(n3077) );
  SDFFRXL d01_reg_32_ ( .D(n6060), .SI(d01[31]), .SE(test_se), .CK(clk), .RN(
        n8933), .Q(d01[32]), .QN(n3076) );
  SDFFRXL d01_reg_31_ ( .D(n6059), .SI(d01[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d01[31]), .QN(n3075) );
  SDFFRXL d01_reg_30_ ( .D(n6058), .SI(d01[29]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d01[30]), .QN(n3074) );
  SDFFRXL d01_reg_29_ ( .D(n6057), .SI(d01[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d01[29]), .QN(n3073) );
  SDFFRXL d01_reg_28_ ( .D(n6056), .SI(d01[27]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d01[28]), .QN(n3072) );
  SDFFRXL d01_reg_27_ ( .D(n6055), .SI(d01[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d01[27]), .QN(n3071) );
  SDFFRXL d01_reg_26_ ( .D(n6054), .SI(d01[25]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d01[26]), .QN(n30701) );
  SDFFRXL d01_reg_25_ ( .D(n6053), .SI(d01[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d01[25]), .QN(n3069) );
  SDFFRXL d01_reg_24_ ( .D(n6052), .SI(d01[23]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d01[24]), .QN(n3068) );
  SDFFRXL d01_reg_23_ ( .D(n6051), .SI(d01[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d01[23]), .QN(n3067) );
  SDFFRXL d01_reg_1_ ( .D(n6029), .SI(n6191), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d01[1]) );
  SDFFRXL d02_reg_0_ ( .D(n5992), .SI(d01[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d02[0]) );
  SDFFRXL d03_reg_0_ ( .D(n5956), .SI(d02[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d03[0]) );
  SDFFRXL d04_reg_0_ ( .D(n5920), .SI(d03[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d04[0]) );
  SDFFRXL d05_reg_1_ ( .D(n5885), .SI(d05[0]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d05[1]) );
  SDFFRXL d06_reg_1_ ( .D(n5849), .SI(d06[0]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d06[1]) );
  SDFFRXL d07_reg_2_ ( .D(n5814), .SI(d07[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d07[2]) );
  SDFFRXL d08_reg_0_ ( .D(n5776), .SI(d07[35]), .SE(test_se), .CK(clk), .RN(
        n9126), .Q(d08[0]) );
  SDFFRXL d09_reg_1_ ( .D(n5741), .SI(d09[0]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d09[1]) );
  SDFFRXL d10_reg_1_ ( .D(n5705), .SI(d10[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d10[1]) );
  SDFFRXL d11_reg_2_ ( .D(n5670), .SI(d11[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d11[2]) );
  SDFFRXL d12_reg_1_ ( .D(n5633), .SI(d12[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d12[1]) );
  SDFFRXL d13_reg_2_ ( .D(n5598), .SI(d13[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d13[2]) );
  SDFFRXL d14_reg_1_ ( .D(n5561), .SI(d14[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d14[1]) );
  SDFFRXL d15_reg_0_ ( .D(n5524), .SI(d14[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d15[0]) );
  SDFFRXL d16_reg_0_ ( .D(n5488), .SI(d15[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d16[0]) );
  SDFFRXL d17_reg_1_ ( .D(n5453), .SI(d17[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d17[1]) );
  SDFFRXL d18_reg_2_ ( .D(n5418), .SI(d18[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d18[2]) );
  SDFFRXL d19_reg_1_ ( .D(n5381), .SI(d19[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d19[1]) );
  SDFFRXL d20_reg_2_ ( .D(n5346), .SI(d20[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d20[2]) );
  SDFFRXL d21_reg_1_ ( .D(n5309), .SI(d21[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d21[1]) );
  SDFFRXL d22_reg_1_ ( .D(n5273), .SI(d22[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d22[1]) );
  SDFFRXL d23_reg_0_ ( .D(n5236), .SI(d22[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d23[0]) );
  SDFFRXL d24_reg_2_ ( .D(n5202), .SI(d24[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d24[2]) );
  SDFFRXL d25_reg_1_ ( .D(n5165), .SI(d25[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d25[1]) );
  SDFFRXL d26_reg_1_ ( .D(n5129), .SI(d26[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d26[1]) );
  SDFFRXL d27_reg_0_ ( .D(n5092), .SI(d26[35]), .SE(test_se), .CK(clk), .RN(
        n9125), .Q(d27[0]) );
  SDFFRXL d28_reg_0_ ( .D(n5056), .SI(d27[35]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d28[0]) );
  SDFFRXL d29_reg_0_ ( .D(n5020), .SI(d28[35]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d29[0]) );
  SDFFRXL d30_reg_1_ ( .D(n5018), .SI(d30[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d30[1]) );
  SDFFRXL d01_reg_22_ ( .D(n6050), .SI(d01[21]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d01[22]) );
  SDFFRXL d01_reg_21_ ( .D(n6049), .SI(d01[20]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d01[21]) );
  SDFFRXL d01_reg_20_ ( .D(n6048), .SI(d01[19]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d01[20]) );
  SDFFRXL d01_reg_19_ ( .D(n6047), .SI(d01[18]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d01[19]) );
  SDFFRXL d01_reg_18_ ( .D(n6046), .SI(d01[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d01[18]) );
  SDFFRXL d01_reg_17_ ( .D(n6045), .SI(d01[16]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d01[17]) );
  SDFFRXL d01_reg_16_ ( .D(n6044), .SI(d01[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d01[16]) );
  SDFFRXL d01_reg_15_ ( .D(n6043), .SI(d01[14]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d01[15]) );
  SDFFRXL d01_reg_14_ ( .D(n6042), .SI(d01[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d01[14]) );
  SDFFRXL d01_reg_13_ ( .D(n6041), .SI(d01[12]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d01[13]) );
  SDFFRXL d01_reg_12_ ( .D(n6040), .SI(d01[11]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d01[12]) );
  SDFFRXL d01_reg_11_ ( .D(n6039), .SI(d01[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d01[11]) );
  SDFFRXL d01_reg_10_ ( .D(n6038), .SI(d01[9]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d01[10]) );
  SDFFRXL d01_reg_9_ ( .D(n6037), .SI(d01[8]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d01[9]) );
  SDFFRXL d01_reg_8_ ( .D(n6036), .SI(d01[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d01[8]) );
  SDFFRXL d01_reg_7_ ( .D(n6035), .SI(d01[6]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d01[7]) );
  SDFFRXL d01_reg_6_ ( .D(n6034), .SI(d01[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d01[6]) );
  SDFFRXL d01_reg_5_ ( .D(n6033), .SI(d01[4]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d01[5]) );
  SDFFRXL d01_reg_4_ ( .D(n6032), .SI(d01[3]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d01[4]) );
  SDFFRXL d01_reg_3_ ( .D(n6031), .SI(d01[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d01[3]) );
  SDFFRXL d01_reg_2_ ( .D(n6030), .SI(d01[1]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d01[2]) );
  SDFFRXL d02_reg_35_ ( .D(n6027), .SI(d02[34]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d02[35]) );
  SDFFRXL d02_reg_34_ ( .D(n6026), .SI(d02[33]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d02[34]) );
  SDFFRXL d02_reg_33_ ( .D(n6025), .SI(d02[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d02[33]) );
  SDFFRXL d02_reg_32_ ( .D(n6024), .SI(d02[31]), .SE(test_se), .CK(clk), .RN(
        n8933), .Q(d02[32]) );
  SDFFRXL d02_reg_31_ ( .D(n6023), .SI(d02[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d02[31]) );
  SDFFRXL d02_reg_30_ ( .D(n6022), .SI(d02[29]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d02[30]) );
  SDFFRXL d02_reg_29_ ( .D(n6021), .SI(d02[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d02[29]) );
  SDFFRXL d02_reg_28_ ( .D(n6020), .SI(d02[27]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d02[28]) );
  SDFFRXL d02_reg_27_ ( .D(n6019), .SI(d02[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d02[27]) );
  SDFFRXL d02_reg_26_ ( .D(n6018), .SI(d02[25]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d02[26]) );
  SDFFRXL d02_reg_25_ ( .D(n6017), .SI(d02[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d02[25]) );
  SDFFRXL d02_reg_24_ ( .D(n6016), .SI(d02[23]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d02[24]) );
  SDFFRXL d02_reg_23_ ( .D(n6015), .SI(d02[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d02[23]) );
  SDFFRXL d02_reg_22_ ( .D(n6014), .SI(d02[21]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d02[22]) );
  SDFFRXL d02_reg_21_ ( .D(n6013), .SI(d02[20]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d02[21]) );
  SDFFRXL d02_reg_20_ ( .D(n6012), .SI(d02[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d02[20]) );
  SDFFRXL d02_reg_19_ ( .D(n6011), .SI(d02[18]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d02[19]) );
  SDFFRXL d02_reg_18_ ( .D(n6010), .SI(d02[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d02[18]) );
  SDFFRXL d02_reg_17_ ( .D(n6009), .SI(d02[16]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d02[17]) );
  SDFFRXL d02_reg_16_ ( .D(n6008), .SI(d02[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d02[16]) );
  SDFFRXL d02_reg_15_ ( .D(n6007), .SI(d02[14]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d02[15]) );
  SDFFRXL d02_reg_14_ ( .D(n6006), .SI(d02[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d02[14]) );
  SDFFRXL d02_reg_13_ ( .D(n6005), .SI(d02[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d02[13]) );
  SDFFRXL d02_reg_12_ ( .D(n6004), .SI(d02[11]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d02[12]) );
  SDFFRXL d02_reg_11_ ( .D(n6003), .SI(d02[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d02[11]) );
  SDFFRXL d02_reg_10_ ( .D(n6002), .SI(d02[9]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d02[10]) );
  SDFFRXL d02_reg_9_ ( .D(n6001), .SI(d02[8]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d02[9]) );
  SDFFRXL d02_reg_8_ ( .D(n6000), .SI(d02[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d02[8]) );
  SDFFRXL d02_reg_7_ ( .D(n5999), .SI(d02[6]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d02[7]) );
  SDFFRXL d02_reg_6_ ( .D(n5998), .SI(d02[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d02[6]) );
  SDFFRXL d02_reg_5_ ( .D(n5997), .SI(d02[4]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d02[5]) );
  SDFFRXL d02_reg_4_ ( .D(n5996), .SI(d02[3]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d02[4]) );
  SDFFRXL d02_reg_3_ ( .D(n5995), .SI(d02[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d02[3]) );
  SDFFRXL d02_reg_2_ ( .D(n5994), .SI(d02[1]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d02[2]) );
  SDFFRXL d02_reg_1_ ( .D(n5993), .SI(d02[0]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d02[1]) );
  SDFFRXL d03_reg_35_ ( .D(n5991), .SI(d03[34]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d03[35]) );
  SDFFRXL d03_reg_34_ ( .D(n5990), .SI(d03[33]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d03[34]) );
  SDFFRXL d03_reg_33_ ( .D(n5989), .SI(d03[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d03[33]) );
  SDFFRXL d03_reg_32_ ( .D(n5988), .SI(d03[31]), .SE(test_se), .CK(clk), .RN(
        n8933), .Q(d03[32]) );
  SDFFRXL d03_reg_31_ ( .D(n5987), .SI(d03[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d03[31]) );
  SDFFRXL d03_reg_30_ ( .D(n5986), .SI(d03[29]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d03[30]) );
  SDFFRXL d03_reg_29_ ( .D(n5985), .SI(d03[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d03[29]) );
  SDFFRXL d03_reg_28_ ( .D(n5984), .SI(d03[27]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d03[28]) );
  SDFFRXL d03_reg_27_ ( .D(n5983), .SI(d03[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d03[27]) );
  SDFFRXL d03_reg_26_ ( .D(n5982), .SI(d03[25]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d03[26]) );
  SDFFRXL d03_reg_25_ ( .D(n5981), .SI(d03[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d03[25]) );
  SDFFRXL d03_reg_24_ ( .D(n5980), .SI(d03[23]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d03[24]) );
  SDFFRXL d03_reg_23_ ( .D(n5979), .SI(d03[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d03[23]) );
  SDFFRXL d03_reg_22_ ( .D(n5978), .SI(d03[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d03[22]) );
  SDFFRXL d03_reg_21_ ( .D(n5977), .SI(d03[20]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d03[21]) );
  SDFFRXL d03_reg_20_ ( .D(n5976), .SI(d03[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d03[20]) );
  SDFFRXL d03_reg_19_ ( .D(n5975), .SI(d03[18]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d03[19]) );
  SDFFRXL d03_reg_18_ ( .D(n5974), .SI(d03[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d03[18]) );
  SDFFRXL d03_reg_17_ ( .D(n5973), .SI(d03[16]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d03[17]) );
  SDFFRXL d03_reg_16_ ( .D(n5972), .SI(d03[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d03[16]) );
  SDFFRXL d03_reg_15_ ( .D(n5971), .SI(d03[14]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d03[15]) );
  SDFFRXL d03_reg_14_ ( .D(n5970), .SI(d03[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d03[14]) );
  SDFFRXL d03_reg_13_ ( .D(n5969), .SI(d03[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d03[13]) );
  SDFFRXL d03_reg_12_ ( .D(n5968), .SI(d03[11]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d03[12]) );
  SDFFRXL d03_reg_11_ ( .D(n5967), .SI(d03[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d03[11]) );
  SDFFRXL d03_reg_10_ ( .D(n5966), .SI(d03[9]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d03[10]) );
  SDFFRXL d03_reg_9_ ( .D(n5965), .SI(d03[8]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d03[9]) );
  SDFFRXL d03_reg_8_ ( .D(n5964), .SI(d03[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d03[8]) );
  SDFFRXL d03_reg_7_ ( .D(n5963), .SI(d03[6]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d03[7]) );
  SDFFRXL d03_reg_6_ ( .D(n5962), .SI(d03[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d03[6]) );
  SDFFRXL d03_reg_5_ ( .D(n5961), .SI(d03[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d03[5]) );
  SDFFRXL d03_reg_4_ ( .D(n5960), .SI(d03[3]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d03[4]) );
  SDFFRXL d03_reg_3_ ( .D(n5959), .SI(d03[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d03[3]) );
  SDFFRXL d03_reg_2_ ( .D(n5958), .SI(d03[1]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d03[2]) );
  SDFFRXL d03_reg_1_ ( .D(n5957), .SI(d03[0]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d03[1]) );
  SDFFRXL d04_reg_35_ ( .D(n5955), .SI(d04[34]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d04[35]) );
  SDFFRXL d04_reg_34_ ( .D(n5954), .SI(d04[33]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d04[34]) );
  SDFFRXL d04_reg_33_ ( .D(n5953), .SI(d04[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d04[33]) );
  SDFFRXL d04_reg_32_ ( .D(n5952), .SI(d04[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d04[32]) );
  SDFFRXL d04_reg_31_ ( .D(n5951), .SI(d04[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d04[31]) );
  SDFFRXL d04_reg_30_ ( .D(n5950), .SI(d04[29]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d04[30]) );
  SDFFRXL d04_reg_29_ ( .D(n5949), .SI(d04[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d04[29]) );
  SDFFRXL d04_reg_28_ ( .D(n5948), .SI(d04[27]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d04[28]) );
  SDFFRXL d04_reg_27_ ( .D(n5947), .SI(d04[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d04[27]) );
  SDFFRXL d04_reg_26_ ( .D(n5946), .SI(d04[25]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d04[26]) );
  SDFFRXL d04_reg_25_ ( .D(n5945), .SI(d04[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d04[25]) );
  SDFFRXL d04_reg_24_ ( .D(n5944), .SI(d04[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d04[24]) );
  SDFFRXL d04_reg_23_ ( .D(n5943), .SI(d04[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d04[23]) );
  SDFFRXL d04_reg_22_ ( .D(n5942), .SI(d04[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d04[22]) );
  SDFFRXL d04_reg_21_ ( .D(n5941), .SI(d04[20]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d04[21]) );
  SDFFRXL d04_reg_20_ ( .D(n5940), .SI(d04[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d04[20]) );
  SDFFRXL d04_reg_19_ ( .D(n5939), .SI(d04[18]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d04[19]) );
  SDFFRXL d04_reg_18_ ( .D(n5938), .SI(d04[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d04[18]) );
  SDFFRXL d04_reg_17_ ( .D(n5937), .SI(d04[16]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d04[17]) );
  SDFFRXL d04_reg_16_ ( .D(n5936), .SI(d04[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d04[16]) );
  SDFFRXL d04_reg_15_ ( .D(n5935), .SI(d04[14]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d04[15]) );
  SDFFRXL d04_reg_14_ ( .D(n5934), .SI(d04[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d04[14]) );
  SDFFRXL d04_reg_13_ ( .D(n5933), .SI(d04[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d04[13]) );
  SDFFRXL d04_reg_12_ ( .D(n5932), .SI(d04[11]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d04[12]) );
  SDFFRXL d04_reg_11_ ( .D(n5931), .SI(d04[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d04[11]) );
  SDFFRXL d04_reg_10_ ( .D(n5930), .SI(d04[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d04[10]) );
  SDFFRXL d04_reg_9_ ( .D(n5929), .SI(d04[8]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d04[9]) );
  SDFFRXL d04_reg_8_ ( .D(n5928), .SI(d04[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d04[8]) );
  SDFFRXL d04_reg_7_ ( .D(n5927), .SI(d04[6]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d04[7]) );
  SDFFRXL d04_reg_6_ ( .D(n5926), .SI(d04[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d04[6]) );
  SDFFRXL d04_reg_5_ ( .D(n5925), .SI(d04[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d04[5]) );
  SDFFRXL d04_reg_4_ ( .D(n5924), .SI(d04[3]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d04[4]) );
  SDFFRXL d04_reg_3_ ( .D(n5923), .SI(d04[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d04[3]) );
  SDFFRXL d04_reg_2_ ( .D(n5922), .SI(d04[1]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d04[2]) );
  SDFFRXL d04_reg_1_ ( .D(n5921), .SI(d04[0]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d04[1]) );
  SDFFRXL d05_reg_35_ ( .D(n5919), .SI(d05[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d05[35]) );
  SDFFRXL d05_reg_34_ ( .D(n5918), .SI(d05[33]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d05[34]) );
  SDFFRXL d05_reg_33_ ( .D(n5917), .SI(d05[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d05[33]) );
  SDFFRXL d05_reg_32_ ( .D(n5916), .SI(d05[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d05[32]) );
  SDFFRXL d05_reg_31_ ( .D(n5915), .SI(d05[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d05[31]) );
  SDFFRXL d05_reg_30_ ( .D(n5914), .SI(d05[29]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d05[30]) );
  SDFFRXL d05_reg_29_ ( .D(n5913), .SI(d05[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d05[29]) );
  SDFFRXL d05_reg_28_ ( .D(n5912), .SI(d05[27]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d05[28]) );
  SDFFRXL d05_reg_27_ ( .D(n5911), .SI(d05[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d05[27]) );
  SDFFRXL d05_reg_26_ ( .D(n5910), .SI(d05[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d05[26]) );
  SDFFRXL d05_reg_25_ ( .D(n5909), .SI(d05[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d05[25]) );
  SDFFRXL d05_reg_24_ ( .D(n5908), .SI(d05[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d05[24]) );
  SDFFRXL d05_reg_23_ ( .D(n5907), .SI(d05[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d05[23]) );
  SDFFRXL d05_reg_22_ ( .D(n5906), .SI(d05[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d05[22]) );
  SDFFRXL d05_reg_21_ ( .D(n5905), .SI(d05[20]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d05[21]) );
  SDFFRXL d05_reg_20_ ( .D(n5904), .SI(d05[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d05[20]) );
  SDFFRXL d05_reg_19_ ( .D(n5903), .SI(d05[18]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d05[19]) );
  SDFFRXL d05_reg_18_ ( .D(n5902), .SI(d05[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d05[18]) );
  SDFFRXL d05_reg_17_ ( .D(n5901), .SI(d05[16]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d05[17]) );
  SDFFRXL d05_reg_16_ ( .D(n5900), .SI(d05[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d05[16]) );
  SDFFRXL d05_reg_15_ ( .D(n5899), .SI(d05[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d05[15]) );
  SDFFRXL d05_reg_14_ ( .D(n5898), .SI(d05[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d05[14]) );
  SDFFRXL d05_reg_13_ ( .D(n5897), .SI(d05[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d05[13]) );
  SDFFRXL d05_reg_12_ ( .D(n5896), .SI(d05[11]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d05[12]) );
  SDFFRXL d05_reg_11_ ( .D(n5895), .SI(d05[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d05[11]) );
  SDFFRXL d05_reg_10_ ( .D(n5894), .SI(d05[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d05[10]) );
  SDFFRXL d05_reg_9_ ( .D(n5893), .SI(d05[8]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d05[9]) );
  SDFFRXL d05_reg_8_ ( .D(n5892), .SI(d05[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d05[8]) );
  SDFFRXL d05_reg_7_ ( .D(n5891), .SI(d05[6]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d05[7]) );
  SDFFRXL d05_reg_6_ ( .D(n5890), .SI(d05[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d05[6]) );
  SDFFRXL d05_reg_5_ ( .D(n5889), .SI(d05[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d05[5]) );
  SDFFRXL d05_reg_4_ ( .D(n5888), .SI(d05[3]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d05[4]) );
  SDFFRXL d05_reg_3_ ( .D(n5887), .SI(d05[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d05[3]) );
  SDFFRXL d05_reg_2_ ( .D(n5886), .SI(d05[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d05[2]) );
  SDFFRXL d06_reg_35_ ( .D(n5883), .SI(d06[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d06[35]) );
  SDFFRXL d06_reg_34_ ( .D(n5882), .SI(d06[33]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d06[34]) );
  SDFFRXL d06_reg_33_ ( .D(n5881), .SI(d06[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d06[33]) );
  SDFFRXL d06_reg_32_ ( .D(n5880), .SI(d06[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d06[32]) );
  SDFFRXL d06_reg_31_ ( .D(n5879), .SI(d06[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d06[31]) );
  SDFFRXL d06_reg_30_ ( .D(n5878), .SI(d06[29]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d06[30]) );
  SDFFRXL d06_reg_29_ ( .D(n5877), .SI(d06[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d06[29]) );
  SDFFRXL d06_reg_28_ ( .D(n5876), .SI(d06[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d06[28]) );
  SDFFRXL d06_reg_27_ ( .D(n5875), .SI(d06[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d06[27]) );
  SDFFRXL d06_reg_26_ ( .D(n5874), .SI(d06[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d06[26]) );
  SDFFRXL d06_reg_25_ ( .D(n5873), .SI(d06[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d06[25]) );
  SDFFRXL d06_reg_24_ ( .D(n5872), .SI(d06[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d06[24]) );
  SDFFRXL d06_reg_23_ ( .D(n5871), .SI(d06[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d06[23]) );
  SDFFRXL d06_reg_22_ ( .D(n5870), .SI(d06[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d06[22]) );
  SDFFRXL d06_reg_21_ ( .D(n5869), .SI(d06[20]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d06[21]) );
  SDFFRXL d06_reg_20_ ( .D(n5868), .SI(d06[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d06[20]) );
  SDFFRXL d06_reg_19_ ( .D(n5867), .SI(d06[18]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d06[19]) );
  SDFFRXL d06_reg_18_ ( .D(n5866), .SI(d06[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d06[18]) );
  SDFFRXL d06_reg_17_ ( .D(n5865), .SI(d06[16]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d06[17]) );
  SDFFRXL d06_reg_16_ ( .D(n5864), .SI(d06[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d06[16]) );
  SDFFRXL d06_reg_15_ ( .D(n5863), .SI(d06[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d06[15]) );
  SDFFRXL d06_reg_14_ ( .D(n5862), .SI(d06[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d06[14]) );
  SDFFRXL d06_reg_13_ ( .D(n5861), .SI(d06[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d06[13]) );
  SDFFRXL d06_reg_12_ ( .D(n5860), .SI(d06[11]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d06[12]) );
  SDFFRXL d06_reg_11_ ( .D(n5859), .SI(d06[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d06[11]) );
  SDFFRXL d06_reg_10_ ( .D(n5858), .SI(d06[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d06[10]) );
  SDFFRXL d06_reg_9_ ( .D(n5857), .SI(d06[8]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d06[9]) );
  SDFFRXL d06_reg_8_ ( .D(n5856), .SI(d06[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d06[8]) );
  SDFFRXL d06_reg_7_ ( .D(n5855), .SI(d06[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d06[7]) );
  SDFFRXL d06_reg_6_ ( .D(n5854), .SI(d06[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d06[6]) );
  SDFFRXL d06_reg_5_ ( .D(n5853), .SI(d06[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d06[5]) );
  SDFFRXL d06_reg_4_ ( .D(n5852), .SI(d06[3]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d06[4]) );
  SDFFRXL d06_reg_3_ ( .D(n5851), .SI(d06[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d06[3]) );
  SDFFRXL d06_reg_2_ ( .D(n5850), .SI(d06[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d06[2]) );
  SDFFRXL d07_reg_35_ ( .D(n5847), .SI(d07[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d07[35]) );
  SDFFRXL d07_reg_34_ ( .D(n5846), .SI(d07[33]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d07[34]) );
  SDFFRXL d07_reg_33_ ( .D(n5845), .SI(d07[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d07[33]) );
  SDFFRXL d07_reg_32_ ( .D(n5844), .SI(d07[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d07[32]) );
  SDFFRXL d07_reg_31_ ( .D(n5843), .SI(d07[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d07[31]) );
  SDFFRXL d07_reg_30_ ( .D(n5842), .SI(d07[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d07[30]) );
  SDFFRXL d07_reg_29_ ( .D(n5841), .SI(d07[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d07[29]) );
  SDFFRXL d07_reg_28_ ( .D(n5840), .SI(d07[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d07[28]) );
  SDFFRXL d07_reg_27_ ( .D(n5839), .SI(d07[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d07[27]) );
  SDFFRXL d07_reg_26_ ( .D(n5838), .SI(d07[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d07[26]) );
  SDFFRXL d07_reg_25_ ( .D(n5837), .SI(d07[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d07[25]) );
  SDFFRXL d07_reg_24_ ( .D(n5836), .SI(d07[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d07[24]) );
  SDFFRXL d07_reg_23_ ( .D(n5835), .SI(d07[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d07[23]) );
  SDFFRXL d07_reg_22_ ( .D(n5834), .SI(d07[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d07[22]) );
  SDFFRXL d07_reg_21_ ( .D(n5833), .SI(d07[20]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d07[21]) );
  SDFFRXL d07_reg_20_ ( .D(n5832), .SI(d07[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d07[20]) );
  SDFFRXL d07_reg_19_ ( .D(n5831), .SI(d07[18]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d07[19]) );
  SDFFRXL d07_reg_18_ ( .D(n5830), .SI(d07[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d07[18]) );
  SDFFRXL d07_reg_17_ ( .D(n5829), .SI(d07[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d07[17]) );
  SDFFRXL d07_reg_16_ ( .D(n5828), .SI(d07[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d07[16]) );
  SDFFRXL d07_reg_15_ ( .D(n5827), .SI(d07[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d07[15]) );
  SDFFRXL d07_reg_14_ ( .D(n5826), .SI(d07[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d07[14]) );
  SDFFRXL d07_reg_13_ ( .D(n5825), .SI(d07[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d07[13]) );
  SDFFRXL d07_reg_12_ ( .D(n5824), .SI(d07[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d07[12]) );
  SDFFRXL d07_reg_11_ ( .D(n5823), .SI(d07[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d07[11]) );
  SDFFRXL d07_reg_10_ ( .D(n5822), .SI(d07[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d07[10]) );
  SDFFRXL d07_reg_9_ ( .D(n5821), .SI(d07[8]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d07[9]) );
  SDFFRXL d07_reg_8_ ( .D(n5820), .SI(d07[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d07[8]) );
  SDFFRXL d07_reg_7_ ( .D(n5819), .SI(d07[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d07[7]) );
  SDFFRXL d07_reg_6_ ( .D(n5818), .SI(d07[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d07[6]) );
  SDFFRXL d07_reg_5_ ( .D(n5817), .SI(d07[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d07[5]) );
  SDFFRXL d07_reg_4_ ( .D(n5816), .SI(d07[3]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d07[4]) );
  SDFFRXL d07_reg_3_ ( .D(n5815), .SI(d07[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d07[3]) );
  SDFFRXL d08_reg_35_ ( .D(n5811), .SI(d08[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d08[35]) );
  SDFFRXL d08_reg_34_ ( .D(n5810), .SI(d08[33]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d08[34]) );
  SDFFRXL d08_reg_33_ ( .D(n5809), .SI(d08[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d08[33]) );
  SDFFRXL d08_reg_32_ ( .D(n5808), .SI(d08[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d08[32]) );
  SDFFRXL d08_reg_31_ ( .D(n5807), .SI(d08[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d08[31]) );
  SDFFRXL d08_reg_30_ ( .D(n5806), .SI(d08[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d08[30]) );
  SDFFRXL d08_reg_29_ ( .D(n5805), .SI(d08[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d08[29]) );
  SDFFRXL d08_reg_28_ ( .D(n5804), .SI(d08[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d08[28]) );
  SDFFRXL d08_reg_27_ ( .D(n5803), .SI(d08[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d08[27]) );
  SDFFRXL d08_reg_26_ ( .D(n5802), .SI(d08[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d08[26]) );
  SDFFRXL d08_reg_25_ ( .D(n5801), .SI(d08[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d08[25]) );
  SDFFRXL d08_reg_24_ ( .D(n5800), .SI(d08[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d08[24]) );
  SDFFRXL d08_reg_23_ ( .D(n5799), .SI(d08[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d08[23]) );
  SDFFRXL d08_reg_22_ ( .D(n5798), .SI(d08[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d08[22]) );
  SDFFRXL d08_reg_21_ ( .D(n5797), .SI(d08[20]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d08[21]) );
  SDFFRXL d08_reg_20_ ( .D(n5796), .SI(d08[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d08[20]) );
  SDFFRXL d08_reg_19_ ( .D(n5795), .SI(d08[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d08[19]) );
  SDFFRXL d08_reg_18_ ( .D(n5794), .SI(d08[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d08[18]) );
  SDFFRXL d08_reg_17_ ( .D(n5793), .SI(d08[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d08[17]) );
  SDFFRXL d08_reg_16_ ( .D(n5792), .SI(d08[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d08[16]) );
  SDFFRXL d08_reg_15_ ( .D(n5791), .SI(d08[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d08[15]) );
  SDFFRXL d08_reg_14_ ( .D(n5790), .SI(d08[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d08[14]) );
  SDFFRXL d08_reg_13_ ( .D(n5789), .SI(d08[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d08[13]) );
  SDFFRXL d08_reg_12_ ( .D(n5788), .SI(d08[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d08[12]) );
  SDFFRXL d08_reg_11_ ( .D(n5787), .SI(d08[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d08[11]) );
  SDFFRXL d08_reg_10_ ( .D(n5786), .SI(d08[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d08[10]) );
  SDFFRXL d08_reg_9_ ( .D(n5785), .SI(d08[8]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d08[9]) );
  SDFFRXL d08_reg_8_ ( .D(n5784), .SI(d08[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d08[8]) );
  SDFFRXL d08_reg_7_ ( .D(n5783), .SI(d08[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d08[7]) );
  SDFFRXL d08_reg_6_ ( .D(n5782), .SI(d08[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d08[6]) );
  SDFFRXL d08_reg_5_ ( .D(n5781), .SI(d08[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d08[5]) );
  SDFFRXL d08_reg_4_ ( .D(n5780), .SI(d08[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d08[4]) );
  SDFFRXL d08_reg_3_ ( .D(n5779), .SI(d08[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d08[3]) );
  SDFFRXL d08_reg_2_ ( .D(n5778), .SI(d08[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d08[2]) );
  SDFFRXL d08_reg_1_ ( .D(n5777), .SI(d08[0]), .SE(test_se), .CK(clk), .RN(
        n9124), .Q(d08[1]) );
  SDFFRXL d09_reg_35_ ( .D(n5775), .SI(d09[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d09[35]) );
  SDFFRXL d09_reg_34_ ( .D(n5774), .SI(d09[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d09[34]) );
  SDFFRXL d09_reg_33_ ( .D(n5773), .SI(d09[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d09[33]) );
  SDFFRXL d09_reg_32_ ( .D(n5772), .SI(d09[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d09[32]) );
  SDFFRXL d09_reg_31_ ( .D(n5771), .SI(d09[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d09[31]) );
  SDFFRXL d09_reg_30_ ( .D(n5770), .SI(d09[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d09[30]) );
  SDFFRXL d09_reg_29_ ( .D(n5769), .SI(d09[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d09[29]) );
  SDFFRXL d09_reg_28_ ( .D(n5768), .SI(d09[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d09[28]) );
  SDFFRXL d09_reg_27_ ( .D(n5767), .SI(d09[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d09[27]) );
  SDFFRXL d09_reg_26_ ( .D(n5766), .SI(d09[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d09[26]) );
  SDFFRXL d09_reg_25_ ( .D(n5765), .SI(d09[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d09[25]) );
  SDFFRXL d09_reg_24_ ( .D(n5764), .SI(d09[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d09[24]) );
  SDFFRXL d09_reg_23_ ( .D(n5763), .SI(d09[22]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d09[23]) );
  SDFFRXL d09_reg_22_ ( .D(n5762), .SI(d09[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d09[22]) );
  SDFFRXL d09_reg_21_ ( .D(n5761), .SI(d09[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d09[21]) );
  SDFFRXL d09_reg_20_ ( .D(n5760), .SI(d09[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d09[20]) );
  SDFFRXL d09_reg_19_ ( .D(n5759), .SI(d09[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d09[19]) );
  SDFFRXL d09_reg_18_ ( .D(n5758), .SI(d09[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d09[18]) );
  SDFFRXL d09_reg_17_ ( .D(n5757), .SI(d09[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d09[17]) );
  SDFFRXL d09_reg_16_ ( .D(n5756), .SI(d09[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d09[16]) );
  SDFFRXL d09_reg_15_ ( .D(n5755), .SI(d09[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d09[15]) );
  SDFFRXL d09_reg_14_ ( .D(n5754), .SI(d09[13]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d09[14]) );
  SDFFRXL d09_reg_13_ ( .D(n5753), .SI(d09[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d09[13]) );
  SDFFRXL d09_reg_12_ ( .D(n5752), .SI(d09[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d09[12]) );
  SDFFRXL d09_reg_11_ ( .D(n5751), .SI(d09[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d09[11]) );
  SDFFRXL d09_reg_10_ ( .D(n5750), .SI(d09[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d09[10]) );
  SDFFRXL d09_reg_9_ ( .D(n5749), .SI(d09[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d09[9]) );
  SDFFRXL d09_reg_8_ ( .D(n5748), .SI(d09[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d09[8]) );
  SDFFRXL d09_reg_7_ ( .D(n5747), .SI(d09[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d09[7]) );
  SDFFRXL d09_reg_6_ ( .D(n5746), .SI(d09[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d09[6]) );
  SDFFRXL d09_reg_5_ ( .D(n5745), .SI(d09[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d09[5]) );
  SDFFRXL d09_reg_4_ ( .D(n5744), .SI(d09[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d09[4]) );
  SDFFRXL d09_reg_3_ ( .D(n5743), .SI(d09[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d09[3]) );
  SDFFRXL d09_reg_2_ ( .D(n5742), .SI(d09[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d09[2]) );
  SDFFRXL d10_reg_35_ ( .D(n5739), .SI(d10[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d10[35]) );
  SDFFRXL d10_reg_34_ ( .D(n5738), .SI(d10[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d10[34]) );
  SDFFRXL d10_reg_33_ ( .D(n5737), .SI(d10[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d10[33]) );
  SDFFRXL d10_reg_32_ ( .D(n5736), .SI(d10[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d10[32]) );
  SDFFRXL d10_reg_31_ ( .D(n5735), .SI(d10[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d10[31]) );
  SDFFRXL d10_reg_30_ ( .D(n5734), .SI(d10[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d10[30]) );
  SDFFRXL d10_reg_29_ ( .D(n5733), .SI(d10[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d10[29]) );
  SDFFRXL d10_reg_28_ ( .D(n5732), .SI(d10[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d10[28]) );
  SDFFRXL d10_reg_27_ ( .D(n5731), .SI(d10[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d10[27]) );
  SDFFRXL d10_reg_26_ ( .D(n5730), .SI(d10[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d10[26]) );
  SDFFRXL d10_reg_25_ ( .D(n5729), .SI(d10[24]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d10[25]) );
  SDFFRXL d10_reg_24_ ( .D(n5728), .SI(d10[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d10[24]) );
  SDFFRXL d10_reg_23_ ( .D(n5727), .SI(d10[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d10[23]) );
  SDFFRXL d10_reg_22_ ( .D(n5726), .SI(d10[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d10[22]) );
  SDFFRXL d10_reg_21_ ( .D(n5725), .SI(d10[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d10[21]) );
  SDFFRXL d10_reg_20_ ( .D(n5724), .SI(d10[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d10[20]) );
  SDFFRXL d10_reg_19_ ( .D(n5723), .SI(d10[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d10[19]) );
  SDFFRXL d10_reg_18_ ( .D(n5722), .SI(d10[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d10[18]) );
  SDFFRXL d10_reg_17_ ( .D(n5721), .SI(d10[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d10[17]) );
  SDFFRXL d10_reg_16_ ( .D(n5720), .SI(d10[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d10[16]) );
  SDFFRXL d10_reg_15_ ( .D(n5719), .SI(d10[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d10[15]) );
  SDFFRXL d10_reg_14_ ( .D(n5718), .SI(d10[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d10[14]) );
  SDFFRXL d10_reg_13_ ( .D(n5717), .SI(d10[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d10[13]) );
  SDFFRXL d10_reg_12_ ( .D(n5716), .SI(d10[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d10[12]) );
  SDFFRXL d10_reg_11_ ( .D(n5715), .SI(d10[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d10[11]) );
  SDFFRXL d10_reg_10_ ( .D(n5714), .SI(d10[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d10[10]) );
  SDFFRXL d10_reg_9_ ( .D(n5713), .SI(d10[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d10[9]) );
  SDFFRXL d10_reg_8_ ( .D(n5712), .SI(d10[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d10[8]) );
  SDFFRXL d10_reg_7_ ( .D(n5711), .SI(d10[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d10[7]) );
  SDFFRXL d10_reg_6_ ( .D(n5710), .SI(d10[5]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d10[6]) );
  SDFFRXL d10_reg_5_ ( .D(n5709), .SI(d10[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d10[5]) );
  SDFFRXL d10_reg_4_ ( .D(n5708), .SI(d10[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d10[4]) );
  SDFFRXL d10_reg_3_ ( .D(n5707), .SI(d10[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d10[3]) );
  SDFFRXL d10_reg_2_ ( .D(n5706), .SI(d10[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d10[2]) );
  SDFFRXL d11_reg_35_ ( .D(n5703), .SI(d11[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d11[35]) );
  SDFFRXL d11_reg_34_ ( .D(n5702), .SI(d11[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d11[34]) );
  SDFFRXL d11_reg_33_ ( .D(n5701), .SI(d11[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d11[33]) );
  SDFFRXL d11_reg_32_ ( .D(n5700), .SI(d11[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d11[32]) );
  SDFFRXL d11_reg_31_ ( .D(n5699), .SI(d11[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d11[31]) );
  SDFFRXL d11_reg_30_ ( .D(n5698), .SI(d11[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d11[30]) );
  SDFFRXL d11_reg_29_ ( .D(n5697), .SI(d11[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d11[29]) );
  SDFFRXL d11_reg_28_ ( .D(n5696), .SI(d11[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d11[28]) );
  SDFFRXL d11_reg_27_ ( .D(n5695), .SI(d11[26]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d11[27]) );
  SDFFRXL d11_reg_26_ ( .D(n5694), .SI(d11[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d11[26]) );
  SDFFRXL d11_reg_25_ ( .D(n5693), .SI(d11[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d11[25]) );
  SDFFRXL d11_reg_24_ ( .D(n5692), .SI(d11[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d11[24]) );
  SDFFRXL d11_reg_23_ ( .D(n5691), .SI(d11[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d11[23]) );
  SDFFRXL d11_reg_22_ ( .D(n5690), .SI(d11[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d11[22]) );
  SDFFRXL d11_reg_21_ ( .D(n5689), .SI(d11[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d11[21]) );
  SDFFRXL d11_reg_20_ ( .D(n5688), .SI(d11[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d11[20]) );
  SDFFRXL d11_reg_19_ ( .D(n5687), .SI(d11[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d11[19]) );
  SDFFRXL d11_reg_18_ ( .D(n5686), .SI(d11[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d11[18]) );
  SDFFRXL d11_reg_17_ ( .D(n5685), .SI(d11[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d11[17]) );
  SDFFRXL d11_reg_16_ ( .D(n5684), .SI(d11[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d11[16]) );
  SDFFRXL d11_reg_15_ ( .D(n5683), .SI(d11[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d11[15]) );
  SDFFRXL d11_reg_14_ ( .D(n5682), .SI(d11[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d11[14]) );
  SDFFRXL d11_reg_13_ ( .D(n5681), .SI(d11[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d11[13]) );
  SDFFRXL d11_reg_12_ ( .D(n5680), .SI(d11[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d11[12]) );
  SDFFRXL d11_reg_11_ ( .D(n5679), .SI(d11[10]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d11[11]) );
  SDFFRXL d11_reg_10_ ( .D(n5678), .SI(d11[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d11[10]) );
  SDFFRXL d11_reg_9_ ( .D(n5677), .SI(d11[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d11[9]) );
  SDFFRXL d11_reg_8_ ( .D(n5676), .SI(d11[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d11[8]) );
  SDFFRXL d11_reg_7_ ( .D(n5675), .SI(d11[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d11[7]) );
  SDFFRXL d11_reg_6_ ( .D(n5674), .SI(d11[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d11[6]) );
  SDFFRXL d11_reg_5_ ( .D(n5673), .SI(d11[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d11[5]) );
  SDFFRXL d11_reg_4_ ( .D(n5672), .SI(d11[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d11[4]) );
  SDFFRXL d11_reg_3_ ( .D(n5671), .SI(d11[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d11[3]) );
  SDFFRXL d12_reg_35_ ( .D(n5667), .SI(d12[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d12[35]) );
  SDFFRXL d12_reg_34_ ( .D(n5666), .SI(d12[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d12[34]) );
  SDFFRXL d12_reg_33_ ( .D(n5665), .SI(d12[32]), .SE(test_se), .CK(clk), .RN(
        n8930), .Q(d12[33]) );
  SDFFRXL d12_reg_32_ ( .D(n5664), .SI(d12[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d12[32]) );
  SDFFRXL d12_reg_31_ ( .D(n5663), .SI(d12[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d12[31]) );
  SDFFRXL d12_reg_30_ ( .D(n5662), .SI(d12[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d12[30]) );
  SDFFRXL d12_reg_29_ ( .D(n5661), .SI(d12[28]), .SE(test_se), .CK(clk), .RN(
        n9056), .Q(d12[29]) );
  SDFFRXL d12_reg_28_ ( .D(n5660), .SI(d12[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d12[28]) );
  SDFFRXL d12_reg_27_ ( .D(n5659), .SI(d12[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d12[27]) );
  SDFFRXL d12_reg_26_ ( .D(n5658), .SI(d12[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d12[26]) );
  SDFFRXL d12_reg_25_ ( .D(n5657), .SI(d12[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d12[25]) );
  SDFFRXL d12_reg_24_ ( .D(n5656), .SI(d12[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d12[24]) );
  SDFFRXL d12_reg_23_ ( .D(n5655), .SI(d12[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d12[23]) );
  SDFFRXL d12_reg_22_ ( .D(n5654), .SI(d12[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d12[22]) );
  SDFFRXL d12_reg_21_ ( .D(n5653), .SI(d12[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d12[21]) );
  SDFFRXL d12_reg_20_ ( .D(n5652), .SI(d12[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d12[20]) );
  SDFFRXL d12_reg_19_ ( .D(n5651), .SI(d12[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d12[19]) );
  SDFFRXL d12_reg_18_ ( .D(n5650), .SI(d12[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d12[18]) );
  SDFFRXL d12_reg_17_ ( .D(n5649), .SI(d12[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d12[17]) );
  SDFFRXL d12_reg_16_ ( .D(n5648), .SI(d12[15]), .SE(test_se), .CK(clk), .RN(
        n9088), .Q(d12[16]) );
  SDFFRXL d12_reg_15_ ( .D(n5647), .SI(d12[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d12[15]) );
  SDFFRXL d12_reg_14_ ( .D(n5646), .SI(d12[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d12[14]) );
  SDFFRXL d12_reg_13_ ( .D(n5645), .SI(d12[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d12[13]) );
  SDFFRXL d12_reg_12_ ( .D(n5644), .SI(d12[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d12[12]) );
  SDFFRXL d12_reg_11_ ( .D(n5643), .SI(d12[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d12[11]) );
  SDFFRXL d12_reg_10_ ( .D(n5642), .SI(d12[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d12[10]) );
  SDFFRXL d12_reg_9_ ( .D(n5641), .SI(d12[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d12[9]) );
  SDFFRXL d12_reg_8_ ( .D(n5640), .SI(d12[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d12[8]) );
  SDFFRXL d12_reg_7_ ( .D(n5639), .SI(d12[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d12[7]) );
  SDFFRXL d12_reg_6_ ( .D(n5638), .SI(d12[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d12[6]) );
  SDFFRXL d12_reg_5_ ( .D(n5637), .SI(d12[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d12[5]) );
  SDFFRXL d12_reg_4_ ( .D(n5636), .SI(d12[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d12[4]) );
  SDFFRXL d12_reg_3_ ( .D(n5635), .SI(d12[2]), .SE(test_se), .CK(clk), .RN(
        n9119), .Q(d12[3]) );
  SDFFRXL d12_reg_2_ ( .D(n5634), .SI(d12[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d12[2]) );
  SDFFRXL d13_reg_35_ ( .D(n5631), .SI(d13[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d13[35]) );
  SDFFRXL d13_reg_34_ ( .D(n5630), .SI(d13[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d13[34]) );
  SDFFRXL d13_reg_33_ ( .D(n5629), .SI(d13[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d13[33]) );
  SDFFRXL d13_reg_32_ ( .D(n5628), .SI(d13[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d13[32]) );
  SDFFRXL d13_reg_31_ ( .D(n5627), .SI(d13[30]), .SE(test_se), .CK(clk), .RN(
        n9051), .Q(d13[31]) );
  SDFFRXL d13_reg_30_ ( .D(n5626), .SI(d13[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d13[30]) );
  SDFFRXL d13_reg_29_ ( .D(n5625), .SI(d13[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d13[29]) );
  SDFFRXL d13_reg_28_ ( .D(n5624), .SI(d13[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d13[28]) );
  SDFFRXL d13_reg_27_ ( .D(n5623), .SI(d13[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d13[27]) );
  SDFFRXL d13_reg_26_ ( .D(n5622), .SI(d13[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d13[26]) );
  SDFFRXL d13_reg_25_ ( .D(n5621), .SI(d13[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d13[25]) );
  SDFFRXL d13_reg_24_ ( .D(n5620), .SI(d13[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d13[24]) );
  SDFFRXL d13_reg_23_ ( .D(n5619), .SI(d13[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d13[23]) );
  SDFFRXL d13_reg_22_ ( .D(n5618), .SI(d13[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d13[22]) );
  SDFFRXL d13_reg_21_ ( .D(n5617), .SI(d13[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d13[21]) );
  SDFFRXL d13_reg_20_ ( .D(n5616), .SI(d13[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d13[20]) );
  SDFFRXL d13_reg_19_ ( .D(n5615), .SI(d13[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d13[19]) );
  SDFFRXL d13_reg_18_ ( .D(n5614), .SI(d13[17]), .SE(test_se), .CK(clk), .RN(
        n9083), .Q(d13[18]) );
  SDFFRXL d13_reg_17_ ( .D(n5613), .SI(d13[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d13[17]) );
  SDFFRXL d13_reg_16_ ( .D(n5612), .SI(d13[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d13[16]) );
  SDFFRXL d13_reg_15_ ( .D(n5611), .SI(d13[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d13[15]) );
  SDFFRXL d13_reg_14_ ( .D(n5610), .SI(d13[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d13[14]) );
  SDFFRXL d13_reg_13_ ( .D(n5609), .SI(d13[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d13[13]) );
  SDFFRXL d13_reg_12_ ( .D(n5608), .SI(d13[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d13[12]) );
  SDFFRXL d13_reg_11_ ( .D(n5607), .SI(d13[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d13[11]) );
  SDFFRXL d13_reg_10_ ( .D(n5606), .SI(d13[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d13[10]) );
  SDFFRXL d13_reg_9_ ( .D(n5605), .SI(d13[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d13[9]) );
  SDFFRXL d13_reg_8_ ( .D(n5604), .SI(d13[7]), .SE(test_se), .CK(clk), .RN(
        n9107), .Q(d13[8]) );
  SDFFRXL d13_reg_7_ ( .D(n5603), .SI(d13[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d13[7]) );
  SDFFRXL d13_reg_6_ ( .D(n5602), .SI(d13[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d13[6]) );
  SDFFRXL d13_reg_5_ ( .D(n5601), .SI(d13[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d13[5]) );
  SDFFRXL d13_reg_4_ ( .D(n5600), .SI(d13[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d13[4]) );
  SDFFRXL d13_reg_3_ ( .D(n5599), .SI(d13[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d13[3]) );
  SDFFRXL d14_reg_35_ ( .D(n5595), .SI(d14[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d14[35]) );
  SDFFRXL d14_reg_34_ ( .D(n5594), .SI(d14[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d14[34]) );
  SDFFRXL d14_reg_33_ ( .D(n5593), .SI(d14[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d14[33]) );
  SDFFRXL d14_reg_32_ ( .D(n5592), .SI(d14[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d14[32]) );
  SDFFRXL d14_reg_31_ ( .D(n5591), .SI(d14[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d14[31]) );
  SDFFRXL d14_reg_30_ ( .D(n5590), .SI(d14[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d14[30]) );
  SDFFRXL d14_reg_29_ ( .D(n5589), .SI(d14[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d14[29]) );
  SDFFRXL d14_reg_28_ ( .D(n5588), .SI(d14[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d14[28]) );
  SDFFRXL d14_reg_27_ ( .D(n5587), .SI(d14[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d14[27]) );
  SDFFRXL d14_reg_26_ ( .D(n5586), .SI(d14[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d14[26]) );
  SDFFRXL d14_reg_25_ ( .D(n5585), .SI(d14[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d14[25]) );
  SDFFRXL d14_reg_24_ ( .D(n5584), .SI(d14[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d14[24]) );
  SDFFRXL d14_reg_23_ ( .D(n5583), .SI(d14[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d14[23]) );
  SDFFRXL d14_reg_22_ ( .D(n5582), .SI(d14[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d14[22]) );
  SDFFRXL d14_reg_21_ ( .D(n5581), .SI(d14[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d14[21]) );
  SDFFRXL d14_reg_20_ ( .D(n5580), .SI(d14[19]), .SE(test_se), .CK(clk), .RN(
        n9078), .Q(d14[20]) );
  SDFFRXL d14_reg_19_ ( .D(n5579), .SI(d14[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d14[19]) );
  SDFFRXL d14_reg_18_ ( .D(n5578), .SI(d14[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d14[18]) );
  SDFFRXL d14_reg_17_ ( .D(n5577), .SI(d14[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d14[17]) );
  SDFFRXL d14_reg_16_ ( .D(n5576), .SI(d14[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d14[16]) );
  SDFFRXL d14_reg_15_ ( .D(n5575), .SI(d14[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d14[15]) );
  SDFFRXL d14_reg_14_ ( .D(n5574), .SI(d14[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d14[14]) );
  SDFFRXL d14_reg_13_ ( .D(n5573), .SI(d14[12]), .SE(test_se), .CK(clk), .RN(
        n9095), .Q(d14[13]) );
  SDFFRXL d14_reg_12_ ( .D(n5572), .SI(d14[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d14[12]) );
  SDFFRXL d14_reg_11_ ( .D(n5571), .SI(d14[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d14[11]) );
  SDFFRXL d14_reg_10_ ( .D(n5570), .SI(d14[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d14[10]) );
  SDFFRXL d14_reg_9_ ( .D(n5569), .SI(d14[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d14[9]) );
  SDFFRXL d14_reg_8_ ( .D(n5568), .SI(d14[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d14[8]) );
  SDFFRXL d14_reg_7_ ( .D(n5567), .SI(d14[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d14[7]) );
  SDFFRXL d14_reg_6_ ( .D(n5566), .SI(d14[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d14[6]) );
  SDFFRXL d14_reg_5_ ( .D(n5565), .SI(d14[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d14[5]) );
  SDFFRXL d14_reg_4_ ( .D(n5564), .SI(d14[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d14[4]) );
  SDFFRXL d14_reg_3_ ( .D(n5563), .SI(d14[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d14[3]) );
  SDFFRXL d14_reg_2_ ( .D(n5562), .SI(d14[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d14[2]) );
  SDFFRXL d15_reg_35_ ( .D(n5559), .SI(d15[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d15[35]) );
  SDFFRXL d15_reg_34_ ( .D(n5558), .SI(d15[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d15[34]) );
  SDFFRXL d15_reg_33_ ( .D(n5557), .SI(d15[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d15[33]) );
  SDFFRXL d15_reg_32_ ( .D(n5556), .SI(d15[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d15[32]) );
  SDFFRXL d15_reg_31_ ( .D(n5555), .SI(d15[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d15[31]) );
  SDFFRXL d15_reg_30_ ( .D(n5554), .SI(d15[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d15[30]) );
  SDFFRXL d15_reg_29_ ( .D(n5553), .SI(d15[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d15[29]) );
  SDFFRXL d15_reg_28_ ( .D(n5552), .SI(d15[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d15[28]) );
  SDFFRXL d15_reg_27_ ( .D(n5551), .SI(d15[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d15[27]) );
  SDFFRXL d15_reg_26_ ( .D(n5550), .SI(d15[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d15[26]) );
  SDFFRXL d15_reg_25_ ( .D(n5549), .SI(d15[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d15[25]) );
  SDFFRXL d15_reg_24_ ( .D(n5548), .SI(d15[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d15[24]) );
  SDFFRXL d15_reg_23_ ( .D(n5547), .SI(d15[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d15[23]) );
  SDFFRXL d15_reg_22_ ( .D(n5546), .SI(d15[21]), .SE(test_se), .CK(clk), .RN(
        n9073), .Q(d15[22]) );
  SDFFRXL d15_reg_21_ ( .D(n5545), .SI(d15[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d15[21]) );
  SDFFRXL d15_reg_20_ ( .D(n5544), .SI(d15[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d15[20]) );
  SDFFRXL d15_reg_19_ ( .D(n5543), .SI(d15[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d15[19]) );
  SDFFRXL d15_reg_18_ ( .D(n5542), .SI(d15[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d15[18]) );
  SDFFRXL d15_reg_17_ ( .D(n5541), .SI(d15[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d15[17]) );
  SDFFRXL d15_reg_16_ ( .D(n5540), .SI(d15[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d15[16]) );
  SDFFRXL d15_reg_15_ ( .D(n5539), .SI(d15[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d15[15]) );
  SDFFRXL d15_reg_14_ ( .D(n5538), .SI(d15[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d15[14]) );
  SDFFRXL d15_reg_13_ ( .D(n5537), .SI(d15[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d15[13]) );
  SDFFRXL d15_reg_12_ ( .D(n5536), .SI(d15[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d15[12]) );
  SDFFRXL d15_reg_11_ ( .D(n5535), .SI(d15[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d15[11]) );
  SDFFRXL d15_reg_10_ ( .D(n5534), .SI(d15[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d15[10]) );
  SDFFRXL d15_reg_9_ ( .D(n5533), .SI(d15[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d15[9]) );
  SDFFRXL d15_reg_8_ ( .D(n5532), .SI(d15[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d15[8]) );
  SDFFRXL d15_reg_7_ ( .D(n5531), .SI(d15[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d15[7]) );
  SDFFRXL d15_reg_6_ ( .D(n5530), .SI(d15[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d15[6]) );
  SDFFRXL d15_reg_5_ ( .D(n5529), .SI(d15[4]), .SE(test_se), .CK(clk), .RN(
        n9114), .Q(d15[5]) );
  SDFFRXL d15_reg_4_ ( .D(n5528), .SI(d15[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d15[4]) );
  SDFFRXL d15_reg_3_ ( .D(n5527), .SI(d15[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d15[3]) );
  SDFFRXL d15_reg_2_ ( .D(n5526), .SI(d15[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d15[2]) );
  SDFFRXL d15_reg_1_ ( .D(n5525), .SI(d15[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d15[1]) );
  SDFFRXL d16_reg_35_ ( .D(n5523), .SI(d16[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d16[35]) );
  SDFFRXL d16_reg_34_ ( .D(n5522), .SI(d16[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d16[34]) );
  SDFFRXL d16_reg_33_ ( .D(n5521), .SI(d16[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d16[33]) );
  SDFFRXL d16_reg_32_ ( .D(n5520), .SI(d16[31]), .SE(test_se), .CK(clk), .RN(
        n8932), .Q(d16[32]) );
  SDFFRXL d16_reg_31_ ( .D(n5519), .SI(d16[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d16[31]) );
  SDFFRXL d16_reg_30_ ( .D(n5518), .SI(d16[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d16[30]) );
  SDFFRXL d16_reg_29_ ( .D(n5517), .SI(d16[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d16[29]) );
  SDFFRXL d16_reg_28_ ( .D(n5516), .SI(d16[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d16[28]) );
  SDFFRXL d16_reg_27_ ( .D(n5515), .SI(d16[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d16[27]) );
  SDFFRXL d16_reg_26_ ( .D(n5514), .SI(d16[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d16[26]) );
  SDFFRXL d16_reg_25_ ( .D(n5513), .SI(d16[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d16[25]) );
  SDFFRXL d16_reg_24_ ( .D(n5512), .SI(d16[23]), .SE(test_se), .CK(clk), .RN(
        n9068), .Q(d16[24]) );
  SDFFRXL d16_reg_23_ ( .D(n5511), .SI(d16[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d16[23]) );
  SDFFRXL d16_reg_22_ ( .D(n5510), .SI(d16[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d16[22]) );
  SDFFRXL d16_reg_21_ ( .D(n5509), .SI(d16[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d16[21]) );
  SDFFRXL d16_reg_20_ ( .D(n5508), .SI(d16[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d16[20]) );
  SDFFRXL d16_reg_19_ ( .D(n5507), .SI(d16[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d16[19]) );
  SDFFRXL d16_reg_18_ ( .D(n5506), .SI(d16[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d16[18]) );
  SDFFRXL d16_reg_17_ ( .D(n5505), .SI(d16[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d16[17]) );
  SDFFRXL d16_reg_16_ ( .D(n5504), .SI(d16[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d16[16]) );
  SDFFRXL d16_reg_15_ ( .D(n5503), .SI(d16[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d16[15]) );
  SDFFRXL d16_reg_14_ ( .D(n5502), .SI(d16[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d16[14]) );
  SDFFRXL d16_reg_13_ ( .D(n5501), .SI(d16[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d16[13]) );
  SDFFRXL d16_reg_12_ ( .D(n5500), .SI(d16[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d16[12]) );
  SDFFRXL d16_reg_11_ ( .D(n5499), .SI(d16[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d16[11]) );
  SDFFRXL d16_reg_10_ ( .D(n5498), .SI(d16[9]), .SE(test_se), .CK(clk), .RN(
        n9102), .Q(d16[10]) );
  SDFFRXL d16_reg_9_ ( .D(n5497), .SI(d16[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d16[9]) );
  SDFFRXL d16_reg_8_ ( .D(n5496), .SI(d16[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d16[8]) );
  SDFFRXL d16_reg_7_ ( .D(n5495), .SI(d16[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d16[7]) );
  SDFFRXL d16_reg_6_ ( .D(n5494), .SI(d16[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d16[6]) );
  SDFFRXL d16_reg_5_ ( .D(n5493), .SI(d16[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d16[5]) );
  SDFFRXL d16_reg_4_ ( .D(n5492), .SI(d16[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d16[4]) );
  SDFFRXL d16_reg_3_ ( .D(n5491), .SI(d16[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d16[3]) );
  SDFFRXL d16_reg_2_ ( .D(n5490), .SI(d16[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d16[2]) );
  SDFFRXL d16_reg_1_ ( .D(n5489), .SI(d16[0]), .SE(test_se), .CK(clk), .RN(
        n9123), .Q(d16[1]) );
  SDFFRXL d17_reg_35_ ( .D(n5487), .SI(d17[34]), .SE(test_se), .CK(clk), .RN(
        n8925), .Q(d17[35]) );
  SDFFRXL d17_reg_34_ ( .D(n5486), .SI(d17[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d17[34]) );
  SDFFRXL d17_reg_33_ ( .D(n5485), .SI(d17[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d17[33]) );
  SDFFRXL d17_reg_32_ ( .D(n5484), .SI(d17[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d17[32]) );
  SDFFRXL d17_reg_31_ ( .D(n5483), .SI(d17[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d17[31]) );
  SDFFRXL d17_reg_30_ ( .D(n5482), .SI(d17[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d17[30]) );
  SDFFRXL d17_reg_29_ ( .D(n5481), .SI(d17[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d17[29]) );
  SDFFRXL d17_reg_28_ ( .D(n5480), .SI(d17[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d17[28]) );
  SDFFRXL d17_reg_27_ ( .D(n5479), .SI(d17[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d17[27]) );
  SDFFRXL d17_reg_26_ ( .D(n5478), .SI(d17[25]), .SE(test_se), .CK(clk), .RN(
        n9063), .Q(d17[26]) );
  SDFFRXL d17_reg_25_ ( .D(n5477), .SI(d17[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d17[25]) );
  SDFFRXL d17_reg_24_ ( .D(n5476), .SI(d17[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d17[24]) );
  SDFFRXL d17_reg_23_ ( .D(n5475), .SI(d17[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d17[23]) );
  SDFFRXL d17_reg_22_ ( .D(n5474), .SI(d17[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d17[22]) );
  SDFFRXL d17_reg_21_ ( .D(n5473), .SI(d17[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d17[21]) );
  SDFFRXL d17_reg_20_ ( .D(n5472), .SI(d17[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d17[20]) );
  SDFFRXL d17_reg_19_ ( .D(n5471), .SI(d17[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d17[19]) );
  SDFFRXL d17_reg_18_ ( .D(n5470), .SI(d17[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d17[18]) );
  SDFFRXL d17_reg_17_ ( .D(n5469), .SI(d17[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d17[17]) );
  SDFFRXL d17_reg_16_ ( .D(n5468), .SI(d17[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d17[16]) );
  SDFFRXL d17_reg_15_ ( .D(n5467), .SI(d17[14]), .SE(test_se), .CK(clk), .RN(
        n9090), .Q(d17[15]) );
  SDFFRXL d17_reg_14_ ( .D(n5466), .SI(d17[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d17[14]) );
  SDFFRXL d17_reg_13_ ( .D(n5465), .SI(d17[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d17[13]) );
  SDFFRXL d17_reg_12_ ( .D(n5464), .SI(d17[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d17[12]) );
  SDFFRXL d17_reg_11_ ( .D(n5463), .SI(d17[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d17[11]) );
  SDFFRXL d17_reg_10_ ( .D(n5462), .SI(d17[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d17[10]) );
  SDFFRXL d17_reg_9_ ( .D(n5461), .SI(d17[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d17[9]) );
  SDFFRXL d17_reg_8_ ( .D(n5460), .SI(d17[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d17[8]) );
  SDFFRXL d17_reg_7_ ( .D(n5459), .SI(d17[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d17[7]) );
  SDFFRXL d17_reg_6_ ( .D(n5458), .SI(d17[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d17[6]) );
  SDFFRXL d17_reg_5_ ( .D(n5457), .SI(d17[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d17[5]) );
  SDFFRXL d17_reg_4_ ( .D(n5456), .SI(d17[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d17[4]) );
  SDFFRXL d17_reg_3_ ( .D(n5455), .SI(d17[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d17[3]) );
  SDFFRXL d17_reg_2_ ( .D(n5454), .SI(d17[1]), .SE(test_se), .CK(clk), .RN(
        n9121), .Q(d17[2]) );
  SDFFRXL d18_reg_35_ ( .D(n5451), .SI(d18[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d18[35]) );
  SDFFRXL d18_reg_34_ ( .D(n5450), .SI(d18[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d18[34]) );
  SDFFRXL d18_reg_33_ ( .D(n5449), .SI(d18[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d18[33]) );
  SDFFRXL d18_reg_32_ ( .D(n5448), .SI(d18[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d18[32]) );
  SDFFRXL d18_reg_31_ ( .D(n5447), .SI(d18[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d18[31]) );
  SDFFRXL d18_reg_30_ ( .D(n5446), .SI(d18[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d18[30]) );
  SDFFRXL d18_reg_29_ ( .D(n5445), .SI(d18[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d18[29]) );
  SDFFRXL d18_reg_28_ ( .D(n5444), .SI(d18[27]), .SE(test_se), .CK(clk), .RN(
        n9058), .Q(d18[28]) );
  SDFFRXL d18_reg_27_ ( .D(n5443), .SI(d18[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d18[27]) );
  SDFFRXL d18_reg_26_ ( .D(n5442), .SI(d18[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d18[26]) );
  SDFFRXL d18_reg_25_ ( .D(n5441), .SI(d18[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d18[25]) );
  SDFFRXL d18_reg_24_ ( .D(n5440), .SI(d18[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d18[24]) );
  SDFFRXL d18_reg_23_ ( .D(n5439), .SI(d18[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d18[23]) );
  SDFFRXL d18_reg_22_ ( .D(n5438), .SI(d18[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d18[22]) );
  SDFFRXL d18_reg_21_ ( .D(n5437), .SI(d18[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d18[21]) );
  SDFFRXL d18_reg_20_ ( .D(n5436), .SI(d18[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d18[20]) );
  SDFFRXL d18_reg_19_ ( .D(n5435), .SI(d18[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d18[19]) );
  SDFFRXL d18_reg_18_ ( .D(n5434), .SI(d18[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d18[18]) );
  SDFFRXL d18_reg_17_ ( .D(n5433), .SI(d18[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d18[17]) );
  SDFFRXL d18_reg_16_ ( .D(n5432), .SI(d18[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d18[16]) );
  SDFFRXL d18_reg_15_ ( .D(n5431), .SI(d18[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d18[15]) );
  SDFFRXL d18_reg_14_ ( .D(n5430), .SI(d18[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d18[14]) );
  SDFFRXL d18_reg_13_ ( .D(n5429), .SI(d18[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d18[13]) );
  SDFFRXL d18_reg_12_ ( .D(n5428), .SI(d18[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d18[12]) );
  SDFFRXL d18_reg_11_ ( .D(n5427), .SI(d18[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d18[11]) );
  SDFFRXL d18_reg_10_ ( .D(n5426), .SI(d18[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d18[10]) );
  SDFFRXL d18_reg_9_ ( .D(n5425), .SI(d18[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d18[9]) );
  SDFFRXL d18_reg_8_ ( .D(n5424), .SI(d18[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d18[8]) );
  SDFFRXL d18_reg_7_ ( .D(n5423), .SI(d18[6]), .SE(test_se), .CK(clk), .RN(
        n9109), .Q(d18[7]) );
  SDFFRXL d18_reg_6_ ( .D(n5422), .SI(d18[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d18[6]) );
  SDFFRXL d18_reg_5_ ( .D(n5421), .SI(d18[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d18[5]) );
  SDFFRXL d18_reg_4_ ( .D(n5420), .SI(d18[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d18[4]) );
  SDFFRXL d18_reg_3_ ( .D(n5419), .SI(d18[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d18[3]) );
  SDFFRXL d19_reg_35_ ( .D(n5415), .SI(d19[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d19[35]) );
  SDFFRXL d19_reg_34_ ( .D(n5414), .SI(d19[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d19[34]) );
  SDFFRXL d19_reg_33_ ( .D(n5413), .SI(d19[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d19[33]) );
  SDFFRXL d19_reg_32_ ( .D(n5412), .SI(d19[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d19[32]) );
  SDFFRXL d19_reg_31_ ( .D(n5411), .SI(d19[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d19[31]) );
  SDFFRXL d19_reg_30_ ( .D(n5410), .SI(d19[29]), .SE(test_se), .CK(clk), .RN(
        n9053), .Q(d19[30]) );
  SDFFRXL d19_reg_29_ ( .D(n5409), .SI(d19[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d19[29]) );
  SDFFRXL d19_reg_28_ ( .D(n5408), .SI(d19[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d19[28]) );
  SDFFRXL d19_reg_27_ ( .D(n5407), .SI(d19[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d19[27]) );
  SDFFRXL d19_reg_26_ ( .D(n5406), .SI(d19[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d19[26]) );
  SDFFRXL d19_reg_25_ ( .D(n5405), .SI(d19[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d19[25]) );
  SDFFRXL d19_reg_24_ ( .D(n5404), .SI(d19[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d19[24]) );
  SDFFRXL d19_reg_23_ ( .D(n5403), .SI(d19[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d19[23]) );
  SDFFRXL d19_reg_22_ ( .D(n5402), .SI(d19[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d19[22]) );
  SDFFRXL d19_reg_21_ ( .D(n5401), .SI(d19[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d19[21]) );
  SDFFRXL d19_reg_20_ ( .D(n5400), .SI(d19[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d19[20]) );
  SDFFRXL d19_reg_19_ ( .D(n5399), .SI(d19[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d19[19]) );
  SDFFRXL d19_reg_18_ ( .D(n5398), .SI(d19[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d19[18]) );
  SDFFRXL d19_reg_17_ ( .D(n5397), .SI(d19[16]), .SE(test_se), .CK(clk), .RN(
        n9085), .Q(d19[17]) );
  SDFFRXL d19_reg_16_ ( .D(n5396), .SI(d19[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d19[16]) );
  SDFFRXL d19_reg_15_ ( .D(n5395), .SI(d19[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d19[15]) );
  SDFFRXL d19_reg_14_ ( .D(n5394), .SI(d19[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d19[14]) );
  SDFFRXL d19_reg_13_ ( .D(n5393), .SI(d19[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d19[13]) );
  SDFFRXL d19_reg_12_ ( .D(n5392), .SI(d19[11]), .SE(test_se), .CK(clk), .RN(
        n9097), .Q(d19[12]) );
  SDFFRXL d19_reg_11_ ( .D(n5391), .SI(d19[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d19[11]) );
  SDFFRXL d19_reg_10_ ( .D(n5390), .SI(d19[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d19[10]) );
  SDFFRXL d19_reg_9_ ( .D(n5389), .SI(d19[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d19[9]) );
  SDFFRXL d19_reg_8_ ( .D(n5388), .SI(d19[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d19[8]) );
  SDFFRXL d19_reg_7_ ( .D(n5387), .SI(d19[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d19[7]) );
  SDFFRXL d19_reg_6_ ( .D(n5386), .SI(d19[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d19[6]) );
  SDFFRXL d19_reg_5_ ( .D(n5385), .SI(d19[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d19[5]) );
  SDFFRXL d19_reg_4_ ( .D(n5384), .SI(d19[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d19[4]) );
  SDFFRXL d19_reg_3_ ( .D(n5383), .SI(d19[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d19[3]) );
  SDFFRXL d19_reg_2_ ( .D(n5382), .SI(d19[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d19[2]) );
  SDFFRXL d20_reg_35_ ( .D(n5379), .SI(d20[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d20[35]) );
  SDFFRXL d20_reg_34_ ( .D(n5378), .SI(d20[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d20[34]) );
  SDFFRXL d20_reg_33_ ( .D(n5377), .SI(d20[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d20[33]) );
  SDFFRXL d20_reg_32_ ( .D(n5376), .SI(d20[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d20[32]) );
  SDFFRXL d20_reg_31_ ( .D(n5375), .SI(d20[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d20[31]) );
  SDFFRXL d20_reg_30_ ( .D(n5374), .SI(d20[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d20[30]) );
  SDFFRXL d20_reg_29_ ( .D(n5373), .SI(d20[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d20[29]) );
  SDFFRXL d20_reg_28_ ( .D(n5372), .SI(d20[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d20[28]) );
  SDFFRXL d20_reg_27_ ( .D(n5371), .SI(d20[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d20[27]) );
  SDFFRXL d20_reg_26_ ( .D(n5370), .SI(d20[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d20[26]) );
  SDFFRXL d20_reg_25_ ( .D(n5369), .SI(d20[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d20[25]) );
  SDFFRXL d20_reg_24_ ( .D(n5368), .SI(d20[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d20[24]) );
  SDFFRXL d20_reg_23_ ( .D(n5367), .SI(d20[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d20[23]) );
  SDFFRXL d20_reg_22_ ( .D(n5366), .SI(d20[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d20[22]) );
  SDFFRXL d20_reg_21_ ( .D(n5365), .SI(d20[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d20[21]) );
  SDFFRXL d20_reg_20_ ( .D(n5364), .SI(d20[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d20[20]) );
  SDFFRXL d20_reg_19_ ( .D(n5363), .SI(d20[18]), .SE(test_se), .CK(clk), .RN(
        n9080), .Q(d20[19]) );
  SDFFRXL d20_reg_18_ ( .D(n5362), .SI(d20[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d20[18]) );
  SDFFRXL d20_reg_17_ ( .D(n5361), .SI(d20[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d20[17]) );
  SDFFRXL d20_reg_16_ ( .D(n5360), .SI(d20[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d20[16]) );
  SDFFRXL d20_reg_15_ ( .D(n5359), .SI(d20[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d20[15]) );
  SDFFRXL d20_reg_14_ ( .D(n5358), .SI(d20[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d20[14]) );
  SDFFRXL d20_reg_13_ ( .D(n5357), .SI(d20[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d20[13]) );
  SDFFRXL d20_reg_12_ ( .D(n5356), .SI(d20[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d20[12]) );
  SDFFRXL d20_reg_11_ ( .D(n5355), .SI(d20[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d20[11]) );
  SDFFRXL d20_reg_10_ ( .D(n5354), .SI(d20[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d20[10]) );
  SDFFRXL d20_reg_9_ ( .D(n5353), .SI(d20[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d20[9]) );
  SDFFRXL d20_reg_8_ ( .D(n5352), .SI(d20[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d20[8]) );
  SDFFRXL d20_reg_7_ ( .D(n5351), .SI(d20[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d20[7]) );
  SDFFRXL d20_reg_6_ ( .D(n5350), .SI(d20[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d20[6]) );
  SDFFRXL d20_reg_5_ ( .D(n5349), .SI(d20[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d20[5]) );
  SDFFRXL d20_reg_4_ ( .D(n5348), .SI(d20[3]), .SE(test_se), .CK(clk), .RN(
        n9116), .Q(d20[4]) );
  SDFFRXL d20_reg_3_ ( .D(n5347), .SI(d20[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d20[3]) );
  SDFFRXL d21_reg_35_ ( .D(n5343), .SI(d21[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d21[35]) );
  SDFFRXL d21_reg_34_ ( .D(n5342), .SI(d21[33]), .SE(test_se), .CK(clk), .RN(
        n8927), .Q(d21[34]) );
  SDFFRXL d21_reg_33_ ( .D(n5341), .SI(d21[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d21[33]) );
  SDFFRXL d21_reg_32_ ( .D(n5340), .SI(d21[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d21[32]) );
  SDFFRXL d21_reg_31_ ( .D(n5339), .SI(d21[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d21[31]) );
  SDFFRXL d21_reg_30_ ( .D(n5338), .SI(d21[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d21[30]) );
  SDFFRXL d21_reg_29_ ( .D(n5337), .SI(d21[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d21[29]) );
  SDFFRXL d21_reg_28_ ( .D(n5336), .SI(d21[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d21[28]) );
  SDFFRXL d21_reg_27_ ( .D(n5335), .SI(d21[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d21[27]) );
  SDFFRXL d21_reg_26_ ( .D(n5334), .SI(d21[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d21[26]) );
  SDFFRXL d21_reg_25_ ( .D(n5333), .SI(d21[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d21[25]) );
  SDFFRXL d21_reg_24_ ( .D(n5332), .SI(d21[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d21[24]) );
  SDFFRXL d21_reg_23_ ( .D(n5331), .SI(d21[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d21[23]) );
  SDFFRXL d21_reg_22_ ( .D(n5330), .SI(d21[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d21[22]) );
  SDFFRXL d21_reg_21_ ( .D(n5329), .SI(d21[20]), .SE(test_se), .CK(clk), .RN(
        n9075), .Q(d21[21]) );
  SDFFRXL d21_reg_20_ ( .D(n5328), .SI(d21[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d21[20]) );
  SDFFRXL d21_reg_19_ ( .D(n5327), .SI(d21[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d21[19]) );
  SDFFRXL d21_reg_18_ ( .D(n5326), .SI(d21[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d21[18]) );
  SDFFRXL d21_reg_17_ ( .D(n5325), .SI(d21[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d21[17]) );
  SDFFRXL d21_reg_16_ ( .D(n5324), .SI(d21[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d21[16]) );
  SDFFRXL d21_reg_15_ ( .D(n5323), .SI(d21[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d21[15]) );
  SDFFRXL d21_reg_14_ ( .D(n5322), .SI(d21[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d21[14]) );
  SDFFRXL d21_reg_13_ ( .D(n5321), .SI(d21[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d21[13]) );
  SDFFRXL d21_reg_12_ ( .D(n5320), .SI(d21[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d21[12]) );
  SDFFRXL d21_reg_11_ ( .D(n5319), .SI(d21[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d21[11]) );
  SDFFRXL d21_reg_10_ ( .D(n5318), .SI(d21[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d21[10]) );
  SDFFRXL d21_reg_9_ ( .D(n5317), .SI(d21[8]), .SE(test_se), .CK(clk), .RN(
        n9104), .Q(d21[9]) );
  SDFFRXL d21_reg_8_ ( .D(n5316), .SI(d21[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d21[8]) );
  SDFFRXL d21_reg_7_ ( .D(n5315), .SI(d21[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d21[7]) );
  SDFFRXL d21_reg_6_ ( .D(n5314), .SI(d21[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d21[6]) );
  SDFFRXL d21_reg_5_ ( .D(n5313), .SI(d21[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d21[5]) );
  SDFFRXL d21_reg_4_ ( .D(n5312), .SI(d21[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d21[4]) );
  SDFFRXL d21_reg_3_ ( .D(n5311), .SI(d21[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d21[3]) );
  SDFFRXL d21_reg_2_ ( .D(n5310), .SI(d21[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d21[2]) );
  SDFFRXL d22_reg_35_ ( .D(n5307), .SI(d22[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d22[35]) );
  SDFFRXL d22_reg_34_ ( .D(n5306), .SI(d22[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d22[34]) );
  SDFFRXL d22_reg_33_ ( .D(n5305), .SI(d22[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d22[33]) );
  SDFFRXL d22_reg_32_ ( .D(n5304), .SI(d22[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d22[32]) );
  SDFFRXL d22_reg_31_ ( .D(n5303), .SI(d22[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d22[31]) );
  SDFFRXL d22_reg_30_ ( .D(n5302), .SI(d22[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d22[30]) );
  SDFFRXL d22_reg_29_ ( .D(n5301), .SI(d22[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d22[29]) );
  SDFFRXL d22_reg_28_ ( .D(n5300), .SI(d22[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d22[28]) );
  SDFFRXL d22_reg_27_ ( .D(n5299), .SI(d22[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d22[27]) );
  SDFFRXL d22_reg_26_ ( .D(n5298), .SI(d22[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d22[26]) );
  SDFFRXL d22_reg_25_ ( .D(n5297), .SI(d22[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d22[25]) );
  SDFFRXL d22_reg_24_ ( .D(n5296), .SI(d22[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d22[24]) );
  SDFFRXL d22_reg_23_ ( .D(n5295), .SI(d22[22]), .SE(test_se), .CK(clk), .RN(
        n9070), .Q(d22[23]) );
  SDFFRXL d22_reg_22_ ( .D(n5294), .SI(d22[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d22[22]) );
  SDFFRXL d22_reg_21_ ( .D(n5293), .SI(d22[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d22[21]) );
  SDFFRXL d22_reg_20_ ( .D(n5292), .SI(d22[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d22[20]) );
  SDFFRXL d22_reg_19_ ( .D(n5291), .SI(d22[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d22[19]) );
  SDFFRXL d22_reg_18_ ( .D(n5290), .SI(d22[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d22[18]) );
  SDFFRXL d22_reg_17_ ( .D(n5289), .SI(d22[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d22[17]) );
  SDFFRXL d22_reg_16_ ( .D(n5288), .SI(d22[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d22[16]) );
  SDFFRXL d22_reg_15_ ( .D(n5287), .SI(d22[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d22[15]) );
  SDFFRXL d22_reg_14_ ( .D(n5286), .SI(d22[13]), .SE(test_se), .CK(clk), .RN(
        n9092), .Q(d22[14]) );
  SDFFRXL d22_reg_13_ ( .D(n5285), .SI(d22[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d22[13]) );
  SDFFRXL d22_reg_12_ ( .D(n5284), .SI(d22[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d22[12]) );
  SDFFRXL d22_reg_11_ ( .D(n5283), .SI(d22[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d22[11]) );
  SDFFRXL d22_reg_10_ ( .D(n5282), .SI(d22[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d22[10]) );
  SDFFRXL d22_reg_9_ ( .D(n5281), .SI(d22[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d22[9]) );
  SDFFRXL d22_reg_8_ ( .D(n5280), .SI(d22[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d22[8]) );
  SDFFRXL d22_reg_7_ ( .D(n5279), .SI(d22[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d22[7]) );
  SDFFRXL d22_reg_6_ ( .D(n5278), .SI(d22[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d22[6]) );
  SDFFRXL d22_reg_5_ ( .D(n5277), .SI(d22[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d22[5]) );
  SDFFRXL d22_reg_4_ ( .D(n5276), .SI(d22[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d22[4]) );
  SDFFRXL d22_reg_3_ ( .D(n5275), .SI(d22[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d22[3]) );
  SDFFRXL d22_reg_2_ ( .D(n5274), .SI(d22[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d22[2]) );
  SDFFRXL d23_reg_35_ ( .D(n5271), .SI(d23[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d23[35]) );
  SDFFRXL d23_reg_34_ ( .D(n5270), .SI(d23[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d23[34]) );
  SDFFRXL d23_reg_33_ ( .D(n5269), .SI(d23[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d23[33]) );
  SDFFRXL d23_reg_32_ ( .D(n5268), .SI(d23[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d23[32]) );
  SDFFRXL d23_reg_31_ ( .D(n5267), .SI(d23[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d23[31]) );
  SDFFRXL d23_reg_30_ ( .D(n5266), .SI(d23[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d23[30]) );
  SDFFRXL d23_reg_29_ ( .D(n5265), .SI(d23[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d23[29]) );
  SDFFRXL d23_reg_28_ ( .D(n5264), .SI(d23[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d23[28]) );
  SDFFRXL d23_reg_27_ ( .D(n5263), .SI(d23[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d23[27]) );
  SDFFRXL d23_reg_26_ ( .D(n5262), .SI(d23[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d23[26]) );
  SDFFRXL d23_reg_25_ ( .D(n5261), .SI(d23[24]), .SE(test_se), .CK(clk), .RN(
        n9065), .Q(d23[25]) );
  SDFFRXL d23_reg_24_ ( .D(n5260), .SI(d23[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d23[24]) );
  SDFFRXL d23_reg_23_ ( .D(n5259), .SI(d23[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d23[23]) );
  SDFFRXL d23_reg_22_ ( .D(n5258), .SI(d23[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d23[22]) );
  SDFFRXL d23_reg_21_ ( .D(n5257), .SI(d23[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d23[21]) );
  SDFFRXL d23_reg_20_ ( .D(n5256), .SI(d23[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d23[20]) );
  SDFFRXL d23_reg_19_ ( .D(n5255), .SI(d23[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d23[19]) );
  SDFFRXL d23_reg_18_ ( .D(n5254), .SI(d23[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d23[18]) );
  SDFFRXL d23_reg_17_ ( .D(n5253), .SI(d23[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d23[17]) );
  SDFFRXL d23_reg_16_ ( .D(n5252), .SI(d23[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d23[16]) );
  SDFFRXL d23_reg_15_ ( .D(n5251), .SI(d23[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d23[15]) );
  SDFFRXL d23_reg_14_ ( .D(n5250), .SI(d23[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d23[14]) );
  SDFFRXL d23_reg_13_ ( .D(n5249), .SI(d23[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d23[13]) );
  SDFFRXL d23_reg_12_ ( .D(n5248), .SI(d23[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d23[12]) );
  SDFFRXL d23_reg_11_ ( .D(n5247), .SI(d23[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d23[11]) );
  SDFFRXL d23_reg_10_ ( .D(n5246), .SI(d23[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d23[10]) );
  SDFFRXL d23_reg_9_ ( .D(n5245), .SI(d23[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d23[9]) );
  SDFFRXL d23_reg_8_ ( .D(n5244), .SI(d23[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d23[8]) );
  SDFFRXL d23_reg_7_ ( .D(n5243), .SI(d23[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d23[7]) );
  SDFFRXL d23_reg_6_ ( .D(n5242), .SI(d23[5]), .SE(test_se), .CK(clk), .RN(
        n9111), .Q(d23[6]) );
  SDFFRXL d23_reg_5_ ( .D(n5241), .SI(d23[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d23[5]) );
  SDFFRXL d23_reg_4_ ( .D(n5240), .SI(d23[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d23[4]) );
  SDFFRXL d23_reg_3_ ( .D(n5239), .SI(d23[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d23[3]) );
  SDFFRXL d23_reg_2_ ( .D(n5238), .SI(d23[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d23[2]) );
  SDFFRXL d23_reg_1_ ( .D(n5237), .SI(d23[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d23[1]) );
  SDFFRXL d24_reg_35_ ( .D(n5235), .SI(d24[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d24[35]) );
  SDFFRXL d24_reg_34_ ( .D(n5234), .SI(d24[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d24[34]) );
  SDFFRXL d24_reg_33_ ( .D(n5233), .SI(d24[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d24[33]) );
  SDFFRXL d24_reg_32_ ( .D(n5232), .SI(d24[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d24[32]) );
  SDFFRXL d24_reg_31_ ( .D(n5231), .SI(d24[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d24[31]) );
  SDFFRXL d24_reg_30_ ( .D(n5230), .SI(d24[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d24[30]) );
  SDFFRXL d24_reg_29_ ( .D(n5229), .SI(d24[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d24[29]) );
  SDFFRXL d24_reg_28_ ( .D(n5228), .SI(d24[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d24[28]) );
  SDFFRXL d24_reg_27_ ( .D(n5227), .SI(d24[26]), .SE(test_se), .CK(clk), .RN(
        n9060), .Q(d24[27]) );
  SDFFRXL d24_reg_26_ ( .D(n5226), .SI(d24[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d24[26]) );
  SDFFRXL d24_reg_25_ ( .D(n5225), .SI(d24[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d24[25]) );
  SDFFRXL d24_reg_24_ ( .D(n5224), .SI(d24[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d24[24]) );
  SDFFRXL d24_reg_23_ ( .D(n5223), .SI(d24[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d24[23]) );
  SDFFRXL d24_reg_22_ ( .D(n5222), .SI(d24[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d24[22]) );
  SDFFRXL d24_reg_21_ ( .D(n5221), .SI(d24[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d24[21]) );
  SDFFRXL d24_reg_20_ ( .D(n5220), .SI(d24[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d24[20]) );
  SDFFRXL d24_reg_19_ ( .D(n5219), .SI(d24[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d24[19]) );
  SDFFRXL d24_reg_18_ ( .D(n5218), .SI(d24[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d24[18]) );
  SDFFRXL d24_reg_17_ ( .D(n5217), .SI(d24[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d24[17]) );
  SDFFRXL d24_reg_16_ ( .D(n5216), .SI(d24[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d24[16]) );
  SDFFRXL d24_reg_15_ ( .D(n5215), .SI(d24[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d24[15]) );
  SDFFRXL d24_reg_14_ ( .D(n5214), .SI(d24[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d24[14]) );
  SDFFRXL d24_reg_13_ ( .D(n5213), .SI(d24[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d24[13]) );
  SDFFRXL d24_reg_12_ ( .D(n5212), .SI(d24[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d24[12]) );
  SDFFRXL d24_reg_11_ ( .D(n5211), .SI(d24[10]), .SE(test_se), .CK(clk), .RN(
        n9099), .Q(d24[11]) );
  SDFFRXL d24_reg_10_ ( .D(n5210), .SI(d24[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d24[10]) );
  SDFFRXL d24_reg_9_ ( .D(n5209), .SI(d24[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d24[9]) );
  SDFFRXL d24_reg_8_ ( .D(n5208), .SI(d24[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d24[8]) );
  SDFFRXL d24_reg_7_ ( .D(n5207), .SI(d24[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d24[7]) );
  SDFFRXL d24_reg_6_ ( .D(n5206), .SI(d24[5]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d24[6]) );
  SDFFRXL d24_reg_5_ ( .D(n5205), .SI(d24[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d24[5]) );
  SDFFRXL d24_reg_4_ ( .D(n5204), .SI(d24[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d24[4]) );
  SDFFRXL d24_reg_3_ ( .D(n5203), .SI(d24[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d24[3]) );
  SDFFRXL d25_reg_35_ ( .D(n5199), .SI(d25[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d25[35]) );
  SDFFRXL d25_reg_34_ ( .D(n5198), .SI(d25[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d25[34]) );
  SDFFRXL d25_reg_33_ ( .D(n5197), .SI(d25[32]), .SE(test_se), .CK(clk), .RN(
        n8929), .Q(d25[33]) );
  SDFFRXL d25_reg_32_ ( .D(n5196), .SI(d25[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d25[32]) );
  SDFFRXL d25_reg_31_ ( .D(n5195), .SI(d25[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d25[31]) );
  SDFFRXL d25_reg_30_ ( .D(n5194), .SI(d25[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d25[30]) );
  SDFFRXL d25_reg_29_ ( .D(n5193), .SI(d25[28]), .SE(test_se), .CK(clk), .RN(
        n9055), .Q(d25[29]) );
  SDFFRXL d25_reg_28_ ( .D(n5192), .SI(d25[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d25[28]) );
  SDFFRXL d25_reg_27_ ( .D(n5191), .SI(d25[26]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d25[27]) );
  SDFFRXL d25_reg_26_ ( .D(n5190), .SI(d25[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d25[26]) );
  SDFFRXL d25_reg_25_ ( .D(n5189), .SI(d25[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d25[25]) );
  SDFFRXL d25_reg_24_ ( .D(n5188), .SI(d25[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d25[24]) );
  SDFFRXL d25_reg_23_ ( .D(n5187), .SI(d25[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d25[23]) );
  SDFFRXL d25_reg_22_ ( .D(n5186), .SI(d25[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d25[22]) );
  SDFFRXL d25_reg_21_ ( .D(n5185), .SI(d25[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d25[21]) );
  SDFFRXL d25_reg_20_ ( .D(n5184), .SI(d25[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d25[20]) );
  SDFFRXL d25_reg_19_ ( .D(n5183), .SI(d25[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d25[19]) );
  SDFFRXL d25_reg_18_ ( .D(n5182), .SI(d25[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d25[18]) );
  SDFFRXL d25_reg_17_ ( .D(n5181), .SI(d25[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d25[17]) );
  SDFFRXL d25_reg_16_ ( .D(n5180), .SI(d25[15]), .SE(test_se), .CK(clk), .RN(
        n9087), .Q(d25[16]) );
  SDFFRXL d25_reg_15_ ( .D(n5179), .SI(d25[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d25[15]) );
  SDFFRXL d25_reg_14_ ( .D(n5178), .SI(d25[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d25[14]) );
  SDFFRXL d25_reg_13_ ( .D(n5177), .SI(d25[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d25[13]) );
  SDFFRXL d25_reg_12_ ( .D(n5176), .SI(d25[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d25[12]) );
  SDFFRXL d25_reg_11_ ( .D(n5175), .SI(d25[10]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d25[11]) );
  SDFFRXL d25_reg_10_ ( .D(n5174), .SI(d25[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d25[10]) );
  SDFFRXL d25_reg_9_ ( .D(n5173), .SI(d25[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d25[9]) );
  SDFFRXL d25_reg_8_ ( .D(n5172), .SI(d25[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d25[8]) );
  SDFFRXL d25_reg_7_ ( .D(n5171), .SI(d25[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d25[7]) );
  SDFFRXL d25_reg_6_ ( .D(n5170), .SI(d25[5]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d25[6]) );
  SDFFRXL d25_reg_5_ ( .D(n5169), .SI(d25[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d25[5]) );
  SDFFRXL d25_reg_4_ ( .D(n5168), .SI(d25[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d25[4]) );
  SDFFRXL d25_reg_3_ ( .D(n5167), .SI(d25[2]), .SE(test_se), .CK(clk), .RN(
        n9118), .Q(d25[3]) );
  SDFFRXL d25_reg_2_ ( .D(n5166), .SI(d25[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d25[2]) );
  SDFFRXL d26_reg_35_ ( .D(n5163), .SI(d26[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d26[35]) );
  SDFFRXL d26_reg_34_ ( .D(n5162), .SI(d26[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d26[34]) );
  SDFFRXL d26_reg_33_ ( .D(n5161), .SI(d26[32]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d26[33]) );
  SDFFRXL d26_reg_32_ ( .D(n5160), .SI(d26[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d26[32]) );
  SDFFRXL d26_reg_31_ ( .D(n5159), .SI(d26[30]), .SE(test_se), .CK(clk), .RN(
        n9050), .Q(d26[31]) );
  SDFFRXL d26_reg_30_ ( .D(n5158), .SI(d26[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d26[30]) );
  SDFFRXL d26_reg_29_ ( .D(n5157), .SI(d26[28]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d26[29]) );
  SDFFRXL d26_reg_28_ ( .D(n5156), .SI(d26[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d26[28]) );
  SDFFRXL d26_reg_27_ ( .D(n5155), .SI(d26[26]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d26[27]) );
  SDFFRXL d26_reg_26_ ( .D(n5154), .SI(d26[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d26[26]) );
  SDFFRXL d26_reg_25_ ( .D(n5153), .SI(d26[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d26[25]) );
  SDFFRXL d26_reg_24_ ( .D(n5152), .SI(d26[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d26[24]) );
  SDFFRXL d26_reg_23_ ( .D(n5151), .SI(d26[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d26[23]) );
  SDFFRXL d26_reg_22_ ( .D(n5150), .SI(d26[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d26[22]) );
  SDFFRXL d26_reg_21_ ( .D(n5149), .SI(d26[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d26[21]) );
  SDFFRXL d26_reg_20_ ( .D(n5148), .SI(d26[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d26[20]) );
  SDFFRXL d26_reg_19_ ( .D(n5147), .SI(d26[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d26[19]) );
  SDFFRXL d26_reg_18_ ( .D(n5146), .SI(d26[17]), .SE(test_se), .CK(clk), .RN(
        n9082), .Q(d26[18]) );
  SDFFRXL d26_reg_17_ ( .D(n5145), .SI(d26[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d26[17]) );
  SDFFRXL d26_reg_16_ ( .D(n5144), .SI(d26[15]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d26[16]) );
  SDFFRXL d26_reg_15_ ( .D(n5143), .SI(d26[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d26[15]) );
  SDFFRXL d26_reg_14_ ( .D(n5142), .SI(d26[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d26[14]) );
  SDFFRXL d26_reg_13_ ( .D(n5141), .SI(d26[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d26[13]) );
  SDFFRXL d26_reg_12_ ( .D(n5140), .SI(d26[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d26[12]) );
  SDFFRXL d26_reg_11_ ( .D(n5139), .SI(d26[10]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d26[11]) );
  SDFFRXL d26_reg_10_ ( .D(n5138), .SI(d26[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d26[10]) );
  SDFFRXL d26_reg_9_ ( .D(n5137), .SI(d26[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d26[9]) );
  SDFFRXL d26_reg_8_ ( .D(n5136), .SI(d26[7]), .SE(test_se), .CK(clk), .RN(
        n9106), .Q(d26[8]) );
  SDFFRXL d26_reg_7_ ( .D(n5135), .SI(d26[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d26[7]) );
  SDFFRXL d26_reg_6_ ( .D(n5134), .SI(d26[5]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d26[6]) );
  SDFFRXL d26_reg_5_ ( .D(n5133), .SI(d26[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d26[5]) );
  SDFFRXL d26_reg_4_ ( .D(n5132), .SI(d26[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d26[4]) );
  SDFFRXL d26_reg_3_ ( .D(n5131), .SI(d26[2]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d26[3]) );
  SDFFRXL d26_reg_2_ ( .D(n5130), .SI(d26[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d26[2]) );
  SDFFRXL d27_reg_35_ ( .D(n5127), .SI(d27[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d27[35]) );
  SDFFRXL d27_reg_34_ ( .D(n5126), .SI(d27[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d27[34]) );
  SDFFRXL d27_reg_33_ ( .D(n5125), .SI(d27[32]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d27[33]) );
  SDFFRXL d27_reg_32_ ( .D(n5124), .SI(d27[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d27[32]) );
  SDFFRXL d27_reg_31_ ( .D(n5123), .SI(d27[30]), .SE(test_se), .CK(clk), .RN(
        n9049), .Q(d27[31]) );
  SDFFRXL d27_reg_30_ ( .D(n5122), .SI(d27[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d27[30]) );
  SDFFRXL d27_reg_29_ ( .D(n5121), .SI(d27[28]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d27[29]) );
  SDFFRXL d27_reg_28_ ( .D(n5120), .SI(d27[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d27[28]) );
  SDFFRXL d27_reg_27_ ( .D(n5119), .SI(d27[26]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d27[27]) );
  SDFFRXL d27_reg_26_ ( .D(n5118), .SI(d27[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d27[26]) );
  SDFFRXL d27_reg_25_ ( .D(n5117), .SI(d27[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d27[25]) );
  SDFFRXL d27_reg_24_ ( .D(n5116), .SI(d27[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d27[24]) );
  SDFFRXL d27_reg_23_ ( .D(n5115), .SI(d27[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d27[23]) );
  SDFFRXL d27_reg_22_ ( .D(n5114), .SI(d27[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d27[22]) );
  SDFFRXL d27_reg_21_ ( .D(n5113), .SI(d27[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d27[21]) );
  SDFFRXL d27_reg_20_ ( .D(n5112), .SI(d27[19]), .SE(test_se), .CK(clk), .RN(
        n9077), .Q(d27[20]) );
  SDFFRXL d27_reg_19_ ( .D(n5111), .SI(d27[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d27[19]) );
  SDFFRXL d27_reg_18_ ( .D(n5110), .SI(d27[17]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d27[18]) );
  SDFFRXL d27_reg_17_ ( .D(n5109), .SI(d27[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d27[17]) );
  SDFFRXL d27_reg_16_ ( .D(n5108), .SI(d27[15]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d27[16]) );
  SDFFRXL d27_reg_15_ ( .D(n5107), .SI(d27[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d27[15]) );
  SDFFRXL d27_reg_14_ ( .D(n5106), .SI(d27[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d27[14]) );
  SDFFRXL d27_reg_13_ ( .D(n5105), .SI(d27[12]), .SE(test_se), .CK(clk), .RN(
        n9094), .Q(d27[13]) );
  SDFFRXL d27_reg_12_ ( .D(n5104), .SI(d27[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d27[12]) );
  SDFFRXL d27_reg_11_ ( .D(n5103), .SI(d27[10]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d27[11]) );
  SDFFRXL d27_reg_10_ ( .D(n5102), .SI(d27[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d27[10]) );
  SDFFRXL d27_reg_9_ ( .D(n5101), .SI(d27[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d27[9]) );
  SDFFRXL d27_reg_8_ ( .D(n5100), .SI(d27[7]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d27[8]) );
  SDFFRXL d27_reg_7_ ( .D(n5099), .SI(d27[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d27[7]) );
  SDFFRXL d27_reg_6_ ( .D(n5098), .SI(d27[5]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d27[6]) );
  SDFFRXL d27_reg_5_ ( .D(n5097), .SI(d27[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d27[5]) );
  SDFFRXL d27_reg_4_ ( .D(n5096), .SI(d27[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d27[4]) );
  SDFFRXL d27_reg_3_ ( .D(n5095), .SI(d27[2]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d27[3]) );
  SDFFRXL d27_reg_2_ ( .D(n5094), .SI(d27[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d27[2]) );
  SDFFRXL d27_reg_1_ ( .D(n5093), .SI(d27[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d27[1]) );
  SDFFRXL d28_reg_35_ ( .D(n5091), .SI(d28[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d28[35]) );
  SDFFRXL d28_reg_34_ ( .D(n5090), .SI(d28[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d28[34]) );
  SDFFRXL d28_reg_33_ ( .D(n5089), .SI(d28[32]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d28[33]) );
  SDFFRXL d28_reg_32_ ( .D(n5088), .SI(d28[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d28[32]) );
  SDFFRXL d28_reg_31_ ( .D(n5087), .SI(d28[30]), .SE(test_se), .CK(clk), .RN(
        n9049), .Q(d28[31]) );
  SDFFRXL d28_reg_30_ ( .D(n5086), .SI(d28[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d28[30]) );
  SDFFRXL d28_reg_29_ ( .D(n5085), .SI(d28[28]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d28[29]) );
  SDFFRXL d28_reg_28_ ( .D(n5084), .SI(d28[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d28[28]) );
  SDFFRXL d28_reg_27_ ( .D(n5083), .SI(d28[26]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d28[27]) );
  SDFFRXL d28_reg_26_ ( .D(n5082), .SI(d28[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d28[26]) );
  SDFFRXL d28_reg_25_ ( .D(n5081), .SI(d28[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d28[25]) );
  SDFFRXL d28_reg_24_ ( .D(n5080), .SI(d28[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d28[24]) );
  SDFFRXL d28_reg_23_ ( .D(n5079), .SI(d28[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d28[23]) );
  SDFFRXL d28_reg_22_ ( .D(n5078), .SI(d28[21]), .SE(test_se), .CK(clk), .RN(
        n9072), .Q(d28[22]) );
  SDFFRXL d28_reg_21_ ( .D(n5077), .SI(d28[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d28[21]) );
  SDFFRXL d28_reg_20_ ( .D(n5076), .SI(d28[19]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d28[20]) );
  SDFFRXL d28_reg_19_ ( .D(n5075), .SI(d28[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d28[19]) );
  SDFFRXL d28_reg_18_ ( .D(n5074), .SI(d28[17]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d28[18]) );
  SDFFRXL d28_reg_17_ ( .D(n5073), .SI(d28[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d28[17]) );
  SDFFRXL d28_reg_16_ ( .D(n5072), .SI(d28[15]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d28[16]) );
  SDFFRXL d28_reg_15_ ( .D(n5071), .SI(d28[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d28[15]) );
  SDFFRXL d28_reg_14_ ( .D(n5070), .SI(d28[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d28[14]) );
  SDFFRXL d28_reg_13_ ( .D(n5069), .SI(d28[12]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d28[13]) );
  SDFFRXL d28_reg_12_ ( .D(n5068), .SI(d28[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d28[12]) );
  SDFFRXL d28_reg_11_ ( .D(n5067), .SI(d28[10]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d28[11]) );
  SDFFRXL d28_reg_10_ ( .D(n5066), .SI(d28[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d28[10]) );
  SDFFRXL d28_reg_9_ ( .D(n5065), .SI(d28[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d28[9]) );
  SDFFRXL d28_reg_8_ ( .D(n5064), .SI(d28[7]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d28[8]) );
  SDFFRXL d28_reg_7_ ( .D(n5063), .SI(d28[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d28[7]) );
  SDFFRXL d28_reg_6_ ( .D(n5062), .SI(d28[5]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d28[6]) );
  SDFFRXL d28_reg_5_ ( .D(n5061), .SI(d28[4]), .SE(test_se), .CK(clk), .RN(
        n9113), .Q(d28[5]) );
  SDFFRXL d28_reg_4_ ( .D(n5060), .SI(d28[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d28[4]) );
  SDFFRXL d28_reg_3_ ( .D(n5059), .SI(d28[2]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d28[3]) );
  SDFFRXL d28_reg_2_ ( .D(n5058), .SI(d28[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d28[2]) );
  SDFFRXL d28_reg_1_ ( .D(n5057), .SI(d28[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d28[1]) );
  SDFFRXL d29_reg_35_ ( .D(n5055), .SI(d29[34]), .SE(test_se), .CK(clk), .RN(
        n8924), .Q(d29[35]) );
  SDFFRXL d29_reg_34_ ( .D(n5054), .SI(d29[33]), .SE(test_se), .CK(clk), .RN(
        n8926), .Q(d29[34]) );
  SDFFRXL d29_reg_33_ ( .D(n5053), .SI(d29[32]), .SE(test_se), .CK(clk), .RN(
        n8928), .Q(d29[33]) );
  SDFFRXL d29_reg_32_ ( .D(n5052), .SI(d29[31]), .SE(test_se), .CK(clk), .RN(
        n8931), .Q(d29[32]) );
  SDFFRXL d29_reg_31_ ( .D(n5051), .SI(d29[30]), .SE(test_se), .CK(clk), .RN(
        n9049), .Q(d29[31]) );
  SDFFRXL d29_reg_30_ ( .D(n5050), .SI(d29[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d29[30]) );
  SDFFRXL d29_reg_29_ ( .D(n5049), .SI(d29[28]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d29[29]) );
  SDFFRXL d29_reg_28_ ( .D(n5048), .SI(d29[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d29[28]) );
  SDFFRXL d29_reg_27_ ( .D(n5047), .SI(d29[26]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d29[27]) );
  SDFFRXL d29_reg_26_ ( .D(n5046), .SI(d29[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d29[26]) );
  SDFFRXL d29_reg_25_ ( .D(n5045), .SI(d29[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d29[25]) );
  SDFFRXL d29_reg_24_ ( .D(n5044), .SI(d29[23]), .SE(test_se), .CK(clk), .RN(
        n9067), .Q(d29[24]) );
  SDFFRXL d29_reg_23_ ( .D(n5043), .SI(d29[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d29[23]) );
  SDFFRXL d29_reg_22_ ( .D(n5042), .SI(d29[21]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d29[22]) );
  SDFFRXL d29_reg_21_ ( .D(n5041), .SI(d29[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d29[21]) );
  SDFFRXL d29_reg_20_ ( .D(n5040), .SI(d29[19]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d29[20]) );
  SDFFRXL d29_reg_19_ ( .D(n5039), .SI(d29[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d29[19]) );
  SDFFRXL d29_reg_18_ ( .D(n5038), .SI(d29[17]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d29[18]) );
  SDFFRXL d29_reg_17_ ( .D(n5037), .SI(d29[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d29[17]) );
  SDFFRXL d29_reg_16_ ( .D(n5036), .SI(d29[15]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d29[16]) );
  SDFFRXL d29_reg_15_ ( .D(n5035), .SI(d29[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d29[15]) );
  SDFFRXL d29_reg_14_ ( .D(n5034), .SI(d29[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d29[14]) );
  SDFFRXL d29_reg_13_ ( .D(n5033), .SI(d29[12]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d29[13]) );
  SDFFRXL d29_reg_12_ ( .D(n5032), .SI(d29[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d29[12]) );
  SDFFRXL d29_reg_11_ ( .D(n5031), .SI(d29[10]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d29[11]) );
  SDFFRXL d29_reg_10_ ( .D(n5030), .SI(d29[9]), .SE(test_se), .CK(clk), .RN(
        n9101), .Q(d29[10]) );
  SDFFRXL d29_reg_9_ ( .D(n5029), .SI(d29[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d29[9]) );
  SDFFRXL d29_reg_8_ ( .D(n5028), .SI(d29[7]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d29[8]) );
  SDFFRXL d29_reg_7_ ( .D(n5027), .SI(d29[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d29[7]) );
  SDFFRXL d29_reg_6_ ( .D(n5026), .SI(d29[5]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d29[6]) );
  SDFFRXL d29_reg_5_ ( .D(n5025), .SI(d29[4]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d29[5]) );
  SDFFRXL d29_reg_4_ ( .D(n5024), .SI(d29[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d29[4]) );
  SDFFRXL d29_reg_3_ ( .D(n5023), .SI(d29[2]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d29[3]) );
  SDFFRXL d29_reg_2_ ( .D(n5022), .SI(d29[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d29[2]) );
  SDFFRXL d29_reg_1_ ( .D(n5021), .SI(d29[0]), .SE(test_se), .CK(clk), .RN(
        n9122), .Q(d29[1]) );
  SDFFRXL d30_reg_2_ ( .D(n5017), .SI(d30[1]), .SE(test_se), .CK(clk), .RN(
        n9120), .Q(d30[2]) );
  SDFFRXL d30_reg_3_ ( .D(n5016), .SI(d30[2]), .SE(test_se), .CK(clk), .RN(
        n9117), .Q(d30[3]) );
  SDFFRXL d30_reg_4_ ( .D(n5015), .SI(d30[3]), .SE(test_se), .CK(clk), .RN(
        n9115), .Q(d30[4]) );
  SDFFRXL d30_reg_5_ ( .D(n5014), .SI(d30[4]), .SE(test_se), .CK(clk), .RN(
        n9112), .Q(d30[5]) );
  SDFFRXL d30_reg_6_ ( .D(n5013), .SI(d30[5]), .SE(test_se), .CK(clk), .RN(
        n9110), .Q(d30[6]) );
  SDFFRXL d30_reg_7_ ( .D(n5012), .SI(d30[6]), .SE(test_se), .CK(clk), .RN(
        n9108), .Q(d30[7]) );
  SDFFRXL d30_reg_8_ ( .D(n5011), .SI(d30[7]), .SE(test_se), .CK(clk), .RN(
        n9105), .Q(d30[8]) );
  SDFFRXL d30_reg_9_ ( .D(n5010), .SI(d30[8]), .SE(test_se), .CK(clk), .RN(
        n9103), .Q(d30[9]) );
  SDFFRXL d30_reg_10_ ( .D(n5009), .SI(d30[9]), .SE(test_se), .CK(clk), .RN(
        n9100), .Q(d30[10]) );
  SDFFRXL d30_reg_11_ ( .D(n5008), .SI(d30[10]), .SE(test_se), .CK(clk), .RN(
        n9098), .Q(d30[11]) );
  SDFFRXL d30_reg_12_ ( .D(n5007), .SI(d30[11]), .SE(test_se), .CK(clk), .RN(
        n9096), .Q(d30[12]) );
  SDFFRXL d30_reg_13_ ( .D(n5006), .SI(d30[12]), .SE(test_se), .CK(clk), .RN(
        n9093), .Q(d30[13]) );
  SDFFRXL d30_reg_14_ ( .D(n5005), .SI(d30[13]), .SE(test_se), .CK(clk), .RN(
        n9091), .Q(d30[14]) );
  SDFFRXL d30_reg_15_ ( .D(n5004), .SI(d30[14]), .SE(test_se), .CK(clk), .RN(
        n9089), .Q(d30[15]) );
  SDFFRXL d30_reg_16_ ( .D(n5003), .SI(d30[15]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d30[16]) );
  SDFFRXL d30_reg_17_ ( .D(n5002), .SI(d30[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d30[17]) );
  SDFFRXL d30_reg_18_ ( .D(n5001), .SI(d30[17]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d30[18]) );
  SDFFRXL d30_reg_19_ ( .D(n5000), .SI(d30[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d30[19]) );
  SDFFRXL d30_reg_20_ ( .D(n4999), .SI(d30[19]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d30[20]) );
  SDFFRXL d30_reg_21_ ( .D(n4998), .SI(d30[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d30[21]) );
  SDFFRXL d30_reg_22_ ( .D(n4997), .SI(d30[21]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d30[22]) );
  SDFFRXL d30_reg_23_ ( .D(n4996), .SI(d30[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d30[23]) );
  SDFFRXL d30_reg_24_ ( .D(n4995), .SI(d30[23]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d30[24]) );
  SDFFRXL d30_reg_25_ ( .D(n4994), .SI(d30[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d30[25]) );
  SDFFRXL d30_reg_26_ ( .D(n4993), .SI(d30[25]), .SE(test_se), .CK(clk), .RN(
        n9062), .Q(d30[26]) );
  SDFFRXL d30_reg_27_ ( .D(n4992), .SI(d30[26]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d30[27]) );
  SDFFRXL d30_reg_28_ ( .D(n4991), .SI(d30[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d30[28]) );
  SDFFRXL d30_reg_29_ ( .D(n4990), .SI(d30[28]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d30[29]) );
  SDFFRXL d30_reg_30_ ( .D(n4989), .SI(d30[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d30[30]) );
  SDFFRXL d30_reg_31_ ( .D(n4988), .SI(d30[30]), .SE(test_se), .CK(clk), .RN(
        n9049), .Q(d30[31]) );
  SDFFRXL d31_reg_16_ ( .D(n4967), .SI(d31[15]), .SE(test_se), .CK(clk), .RN(
        n9086), .Q(d31[16]) );
  SDFFRXL d31_reg_17_ ( .D(n4966), .SI(d31[16]), .SE(test_se), .CK(clk), .RN(
        n9084), .Q(d31[17]) );
  SDFFRXL d31_reg_18_ ( .D(n4965), .SI(d31[17]), .SE(test_se), .CK(clk), .RN(
        n9081), .Q(d31[18]) );
  SDFFRXL d31_reg_19_ ( .D(n4964), .SI(d31[18]), .SE(test_se), .CK(clk), .RN(
        n9079), .Q(d31[19]) );
  SDFFRXL d31_reg_20_ ( .D(n4963), .SI(d31[19]), .SE(test_se), .CK(clk), .RN(
        n9076), .Q(d31[20]) );
  SDFFRXL d31_reg_21_ ( .D(n4962), .SI(d31[20]), .SE(test_se), .CK(clk), .RN(
        n9074), .Q(d31[21]) );
  SDFFRXL d31_reg_22_ ( .D(n4961), .SI(d31[21]), .SE(test_se), .CK(clk), .RN(
        n9071), .Q(d31[22]) );
  SDFFRXL d31_reg_23_ ( .D(n4960), .SI(d31[22]), .SE(test_se), .CK(clk), .RN(
        n9069), .Q(d31[23]) );
  SDFFRXL d31_reg_24_ ( .D(n4959), .SI(d31[23]), .SE(test_se), .CK(clk), .RN(
        n9066), .Q(d31[24]) );
  SDFFRXL d31_reg_25_ ( .D(n4958), .SI(d31[24]), .SE(test_se), .CK(clk), .RN(
        n9064), .Q(d31[25]) );
  SDFFRXL d31_reg_26_ ( .D(n4957), .SI(d31[25]), .SE(test_se), .CK(clk), .RN(
        n9061), .Q(d31[26]) );
  SDFFRXL d31_reg_27_ ( .D(n4956), .SI(d31[26]), .SE(test_se), .CK(clk), .RN(
        n9059), .Q(d31[27]) );
  SDFFRXL d31_reg_28_ ( .D(n4955), .SI(d31[27]), .SE(test_se), .CK(clk), .RN(
        n9057), .Q(d31[28]) );
  SDFFRXL d31_reg_29_ ( .D(n4954), .SI(d31[28]), .SE(test_se), .CK(clk), .RN(
        n9054), .Q(d31[29]) );
  SDFFRXL d31_reg_30_ ( .D(n4953), .SI(d31[29]), .SE(test_se), .CK(clk), .RN(
        n9052), .Q(d31[30]) );
  SDFFRXL d31_reg_31_ ( .D(n4952), .SI(d31[30]), .SE(test_se), .CK(clk), .RN(
        n9049), .Q(d31[31]) );
  SDFFRXL BF2II_a00_r_reg_0_ ( .D(n4800), .SI(N128), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(N130), .QN(n6110) );
  SDFFRXL BF2I_b_s_reg ( .D(counter[1]), .SI(n6247), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(BF2I_b_s), .QN(n6111) );
  SDFFRXL BF2I_a00_r_reg_0_ ( .D(n4928), .SI(n11091), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(BF2I_a_xr_n[0]), .QN(n1944) );
  SDFFRXL BF2I_b00_r_reg_0_ ( .D(n4678), .SI(BF2I_b_xi_n[31]), .SE(test_se), 
        .CK(clk), .RN(n9048), .Q(BF2I_b_xr_n[0]), .QN(n1725) );
  SDFFRXL BF2I_b00_i_reg_0_ ( .D(n4614), .SI(n6192), .SE(test_se), .CK(clk), 
        .RN(n9048), .Q(BF2I_b_xi_n[0]), .QN(n1661) );
  SDFFRXL fft_d14_reg_31_ ( .D(N1048), .SI(fft_d14[30]), .SE(test_se), .CK(clk), .RN(n8983), .Q(fft_d14[31]) );
  SDFFRXL fft_d14_reg_30_ ( .D(N1047), .SI(fft_d14[29]), .SE(test_se), .CK(clk), .RN(n8978), .Q(fft_d14[30]) );
  SDFFRXL fft_d14_reg_29_ ( .D(N1046), .SI(fft_d14[28]), .SE(test_se), .CK(clk), .RN(n8973), .Q(fft_d14[29]) );
  SDFFRXL fft_d14_reg_28_ ( .D(N1045), .SI(fft_d14[27]), .SE(test_se), .CK(clk), .RN(n8968), .Q(fft_d14[28]) );
  SDFFRXL fft_d14_reg_27_ ( .D(N1044), .SI(fft_d14[26]), .SE(test_se), .CK(clk), .RN(n8964), .Q(fft_d14[27]) );
  SDFFRXL fft_d14_reg_26_ ( .D(N1043), .SI(fft_d14[25]), .SE(test_se), .CK(clk), .RN(n8959), .Q(fft_d14[26]) );
  SDFFRXL fft_d14_reg_25_ ( .D(N1042), .SI(fft_d14[24]), .SE(test_se), .CK(clk), .RN(n8954), .Q(fft_d14[25]) );
  SDFFRXL fft_d14_reg_24_ ( .D(N1041), .SI(fft_d14[23]), .SE(test_se), .CK(clk), .RN(n8949), .Q(fft_d14[24]) );
  SDFFRXL fft_d14_reg_23_ ( .D(N1040), .SI(fft_d14[22]), .SE(test_se), .CK(clk), .RN(n8944), .Q(fft_d14[23]) );
  SDFFRXL fft_d14_reg_22_ ( .D(N1039), .SI(fft_d14[21]), .SE(test_se), .CK(clk), .RN(n8939), .Q(fft_d14[22]) );
  SDFFRXL fft_d14_reg_21_ ( .D(N1038), .SI(fft_d14[20]), .SE(test_se), .CK(clk), .RN(n8991), .Q(fft_d14[21]) );
  SDFFRXL fft_d14_reg_20_ ( .D(N1037), .SI(fft_d14[19]), .SE(test_se), .CK(clk), .RN(n8996), .Q(fft_d14[20]) );
  SDFFRXL fft_d14_reg_19_ ( .D(N1036), .SI(fft_d14[18]), .SE(test_se), .CK(clk), .RN(n9002), .Q(fft_d14[19]) );
  SDFFRXL fft_d14_reg_18_ ( .D(N1035), .SI(fft_d14[17]), .SE(test_se), .CK(clk), .RN(n9007), .Q(fft_d14[18]) );
  SDFFRXL fft_d14_reg_17_ ( .D(N1034), .SI(fft_d14[16]), .SE(test_se), .CK(clk), .RN(n9012), .Q(fft_d14[17]) );
  SDFFRXL fft_d14_reg_16_ ( .D(N1033), .SI(fft_d14[15]), .SE(test_se), .CK(clk), .RN(n9017), .Q(fft_d14[16]) );
  SDFFRXL fft_d14_reg_15_ ( .D(N1032), .SI(fft_d14[14]), .SE(test_se), .CK(clk), .RN(n8981), .Q(fft_d14[15]) );
  SDFFRXL fft_d14_reg_14_ ( .D(N1031), .SI(fft_d14[13]), .SE(test_se), .CK(clk), .RN(n8976), .Q(fft_d14[14]) );
  SDFFRXL fft_d14_reg_13_ ( .D(N1030), .SI(fft_d14[12]), .SE(test_se), .CK(clk), .RN(n8971), .Q(fft_d14[13]) );
  SDFFRXL fft_d14_reg_12_ ( .D(N1029), .SI(fft_d14[11]), .SE(test_se), .CK(clk), .RN(n8966), .Q(fft_d14[12]) );
  SDFFRXL fft_d14_reg_11_ ( .D(N1028), .SI(fft_d14[10]), .SE(test_se), .CK(clk), .RN(n8961), .Q(fft_d14[11]) );
  SDFFRXL fft_d14_reg_10_ ( .D(N1027), .SI(fft_d14[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d14[10]) );
  SDFFRXL fft_d14_reg_9_ ( .D(N1026), .SI(fft_d14[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d14[9]) );
  SDFFRXL fft_d14_reg_8_ ( .D(N1025), .SI(fft_d14[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d14[8]) );
  SDFFRXL fft_d14_reg_7_ ( .D(N1024), .SI(fft_d14[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d14[7]) );
  SDFFRXL fft_d14_reg_6_ ( .D(N1023), .SI(fft_d14[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d14[6]) );
  SDFFRXL fft_d14_reg_5_ ( .D(N1022), .SI(fft_d14[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d14[5]) );
  SDFFRXL fft_d14_reg_4_ ( .D(N1021), .SI(fft_d14[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d14[4]) );
  SDFFRXL fft_d14_reg_3_ ( .D(N1020), .SI(fft_d14[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d14[3]) );
  SDFFRXL fft_d14_reg_2_ ( .D(N1019), .SI(fft_d14[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d14[2]) );
  SDFFRXL fft_d14_reg_1_ ( .D(N1018), .SI(fft_d14[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d14[1]) );
  SDFFRXL fft_d14_reg_0_ ( .D(N1017), .SI(n10514), .SE(test_se), .CK(clk), 
        .RN(n9015), .Q(fft_d14[0]) );
  SDFFRXL fft_d15_reg_31_ ( .D(N1080), .SI(fft_d15[30]), .SE(test_se), .CK(clk), .RN(n8983), .Q(fft_d15[31]) );
  SDFFRXL fft_d15_reg_30_ ( .D(N1079), .SI(fft_d15[29]), .SE(test_se), .CK(clk), .RN(n8978), .Q(fft_d15[30]) );
  SDFFRXL fft_d15_reg_29_ ( .D(N1078), .SI(fft_d15[28]), .SE(test_se), .CK(clk), .RN(n8973), .Q(fft_d15[29]) );
  SDFFRXL fft_d15_reg_28_ ( .D(N1077), .SI(fft_d15[27]), .SE(test_se), .CK(clk), .RN(n8968), .Q(fft_d15[28]) );
  SDFFRXL fft_d15_reg_27_ ( .D(N1076), .SI(fft_d15[26]), .SE(test_se), .CK(clk), .RN(n8963), .Q(fft_d15[27]) );
  SDFFRXL fft_d15_reg_26_ ( .D(N1075), .SI(fft_d15[25]), .SE(test_se), .CK(clk), .RN(n8958), .Q(fft_d15[26]) );
  SDFFRXL fft_d15_reg_25_ ( .D(N1074), .SI(fft_d15[24]), .SE(test_se), .CK(clk), .RN(n8953), .Q(fft_d15[25]) );
  SDFFRXL fft_d15_reg_24_ ( .D(N1073), .SI(fft_d15[23]), .SE(test_se), .CK(clk), .RN(n8948), .Q(fft_d15[24]) );
  SDFFRXL fft_d15_reg_23_ ( .D(N1072), .SI(fft_d15[22]), .SE(test_se), .CK(clk), .RN(n8943), .Q(fft_d15[23]) );
  SDFFRXL fft_d15_reg_22_ ( .D(N1071), .SI(fft_d15[21]), .SE(test_se), .CK(clk), .RN(n8938), .Q(fft_d15[22]) );
  SDFFRXL fft_d15_reg_21_ ( .D(N1070), .SI(fft_d15[20]), .SE(test_se), .CK(clk), .RN(n8991), .Q(fft_d15[21]) );
  SDFFRXL fft_d15_reg_20_ ( .D(N1069), .SI(fft_d15[19]), .SE(test_se), .CK(clk), .RN(n8996), .Q(fft_d15[20]) );
  SDFFRXL fft_d15_reg_19_ ( .D(N1068), .SI(fft_d15[18]), .SE(test_se), .CK(clk), .RN(n9001), .Q(fft_d15[19]) );
  SDFFRXL fft_d15_reg_18_ ( .D(N1067), .SI(fft_d15[17]), .SE(test_se), .CK(clk), .RN(n9006), .Q(fft_d15[18]) );
  SDFFRXL fft_d15_reg_17_ ( .D(N1066), .SI(fft_d15[16]), .SE(test_se), .CK(clk), .RN(n9012), .Q(fft_d15[17]) );
  SDFFRXL fft_d15_reg_16_ ( .D(N1065), .SI(fft_d15[15]), .SE(test_se), .CK(clk), .RN(n9017), .Q(fft_d15[16]) );
  SDFFRXL fft_d15_reg_15_ ( .D(N1064), .SI(fft_d15[14]), .SE(test_se), .CK(clk), .RN(n8980), .Q(fft_d15[15]) );
  SDFFRXL fft_d15_reg_14_ ( .D(N1063), .SI(fft_d15[13]), .SE(test_se), .CK(clk), .RN(n8975), .Q(fft_d15[14]) );
  SDFFRXL fft_d15_reg_13_ ( .D(N1062), .SI(fft_d15[12]), .SE(test_se), .CK(clk), .RN(n8970), .Q(fft_d15[13]) );
  SDFFRXL fft_d15_reg_12_ ( .D(N1061), .SI(fft_d15[11]), .SE(test_se), .CK(clk), .RN(n8965), .Q(fft_d15[12]) );
  SDFFRXL fft_d15_reg_11_ ( .D(N1060), .SI(fft_d15[10]), .SE(test_se), .CK(clk), .RN(n8960), .Q(fft_d15[11]) );
  SDFFRXL fft_d15_reg_10_ ( .D(N1059), .SI(fft_d15[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d15[10]) );
  SDFFRXL fft_d15_reg_9_ ( .D(N1058), .SI(fft_d15[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d15[9]) );
  SDFFRXL fft_d15_reg_8_ ( .D(N1057), .SI(fft_d15[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d15[8]) );
  SDFFRXL fft_d15_reg_7_ ( .D(N1056), .SI(fft_d15[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d15[7]) );
  SDFFRXL fft_d15_reg_6_ ( .D(N1055), .SI(fft_d15[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d15[6]) );
  SDFFRXL fft_d15_reg_5_ ( .D(N1054), .SI(fft_d15[4]), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(fft_d15[5]) );
  SDFFRXL fft_d15_reg_4_ ( .D(N1053), .SI(fft_d15[3]), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(fft_d15[4]) );
  SDFFRXL fft_d15_reg_3_ ( .D(N1052), .SI(fft_d15[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d15[3]) );
  SDFFRXL fft_d15_reg_2_ ( .D(N1051), .SI(fft_d15[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d15[2]) );
  SDFFRXL fft_d15_reg_1_ ( .D(N1050), .SI(fft_d15[0]), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(fft_d15[1]) );
  SDFFRXL fft_d15_reg_0_ ( .D(N1049), .SI(fft_d15_q[31]), .SE(test_se), .CK(
        clk), .RN(n9014), .Q(fft_d15[0]) );
  SDFFRXL fft_valid_reg ( .D(n10478), .SI(n10482), .SE(test_se), .CK(clk), 
        .RN(n9127), .Q(fft_valid) );
  SDFFRXL fft_d0_reg_31_ ( .D(N600), .SI(fft_d0[30]), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(fft_d0[31]) );
  SDFFRXL fft_d0_reg_30_ ( .D(N599), .SI(fft_d0[29]), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(fft_d0[30]) );
  SDFFRXL fft_d0_reg_29_ ( .D(N598), .SI(fft_d0[28]), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(fft_d0[29]) );
  SDFFRXL fft_d0_reg_28_ ( .D(N597), .SI(fft_d0[27]), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(fft_d0[28]) );
  SDFFRXL fft_d0_reg_27_ ( .D(N596), .SI(fft_d0[26]), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(fft_d0[27]) );
  SDFFRXL fft_d0_reg_26_ ( .D(N595), .SI(fft_d0[25]), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(fft_d0[26]) );
  SDFFRXL fft_d0_reg_25_ ( .D(N594), .SI(fft_d0[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d0[25]) );
  SDFFRXL fft_d0_reg_24_ ( .D(N593), .SI(fft_d0[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d0[24]) );
  SDFFRXL fft_d0_reg_23_ ( .D(N592), .SI(fft_d0[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d0[23]) );
  SDFFRXL fft_d0_reg_22_ ( .D(N591), .SI(fft_d0[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d0[22]) );
  SDFFRXL fft_d0_reg_21_ ( .D(N590), .SI(fft_d0[20]), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(fft_d0[21]) );
  SDFFRXL fft_d0_reg_20_ ( .D(N589), .SI(fft_d0[19]), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(fft_d0[20]) );
  SDFFRXL fft_d0_reg_19_ ( .D(N588), .SI(fft_d0[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d0[19]) );
  SDFFRXL fft_d0_reg_18_ ( .D(N587), .SI(fft_d0[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d0[18]) );
  SDFFRXL fft_d0_reg_17_ ( .D(N586), .SI(fft_d0[16]), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(fft_d0[17]) );
  SDFFRXL fft_d0_reg_16_ ( .D(N585), .SI(fft_d0[15]), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(fft_d0[16]) );
  SDFFRXL fft_d0_reg_15_ ( .D(N584), .SI(fft_d0[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d0[15]) );
  SDFFRXL fft_d0_reg_14_ ( .D(N583), .SI(fft_d0[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d0[14]) );
  SDFFRXL fft_d0_reg_13_ ( .D(N582), .SI(fft_d0[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d0[13]) );
  SDFFRXL fft_d0_reg_12_ ( .D(N581), .SI(fft_d0[11]), .SE(test_se), .CK(clk), 
        .RN(n8967), .Q(fft_d0[12]) );
  SDFFRXL fft_d0_reg_11_ ( .D(N580), .SI(fft_d0[10]), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(fft_d0[11]) );
  SDFFRXL fft_d0_reg_10_ ( .D(N579), .SI(fft_d0[9]), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(fft_d0[10]) );
  SDFFRXL fft_d0_reg_9_ ( .D(N578), .SI(fft_d0[8]), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(fft_d0[9]) );
  SDFFRXL fft_d0_reg_8_ ( .D(N577), .SI(fft_d0[7]), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(fft_d0[8]) );
  SDFFRXL fft_d0_reg_7_ ( .D(N576), .SI(fft_d0[6]), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(fft_d0[7]) );
  SDFFRXL fft_d0_reg_6_ ( .D(N575), .SI(fft_d0[5]), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(fft_d0[6]) );
  SDFFRXL fft_d0_reg_5_ ( .D(N574), .SI(fft_d0[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d0[5]) );
  SDFFRXL fft_d0_reg_4_ ( .D(N573), .SI(fft_d0[3]), .SE(test_se), .CK(clk), 
        .RN(n8995), .Q(fft_d0[4]) );
  SDFFRXL fft_d0_reg_3_ ( .D(N572), .SI(fft_d0[2]), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(fft_d0[3]) );
  SDFFRXL fft_d0_reg_2_ ( .D(N571), .SI(fft_d0[1]), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(fft_d0[2]) );
  SDFFRXL fft_d0_reg_1_ ( .D(N570), .SI(fft_d0[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d0[1]) );
  SDFFRXL fft_d0_reg_0_ ( .D(N569), .SI(n10962), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d0[0]) );
  SDFFRXL fft_d1_reg_31_ ( .D(N632), .SI(fft_d1[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d1[31]) );
  SDFFRXL fft_d1_reg_30_ ( .D(N631), .SI(fft_d1[29]), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(fft_d1[30]) );
  SDFFRXL fft_d1_reg_29_ ( .D(N630), .SI(fft_d1[28]), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(fft_d1[29]) );
  SDFFRXL fft_d1_reg_28_ ( .D(N629), .SI(fft_d1[27]), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(fft_d1[28]) );
  SDFFRXL fft_d1_reg_27_ ( .D(N628), .SI(fft_d1[26]), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(fft_d1[27]) );
  SDFFRXL fft_d1_reg_26_ ( .D(N627), .SI(fft_d1[25]), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(fft_d1[26]) );
  SDFFRXL fft_d1_reg_25_ ( .D(N626), .SI(fft_d1[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d1[25]) );
  SDFFRXL fft_d1_reg_24_ ( .D(N625), .SI(fft_d1[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d1[24]) );
  SDFFRXL fft_d1_reg_23_ ( .D(N624), .SI(fft_d1[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d1[23]) );
  SDFFRXL fft_d1_reg_22_ ( .D(N623), .SI(fft_d1[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d1[22]) );
  SDFFRXL fft_d1_reg_21_ ( .D(N622), .SI(fft_d1[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d1[21]) );
  SDFFRXL fft_d1_reg_20_ ( .D(N621), .SI(fft_d1[19]), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(fft_d1[20]) );
  SDFFRXL fft_d1_reg_19_ ( .D(N620), .SI(fft_d1[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d1[19]) );
  SDFFRXL fft_d1_reg_18_ ( .D(N619), .SI(fft_d1[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d1[18]) );
  SDFFRXL fft_d1_reg_17_ ( .D(N618), .SI(fft_d1[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d1[17]) );
  SDFFRXL fft_d1_reg_16_ ( .D(N617), .SI(fft_d1[15]), .SE(test_se), .CK(clk), 
        .RN(n9017), .Q(fft_d1[16]) );
  SDFFRXL fft_d1_reg_15_ ( .D(N616), .SI(fft_d1[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d1[15]) );
  SDFFRXL fft_d1_reg_14_ ( .D(N615), .SI(fft_d1[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d1[14]) );
  SDFFRXL fft_d1_reg_13_ ( .D(N614), .SI(fft_d1[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d1[13]) );
  SDFFRXL fft_d1_reg_12_ ( .D(N613), .SI(fft_d1[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d1[12]) );
  SDFFRXL fft_d1_reg_11_ ( .D(N612), .SI(fft_d1[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d1[11]) );
  SDFFRXL fft_d1_reg_10_ ( .D(N611), .SI(fft_d1[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d1[10]) );
  SDFFRXL fft_d1_reg_9_ ( .D(N610), .SI(fft_d1[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d1[9]) );
  SDFFRXL fft_d1_reg_8_ ( .D(N609), .SI(fft_d1[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d1[8]) );
  SDFFRXL fft_d1_reg_7_ ( .D(N608), .SI(fft_d1[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d1[7]) );
  SDFFRXL fft_d1_reg_6_ ( .D(N607), .SI(fft_d1[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d1[6]) );
  SDFFRXL fft_d1_reg_5_ ( .D(N606), .SI(fft_d1[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d1[5]) );
  SDFFRXL fft_d1_reg_4_ ( .D(N605), .SI(fft_d1[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d1[4]) );
  SDFFRXL fft_d1_reg_3_ ( .D(N604), .SI(fft_d1[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d1[3]) );
  SDFFRXL fft_d1_reg_2_ ( .D(N603), .SI(fft_d1[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d1[2]) );
  SDFFRXL fft_d1_reg_1_ ( .D(N602), .SI(fft_d1[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d1[1]) );
  SDFFRXL fft_d1_reg_0_ ( .D(N601), .SI(n10930), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d1[0]) );
  SDFFRXL fft_d2_reg_31_ ( .D(N664), .SI(fft_d2[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d2[31]) );
  SDFFRXL fft_d2_reg_30_ ( .D(N663), .SI(fft_d2[29]), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(fft_d2[30]) );
  SDFFRXL fft_d2_reg_29_ ( .D(N662), .SI(fft_d2[28]), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(fft_d2[29]) );
  SDFFRXL fft_d2_reg_28_ ( .D(N661), .SI(fft_d2[27]), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(fft_d2[28]) );
  SDFFRXL fft_d2_reg_27_ ( .D(N660), .SI(fft_d2[26]), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(fft_d2[27]) );
  SDFFRXL fft_d2_reg_26_ ( .D(N659), .SI(fft_d2[25]), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(fft_d2[26]) );
  SDFFRXL fft_d2_reg_25_ ( .D(N658), .SI(fft_d2[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d2[25]) );
  SDFFRXL fft_d2_reg_24_ ( .D(N657), .SI(fft_d2[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d2[24]) );
  SDFFRXL fft_d2_reg_23_ ( .D(N656), .SI(fft_d2[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d2[23]) );
  SDFFRXL fft_d2_reg_22_ ( .D(N655), .SI(fft_d2[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d2[22]) );
  SDFFRXL fft_d2_reg_21_ ( .D(N654), .SI(fft_d2[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d2[21]) );
  SDFFRXL fft_d2_reg_20_ ( .D(N653), .SI(fft_d2[19]), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(fft_d2[20]) );
  SDFFRXL fft_d2_reg_19_ ( .D(N652), .SI(fft_d2[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d2[19]) );
  SDFFRXL fft_d2_reg_18_ ( .D(N651), .SI(fft_d2[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d2[18]) );
  SDFFRXL fft_d2_reg_17_ ( .D(N650), .SI(fft_d2[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d2[17]) );
  SDFFRXL fft_d2_reg_16_ ( .D(N649), .SI(fft_d2[15]), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(fft_d2[16]) );
  SDFFRXL fft_d2_reg_15_ ( .D(N648), .SI(fft_d2[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d2[15]) );
  SDFFRXL fft_d2_reg_14_ ( .D(N647), .SI(fft_d2[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d2[14]) );
  SDFFRXL fft_d2_reg_13_ ( .D(N646), .SI(fft_d2[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d2[13]) );
  SDFFRXL fft_d2_reg_12_ ( .D(N645), .SI(fft_d2[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d2[12]) );
  SDFFRXL fft_d2_reg_11_ ( .D(N644), .SI(fft_d2[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d2[11]) );
  SDFFRXL fft_d2_reg_10_ ( .D(N643), .SI(fft_d2[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d2[10]) );
  SDFFRXL fft_d2_reg_9_ ( .D(N642), .SI(fft_d2[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d2[9]) );
  SDFFRXL fft_d2_reg_8_ ( .D(N641), .SI(fft_d2[7]), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(fft_d2[8]) );
  SDFFRXL fft_d2_reg_7_ ( .D(N640), .SI(fft_d2[6]), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(fft_d2[7]) );
  SDFFRXL fft_d2_reg_6_ ( .D(N639), .SI(fft_d2[5]), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(fft_d2[6]) );
  SDFFRXL fft_d2_reg_5_ ( .D(N638), .SI(fft_d2[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d2[5]) );
  SDFFRXL fft_d2_reg_4_ ( .D(N637), .SI(fft_d2[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d2[4]) );
  SDFFRXL fft_d2_reg_3_ ( .D(N636), .SI(fft_d2[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d2[3]) );
  SDFFRXL fft_d2_reg_2_ ( .D(N635), .SI(fft_d2[1]), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(fft_d2[2]) );
  SDFFRXL fft_d2_reg_1_ ( .D(N634), .SI(fft_d2[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d2[1]) );
  SDFFRXL fft_d2_reg_0_ ( .D(N633), .SI(n10898), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d2[0]) );
  SDFFRXL fft_d3_reg_31_ ( .D(N696), .SI(fft_d3[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d3[31]) );
  SDFFRXL fft_d3_reg_30_ ( .D(N695), .SI(fft_d3[29]), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(fft_d3[30]) );
  SDFFRXL fft_d3_reg_29_ ( .D(N694), .SI(fft_d3[28]), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(fft_d3[29]) );
  SDFFRXL fft_d3_reg_28_ ( .D(N693), .SI(fft_d3[27]), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(fft_d3[28]) );
  SDFFRXL fft_d3_reg_27_ ( .D(N692), .SI(fft_d3[26]), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(fft_d3[27]) );
  SDFFRXL fft_d3_reg_26_ ( .D(N691), .SI(fft_d3[25]), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(fft_d3[26]) );
  SDFFRXL fft_d3_reg_25_ ( .D(N690), .SI(fft_d3[24]), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(fft_d3[25]) );
  SDFFRXL fft_d3_reg_24_ ( .D(N689), .SI(fft_d3[23]), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(fft_d3[24]) );
  SDFFRXL fft_d3_reg_23_ ( .D(N688), .SI(fft_d3[22]), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(fft_d3[23]) );
  SDFFRXL fft_d3_reg_22_ ( .D(N687), .SI(fft_d3[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d3[22]) );
  SDFFRXL fft_d3_reg_21_ ( .D(N686), .SI(fft_d3[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d3[21]) );
  SDFFRXL fft_d3_reg_20_ ( .D(N685), .SI(fft_d3[19]), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(fft_d3[20]) );
  SDFFRXL fft_d3_reg_19_ ( .D(N684), .SI(fft_d3[18]), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(fft_d3[19]) );
  SDFFRXL fft_d3_reg_18_ ( .D(N683), .SI(fft_d3[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d3[18]) );
  SDFFRXL fft_d3_reg_17_ ( .D(N682), .SI(fft_d3[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d3[17]) );
  SDFFRXL fft_d3_reg_16_ ( .D(N681), .SI(fft_d3[15]), .SE(test_se), .CK(clk), 
        .RN(n9017), .Q(fft_d3[16]) );
  SDFFRXL fft_d3_reg_15_ ( .D(N680), .SI(fft_d3[14]), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(fft_d3[15]) );
  SDFFRXL fft_d3_reg_14_ ( .D(N679), .SI(fft_d3[13]), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(fft_d3[14]) );
  SDFFRXL fft_d3_reg_13_ ( .D(N678), .SI(fft_d3[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d3[13]) );
  SDFFRXL fft_d3_reg_12_ ( .D(N677), .SI(fft_d3[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d3[12]) );
  SDFFRXL fft_d3_reg_11_ ( .D(N676), .SI(fft_d3[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d3[11]) );
  SDFFRXL fft_d3_reg_10_ ( .D(N675), .SI(fft_d3[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d3[10]) );
  SDFFRXL fft_d3_reg_9_ ( .D(N674), .SI(fft_d3[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d3[9]) );
  SDFFRXL fft_d3_reg_8_ ( .D(N673), .SI(fft_d3[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d3[8]) );
  SDFFRXL fft_d3_reg_7_ ( .D(N672), .SI(fft_d3[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d3[7]) );
  SDFFRXL fft_d3_reg_6_ ( .D(N671), .SI(fft_d3[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d3[6]) );
  SDFFRXL fft_d3_reg_5_ ( .D(N670), .SI(fft_d3[4]), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(fft_d3[5]) );
  SDFFRXL fft_d3_reg_4_ ( .D(N669), .SI(fft_d3[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d3[4]) );
  SDFFRXL fft_d3_reg_3_ ( .D(N668), .SI(fft_d3[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d3[3]) );
  SDFFRXL fft_d3_reg_2_ ( .D(N667), .SI(fft_d3[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d3[2]) );
  SDFFRXL fft_d3_reg_1_ ( .D(N666), .SI(fft_d3[0]), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(fft_d3[1]) );
  SDFFRXL fft_d3_reg_0_ ( .D(N665), .SI(n10866), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d3[0]) );
  SDFFRXL fft_d4_reg_31_ ( .D(N728), .SI(fft_d4[30]), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(fft_d4[31]) );
  SDFFRXL fft_d4_reg_30_ ( .D(N727), .SI(fft_d4[29]), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(fft_d4[30]) );
  SDFFRXL fft_d4_reg_29_ ( .D(N726), .SI(fft_d4[28]), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(fft_d4[29]) );
  SDFFRXL fft_d4_reg_28_ ( .D(N725), .SI(fft_d4[27]), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(fft_d4[28]) );
  SDFFRXL fft_d4_reg_27_ ( .D(N724), .SI(fft_d4[26]), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(fft_d4[27]) );
  SDFFRXL fft_d4_reg_26_ ( .D(N723), .SI(fft_d4[25]), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(fft_d4[26]) );
  SDFFRXL fft_d4_reg_25_ ( .D(N722), .SI(fft_d4[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d4[25]) );
  SDFFRXL fft_d4_reg_24_ ( .D(N721), .SI(fft_d4[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d4[24]) );
  SDFFRXL fft_d4_reg_23_ ( .D(N720), .SI(fft_d4[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d4[23]) );
  SDFFRXL fft_d4_reg_22_ ( .D(N719), .SI(fft_d4[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d4[22]) );
  SDFFRXL fft_d4_reg_21_ ( .D(N718), .SI(fft_d4[20]), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(fft_d4[21]) );
  SDFFRXL fft_d4_reg_20_ ( .D(N717), .SI(fft_d4[19]), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(fft_d4[20]) );
  SDFFRXL fft_d4_reg_19_ ( .D(N716), .SI(fft_d4[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d4[19]) );
  SDFFRXL fft_d4_reg_18_ ( .D(N715), .SI(fft_d4[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d4[18]) );
  SDFFRXL fft_d4_reg_17_ ( .D(N714), .SI(fft_d4[16]), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(fft_d4[17]) );
  SDFFRXL fft_d4_reg_16_ ( .D(N713), .SI(fft_d4[15]), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(fft_d4[16]) );
  SDFFRXL fft_d4_reg_15_ ( .D(N712), .SI(fft_d4[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d4[15]) );
  SDFFRXL fft_d4_reg_14_ ( .D(N711), .SI(fft_d4[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d4[14]) );
  SDFFRXL fft_d4_reg_13_ ( .D(N710), .SI(fft_d4[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d4[13]) );
  SDFFRXL fft_d4_reg_12_ ( .D(N709), .SI(fft_d4[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d4[12]) );
  SDFFRXL fft_d4_reg_11_ ( .D(N708), .SI(fft_d4[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d4[11]) );
  SDFFRXL fft_d4_reg_10_ ( .D(N707), .SI(fft_d4[9]), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(fft_d4[10]) );
  SDFFRXL fft_d4_reg_9_ ( .D(N706), .SI(fft_d4[8]), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(fft_d4[9]) );
  SDFFRXL fft_d4_reg_8_ ( .D(N705), .SI(fft_d4[7]), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(fft_d4[8]) );
  SDFFRXL fft_d4_reg_7_ ( .D(N704), .SI(fft_d4[6]), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(fft_d4[7]) );
  SDFFRXL fft_d4_reg_6_ ( .D(N703), .SI(fft_d4[5]), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(fft_d4[6]) );
  SDFFRXL fft_d4_reg_5_ ( .D(N702), .SI(fft_d4[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d4[5]) );
  SDFFRXL fft_d4_reg_4_ ( .D(N701), .SI(fft_d4[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d4[4]) );
  SDFFRXL fft_d4_reg_3_ ( .D(N700), .SI(fft_d4[2]), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(fft_d4[3]) );
  SDFFRXL fft_d4_reg_2_ ( .D(N699), .SI(fft_d4[1]), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(fft_d4[2]) );
  SDFFRXL fft_d4_reg_1_ ( .D(N698), .SI(fft_d4[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d4[1]) );
  SDFFRXL fft_d4_reg_0_ ( .D(N697), .SI(n10834), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d4[0]) );
  SDFFRXL fft_d5_reg_31_ ( .D(N760), .SI(fft_d5[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d5[31]) );
  SDFFRXL fft_d5_reg_30_ ( .D(N759), .SI(fft_d5[29]), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(fft_d5[30]) );
  SDFFRXL fft_d5_reg_29_ ( .D(N758), .SI(fft_d5[28]), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(fft_d5[29]) );
  SDFFRXL fft_d5_reg_28_ ( .D(N757), .SI(fft_d5[27]), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(fft_d5[28]) );
  SDFFRXL fft_d5_reg_27_ ( .D(N756), .SI(fft_d5[26]), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(fft_d5[27]) );
  SDFFRXL fft_d5_reg_26_ ( .D(N755), .SI(fft_d5[25]), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(fft_d5[26]) );
  SDFFRXL fft_d5_reg_25_ ( .D(N754), .SI(fft_d5[24]), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(fft_d5[25]) );
  SDFFRXL fft_d5_reg_24_ ( .D(N753), .SI(fft_d5[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d5[24]) );
  SDFFRXL fft_d5_reg_23_ ( .D(N752), .SI(fft_d5[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d5[23]) );
  SDFFRXL fft_d5_reg_22_ ( .D(N751), .SI(fft_d5[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d5[22]) );
  SDFFRXL fft_d5_reg_21_ ( .D(N750), .SI(fft_d5[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d5[21]) );
  SDFFRXL fft_d5_reg_20_ ( .D(N749), .SI(fft_d5[19]), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(fft_d5[20]) );
  SDFFRXL fft_d5_reg_19_ ( .D(N748), .SI(fft_d5[18]), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(fft_d5[19]) );
  SDFFRXL fft_d5_reg_18_ ( .D(N747), .SI(fft_d5[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d5[18]) );
  SDFFRXL fft_d5_reg_17_ ( .D(N746), .SI(fft_d5[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d5[17]) );
  SDFFRXL fft_d5_reg_16_ ( .D(N745), .SI(fft_d5[15]), .SE(test_se), .CK(clk), 
        .RN(n9017), .Q(fft_d5[16]) );
  SDFFRXL fft_d5_reg_15_ ( .D(N744), .SI(fft_d5[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d5[15]) );
  SDFFRXL fft_d5_reg_14_ ( .D(N743), .SI(fft_d5[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d5[14]) );
  SDFFRXL fft_d5_reg_13_ ( .D(N742), .SI(fft_d5[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d5[13]) );
  SDFFRXL fft_d5_reg_12_ ( .D(N741), .SI(fft_d5[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d5[12]) );
  SDFFRXL fft_d5_reg_11_ ( .D(N740), .SI(fft_d5[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d5[11]) );
  SDFFRXL fft_d5_reg_10_ ( .D(N739), .SI(fft_d5[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d5[10]) );
  SDFFRXL fft_d5_reg_9_ ( .D(N738), .SI(fft_d5[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d5[9]) );
  SDFFRXL fft_d5_reg_8_ ( .D(N737), .SI(fft_d5[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d5[8]) );
  SDFFRXL fft_d5_reg_7_ ( .D(N736), .SI(fft_d5[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d5[7]) );
  SDFFRXL fft_d5_reg_6_ ( .D(N735), .SI(fft_d5[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d5[6]) );
  SDFFRXL fft_d5_reg_5_ ( .D(N734), .SI(fft_d5[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d5[5]) );
  SDFFRXL fft_d5_reg_4_ ( .D(N733), .SI(fft_d5[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d5[4]) );
  SDFFRXL fft_d5_reg_3_ ( .D(N732), .SI(fft_d5[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d5[3]) );
  SDFFRXL fft_d5_reg_2_ ( .D(N731), .SI(fft_d5[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d5[2]) );
  SDFFRXL fft_d5_reg_1_ ( .D(N730), .SI(fft_d5[0]), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(fft_d5[1]) );
  SDFFRXL fft_d5_reg_0_ ( .D(N729), .SI(n10802), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d5[0]) );
  SDFFRXL fft_d6_reg_31_ ( .D(N792), .SI(fft_d6[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d6[31]) );
  SDFFRXL fft_d6_reg_30_ ( .D(N791), .SI(fft_d6[29]), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(fft_d6[30]) );
  SDFFRXL fft_d6_reg_29_ ( .D(N790), .SI(fft_d6[28]), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(fft_d6[29]) );
  SDFFRXL fft_d6_reg_28_ ( .D(N789), .SI(fft_d6[27]), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(fft_d6[28]) );
  SDFFRXL fft_d6_reg_27_ ( .D(N788), .SI(fft_d6[26]), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(fft_d6[27]) );
  SDFFRXL fft_d6_reg_26_ ( .D(N787), .SI(fft_d6[25]), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(fft_d6[26]) );
  SDFFRXL fft_d6_reg_25_ ( .D(N786), .SI(fft_d6[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d6[25]) );
  SDFFRXL fft_d6_reg_24_ ( .D(N785), .SI(fft_d6[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d6[24]) );
  SDFFRXL fft_d6_reg_23_ ( .D(N784), .SI(fft_d6[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d6[23]) );
  SDFFRXL fft_d6_reg_22_ ( .D(N783), .SI(fft_d6[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d6[22]) );
  SDFFRXL fft_d6_reg_21_ ( .D(N782), .SI(fft_d6[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d6[21]) );
  SDFFRXL fft_d6_reg_20_ ( .D(N781), .SI(fft_d6[19]), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(fft_d6[20]) );
  SDFFRXL fft_d6_reg_19_ ( .D(N780), .SI(fft_d6[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d6[19]) );
  SDFFRXL fft_d6_reg_18_ ( .D(N779), .SI(fft_d6[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d6[18]) );
  SDFFRXL fft_d6_reg_17_ ( .D(N778), .SI(fft_d6[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d6[17]) );
  SDFFRXL fft_d6_reg_16_ ( .D(N777), .SI(fft_d6[15]), .SE(test_se), .CK(clk), 
        .RN(n9017), .Q(fft_d6[16]) );
  SDFFRXL fft_d6_reg_15_ ( .D(N776), .SI(fft_d6[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d6[15]) );
  SDFFRXL fft_d6_reg_14_ ( .D(N775), .SI(fft_d6[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d6[14]) );
  SDFFRXL fft_d6_reg_13_ ( .D(N774), .SI(fft_d6[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d6[13]) );
  SDFFRXL fft_d6_reg_12_ ( .D(N773), .SI(fft_d6[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d6[12]) );
  SDFFRXL fft_d6_reg_11_ ( .D(N772), .SI(fft_d6[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d6[11]) );
  SDFFRXL fft_d6_reg_10_ ( .D(N771), .SI(fft_d6[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d6[10]) );
  SDFFRXL fft_d6_reg_9_ ( .D(N770), .SI(fft_d6[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d6[9]) );
  SDFFRXL fft_d6_reg_8_ ( .D(N769), .SI(fft_d6[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d6[8]) );
  SDFFRXL fft_d6_reg_7_ ( .D(N768), .SI(fft_d6[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d6[7]) );
  SDFFRXL fft_d6_reg_6_ ( .D(N767), .SI(fft_d6[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d6[6]) );
  SDFFRXL fft_d6_reg_5_ ( .D(N766), .SI(fft_d6[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d6[5]) );
  SDFFRXL fft_d6_reg_4_ ( .D(N765), .SI(fft_d6[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d6[4]) );
  SDFFRXL fft_d6_reg_3_ ( .D(N764), .SI(fft_d6[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d6[3]) );
  SDFFRXL fft_d6_reg_2_ ( .D(N763), .SI(fft_d6[1]), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(fft_d6[2]) );
  SDFFRXL fft_d6_reg_1_ ( .D(N762), .SI(fft_d6[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d6[1]) );
  SDFFRXL fft_d6_reg_0_ ( .D(N761), .SI(n10770), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d6[0]) );
  SDFFRXL fft_d7_reg_31_ ( .D(N824), .SI(fft_d7[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d7[31]) );
  SDFFRXL fft_d7_reg_30_ ( .D(N823), .SI(fft_d7[29]), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(fft_d7[30]) );
  SDFFRXL fft_d7_reg_29_ ( .D(N822), .SI(fft_d7[28]), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(fft_d7[29]) );
  SDFFRXL fft_d7_reg_28_ ( .D(N821), .SI(fft_d7[27]), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(fft_d7[28]) );
  SDFFRXL fft_d7_reg_27_ ( .D(N820), .SI(fft_d7[26]), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(fft_d7[27]) );
  SDFFRXL fft_d7_reg_26_ ( .D(N819), .SI(fft_d7[25]), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(fft_d7[26]) );
  SDFFRXL fft_d7_reg_25_ ( .D(N818), .SI(fft_d7[24]), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(fft_d7[25]) );
  SDFFRXL fft_d7_reg_24_ ( .D(N817), .SI(fft_d7[23]), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(fft_d7[24]) );
  SDFFRXL fft_d7_reg_23_ ( .D(N816), .SI(fft_d7[22]), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(fft_d7[23]) );
  SDFFRXL fft_d7_reg_22_ ( .D(N815), .SI(fft_d7[21]), .SE(test_se), .CK(clk), 
        .RN(n8938), .Q(fft_d7[22]) );
  SDFFRXL fft_d7_reg_21_ ( .D(N814), .SI(fft_d7[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d7[21]) );
  SDFFRXL fft_d7_reg_20_ ( .D(N813), .SI(fft_d7[19]), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(fft_d7[20]) );
  SDFFRXL fft_d7_reg_19_ ( .D(N812), .SI(fft_d7[18]), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(fft_d7[19]) );
  SDFFRXL fft_d7_reg_18_ ( .D(N811), .SI(fft_d7[17]), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(fft_d7[18]) );
  SDFFRXL fft_d7_reg_17_ ( .D(N810), .SI(fft_d7[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d7[17]) );
  SDFFRXL fft_d7_reg_16_ ( .D(N809), .SI(fft_d7[15]), .SE(test_se), .CK(clk), 
        .RN(n9017), .Q(fft_d7[16]) );
  SDFFRXL fft_d7_reg_15_ ( .D(N808), .SI(fft_d7[14]), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(fft_d7[15]) );
  SDFFRXL fft_d7_reg_14_ ( .D(N807), .SI(fft_d7[13]), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(fft_d7[14]) );
  SDFFRXL fft_d7_reg_13_ ( .D(N806), .SI(fft_d7[12]), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(fft_d7[13]) );
  SDFFRXL fft_d7_reg_12_ ( .D(N805), .SI(fft_d7[11]), .SE(test_se), .CK(clk), 
        .RN(n8965), .Q(fft_d7[12]) );
  SDFFRXL fft_d7_reg_11_ ( .D(N804), .SI(fft_d7[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d7[11]) );
  SDFFRXL fft_d7_reg_10_ ( .D(N803), .SI(fft_d7[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d7[10]) );
  SDFFRXL fft_d7_reg_9_ ( .D(N802), .SI(fft_d7[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d7[9]) );
  SDFFRXL fft_d7_reg_8_ ( .D(N801), .SI(fft_d7[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d7[8]) );
  SDFFRXL fft_d7_reg_7_ ( .D(N800), .SI(fft_d7[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d7[7]) );
  SDFFRXL fft_d7_reg_6_ ( .D(N799), .SI(fft_d7[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d7[6]) );
  SDFFRXL fft_d7_reg_5_ ( .D(N798), .SI(fft_d7[4]), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(fft_d7[5]) );
  SDFFRXL fft_d7_reg_4_ ( .D(N797), .SI(fft_d7[3]), .SE(test_se), .CK(clk), 
        .RN(n8993), .Q(fft_d7[4]) );
  SDFFRXL fft_d7_reg_3_ ( .D(N796), .SI(fft_d7[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d7[3]) );
  SDFFRXL fft_d7_reg_2_ ( .D(N795), .SI(fft_d7[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d7[2]) );
  SDFFRXL fft_d7_reg_1_ ( .D(N794), .SI(fft_d7[0]), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(fft_d7[1]) );
  SDFFRXL fft_d7_reg_0_ ( .D(N793), .SI(n10738), .SE(test_se), .CK(clk), .RN(
        n9014), .Q(fft_d7[0]) );
  SDFFRXL fft_d8_reg_31_ ( .D(N856), .SI(fft_d8[30]), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(fft_d8[31]) );
  SDFFRXL fft_d8_reg_30_ ( .D(N855), .SI(fft_d8[29]), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(fft_d8[30]) );
  SDFFRXL fft_d8_reg_29_ ( .D(N854), .SI(fft_d8[28]), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(fft_d8[29]) );
  SDFFRXL fft_d8_reg_28_ ( .D(N853), .SI(fft_d8[27]), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(fft_d8[28]) );
  SDFFRXL fft_d8_reg_27_ ( .D(N852), .SI(fft_d8[26]), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(fft_d8[27]) );
  SDFFRXL fft_d8_reg_26_ ( .D(N851), .SI(fft_d8[25]), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(fft_d8[26]) );
  SDFFRXL fft_d8_reg_25_ ( .D(N850), .SI(fft_d8[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d8[25]) );
  SDFFRXL fft_d8_reg_24_ ( .D(N849), .SI(fft_d8[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d8[24]) );
  SDFFRXL fft_d8_reg_23_ ( .D(N848), .SI(fft_d8[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d8[23]) );
  SDFFRXL fft_d8_reg_22_ ( .D(N847), .SI(fft_d8[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d8[22]) );
  SDFFRXL fft_d8_reg_21_ ( .D(N846), .SI(fft_d8[20]), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(fft_d8[21]) );
  SDFFRXL fft_d8_reg_20_ ( .D(N845), .SI(fft_d8[19]), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(fft_d8[20]) );
  SDFFRXL fft_d8_reg_19_ ( .D(N844), .SI(fft_d8[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d8[19]) );
  SDFFRXL fft_d8_reg_18_ ( .D(N843), .SI(fft_d8[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d8[18]) );
  SDFFRXL fft_d8_reg_17_ ( .D(N842), .SI(fft_d8[16]), .SE(test_se), .CK(clk), 
        .RN(n9013), .Q(fft_d8[17]) );
  SDFFRXL fft_d8_reg_16_ ( .D(N841), .SI(fft_d8[15]), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(fft_d8[16]) );
  SDFFRXL fft_d8_reg_15_ ( .D(N840), .SI(fft_d8[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d8[15]) );
  SDFFRXL fft_d8_reg_14_ ( .D(N839), .SI(fft_d8[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d8[14]) );
  SDFFRXL fft_d8_reg_13_ ( .D(N838), .SI(fft_d8[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d8[13]) );
  SDFFRXL fft_d8_reg_12_ ( .D(N837), .SI(fft_d8[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d8[12]) );
  SDFFRXL fft_d8_reg_11_ ( .D(N836), .SI(fft_d8[10]), .SE(test_se), .CK(clk), 
        .RN(n8962), .Q(fft_d8[11]) );
  SDFFRXL fft_d8_reg_10_ ( .D(N835), .SI(fft_d8[9]), .SE(test_se), .CK(clk), 
        .RN(n8957), .Q(fft_d8[10]) );
  SDFFRXL fft_d8_reg_9_ ( .D(N834), .SI(fft_d8[8]), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(fft_d8[9]) );
  SDFFRXL fft_d8_reg_8_ ( .D(N833), .SI(fft_d8[7]), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(fft_d8[8]) );
  SDFFRXL fft_d8_reg_7_ ( .D(N832), .SI(fft_d8[6]), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(fft_d8[7]) );
  SDFFRXL fft_d8_reg_6_ ( .D(N831), .SI(fft_d8[5]), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(fft_d8[6]) );
  SDFFRXL fft_d8_reg_5_ ( .D(N830), .SI(fft_d8[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d8[5]) );
  SDFFRXL fft_d8_reg_4_ ( .D(N829), .SI(fft_d8[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d8[4]) );
  SDFFRXL fft_d8_reg_3_ ( .D(N828), .SI(fft_d8[2]), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(fft_d8[3]) );
  SDFFRXL fft_d8_reg_2_ ( .D(N827), .SI(fft_d8[1]), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(fft_d8[2]) );
  SDFFRXL fft_d8_reg_1_ ( .D(N826), .SI(fft_d8[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d8[1]) );
  SDFFRXL fft_d8_reg_0_ ( .D(N825), .SI(n10706), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d8[0]) );
  SDFFRXL fft_d9_reg_31_ ( .D(N888), .SI(fft_d9[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d9[31]) );
  SDFFRXL fft_d9_reg_30_ ( .D(N887), .SI(fft_d9[29]), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(fft_d9[30]) );
  SDFFRXL fft_d9_reg_29_ ( .D(N886), .SI(fft_d9[28]), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(fft_d9[29]) );
  SDFFRXL fft_d9_reg_28_ ( .D(N885), .SI(fft_d9[27]), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(fft_d9[28]) );
  SDFFRXL fft_d9_reg_27_ ( .D(N884), .SI(fft_d9[26]), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(fft_d9[27]) );
  SDFFRXL fft_d9_reg_26_ ( .D(N883), .SI(fft_d9[25]), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(fft_d9[26]) );
  SDFFRXL fft_d9_reg_25_ ( .D(N882), .SI(fft_d9[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d9[25]) );
  SDFFRXL fft_d9_reg_24_ ( .D(N881), .SI(fft_d9[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d9[24]) );
  SDFFRXL fft_d9_reg_23_ ( .D(N880), .SI(fft_d9[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d9[23]) );
  SDFFRXL fft_d9_reg_22_ ( .D(N879), .SI(fft_d9[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d9[22]) );
  SDFFRXL fft_d9_reg_21_ ( .D(N878), .SI(fft_d9[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d9[21]) );
  SDFFRXL fft_d9_reg_20_ ( .D(N877), .SI(fft_d9[19]), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(fft_d9[20]) );
  SDFFRXL fft_d9_reg_19_ ( .D(N876), .SI(fft_d9[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d9[19]) );
  SDFFRXL fft_d9_reg_18_ ( .D(N875), .SI(fft_d9[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d9[18]) );
  SDFFRXL fft_d9_reg_17_ ( .D(N874), .SI(fft_d9[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d9[17]) );
  SDFFRXL fft_d9_reg_16_ ( .D(N873), .SI(fft_d9[15]), .SE(test_se), .CK(clk), 
        .RN(n9017), .Q(fft_d9[16]) );
  SDFFRXL fft_d9_reg_15_ ( .D(N872), .SI(fft_d9[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d9[15]) );
  SDFFRXL fft_d9_reg_14_ ( .D(N871), .SI(fft_d9[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d9[14]) );
  SDFFRXL fft_d9_reg_13_ ( .D(N870), .SI(fft_d9[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d9[13]) );
  SDFFRXL fft_d9_reg_12_ ( .D(N869), .SI(fft_d9[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d9[12]) );
  SDFFRXL fft_d9_reg_11_ ( .D(N868), .SI(fft_d9[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d9[11]) );
  SDFFRXL fft_d9_reg_10_ ( .D(N867), .SI(fft_d9[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d9[10]) );
  SDFFRXL fft_d9_reg_9_ ( .D(N866), .SI(fft_d9[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d9[9]) );
  SDFFRXL fft_d9_reg_8_ ( .D(N865), .SI(fft_d9[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d9[8]) );
  SDFFRXL fft_d9_reg_7_ ( .D(N864), .SI(fft_d9[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d9[7]) );
  SDFFRXL fft_d9_reg_6_ ( .D(N863), .SI(fft_d9[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d9[6]) );
  SDFFRXL fft_d9_reg_5_ ( .D(N862), .SI(fft_d9[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d9[5]) );
  SDFFRXL fft_d9_reg_4_ ( .D(N861), .SI(fft_d9[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d9[4]) );
  SDFFRXL fft_d9_reg_3_ ( .D(N860), .SI(fft_d9[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d9[3]) );
  SDFFRXL fft_d9_reg_2_ ( .D(N859), .SI(fft_d9[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d9[2]) );
  SDFFRXL fft_d9_reg_1_ ( .D(N858), .SI(fft_d9[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d9[1]) );
  SDFFRXL fft_d9_reg_0_ ( .D(N857), .SI(n10674), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d9[0]) );
  SDFFRXL fft_d10_reg_31_ ( .D(N920), .SI(fft_d10[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d10[31]) );
  SDFFRXL fft_d10_reg_30_ ( .D(N919), .SI(fft_d10[29]), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(fft_d10[30]) );
  SDFFRXL fft_d10_reg_29_ ( .D(N918), .SI(fft_d10[28]), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(fft_d10[29]) );
  SDFFRXL fft_d10_reg_28_ ( .D(N917), .SI(fft_d10[27]), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(fft_d10[28]) );
  SDFFRXL fft_d10_reg_27_ ( .D(N916), .SI(fft_d10[26]), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(fft_d10[27]) );
  SDFFRXL fft_d10_reg_26_ ( .D(N915), .SI(fft_d10[25]), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(fft_d10[26]) );
  SDFFRXL fft_d10_reg_25_ ( .D(N914), .SI(fft_d10[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d10[25]) );
  SDFFRXL fft_d10_reg_24_ ( .D(N913), .SI(fft_d10[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d10[24]) );
  SDFFRXL fft_d10_reg_23_ ( .D(N912), .SI(fft_d10[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d10[23]) );
  SDFFRXL fft_d10_reg_22_ ( .D(N911), .SI(fft_d10[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d10[22]) );
  SDFFRXL fft_d10_reg_21_ ( .D(N910), .SI(fft_d10[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d10[21]) );
  SDFFRXL fft_d10_reg_20_ ( .D(N909), .SI(fft_d10[19]), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(fft_d10[20]) );
  SDFFRXL fft_d10_reg_19_ ( .D(N908), .SI(fft_d10[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d10[19]) );
  SDFFRXL fft_d10_reg_18_ ( .D(N907), .SI(fft_d10[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d10[18]) );
  SDFFRXL fft_d10_reg_17_ ( .D(N906), .SI(fft_d10[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d10[17]) );
  SDFFRXL fft_d10_reg_16_ ( .D(N905), .SI(fft_d10[15]), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(fft_d10[16]) );
  SDFFRXL fft_d10_reg_15_ ( .D(N904), .SI(fft_d10[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d10[15]) );
  SDFFRXL fft_d10_reg_14_ ( .D(N903), .SI(fft_d10[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d10[14]) );
  SDFFRXL fft_d10_reg_13_ ( .D(N902), .SI(fft_d10[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d10[13]) );
  SDFFRXL fft_d10_reg_12_ ( .D(N901), .SI(fft_d10[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d10[12]) );
  SDFFRXL fft_d10_reg_11_ ( .D(N900), .SI(fft_d10[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d10[11]) );
  SDFFRXL fft_d10_reg_10_ ( .D(N899), .SI(fft_d10[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d10[10]) );
  SDFFRXL fft_d10_reg_9_ ( .D(N898), .SI(fft_d10[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d10[9]) );
  SDFFRXL fft_d10_reg_8_ ( .D(N897), .SI(fft_d10[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d10[8]) );
  SDFFRXL fft_d10_reg_7_ ( .D(N896), .SI(fft_d10[6]), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(fft_d10[7]) );
  SDFFRXL fft_d10_reg_6_ ( .D(N895), .SI(fft_d10[5]), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(fft_d10[6]) );
  SDFFRXL fft_d10_reg_5_ ( .D(N894), .SI(fft_d10[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d10[5]) );
  SDFFRXL fft_d10_reg_4_ ( .D(N893), .SI(fft_d10[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d10[4]) );
  SDFFRXL fft_d10_reg_3_ ( .D(N892), .SI(fft_d10[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d10[3]) );
  SDFFRXL fft_d10_reg_2_ ( .D(N891), .SI(fft_d10[1]), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(fft_d10[2]) );
  SDFFRXL fft_d10_reg_1_ ( .D(N890), .SI(fft_d10[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d10[1]) );
  SDFFRXL fft_d10_reg_0_ ( .D(N889), .SI(n10642), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d10[0]) );
  SDFFRXL fft_d11_reg_31_ ( .D(N952), .SI(fft_d11[30]), .SE(test_se), .CK(clk), 
        .RN(n8983), .Q(fft_d11[31]) );
  SDFFRXL fft_d11_reg_30_ ( .D(N951), .SI(fft_d11[29]), .SE(test_se), .CK(clk), 
        .RN(n8978), .Q(fft_d11[30]) );
  SDFFRXL fft_d11_reg_29_ ( .D(N950), .SI(fft_d11[28]), .SE(test_se), .CK(clk), 
        .RN(n8973), .Q(fft_d11[29]) );
  SDFFRXL fft_d11_reg_28_ ( .D(N949), .SI(fft_d11[27]), .SE(test_se), .CK(clk), 
        .RN(n8968), .Q(fft_d11[28]) );
  SDFFRXL fft_d11_reg_27_ ( .D(N948), .SI(fft_d11[26]), .SE(test_se), .CK(clk), 
        .RN(n8963), .Q(fft_d11[27]) );
  SDFFRXL fft_d11_reg_26_ ( .D(N947), .SI(fft_d11[25]), .SE(test_se), .CK(clk), 
        .RN(n8958), .Q(fft_d11[26]) );
  SDFFRXL fft_d11_reg_25_ ( .D(N946), .SI(fft_d11[24]), .SE(test_se), .CK(clk), 
        .RN(n8953), .Q(fft_d11[25]) );
  SDFFRXL fft_d11_reg_24_ ( .D(N945), .SI(fft_d11[23]), .SE(test_se), .CK(clk), 
        .RN(n8948), .Q(fft_d11[24]) );
  SDFFRXL fft_d11_reg_23_ ( .D(N944), .SI(fft_d11[22]), .SE(test_se), .CK(clk), 
        .RN(n8943), .Q(fft_d11[23]) );
  SDFFRXL fft_d11_reg_22_ ( .D(N943), .SI(fft_d11[21]), .SE(test_se), .CK(clk), 
        .RN(n8938), .Q(fft_d11[22]) );
  SDFFRXL fft_d11_reg_21_ ( .D(N942), .SI(fft_d11[20]), .SE(test_se), .CK(clk), 
        .RN(n8991), .Q(fft_d11[21]) );
  SDFFRXL fft_d11_reg_20_ ( .D(N941), .SI(fft_d11[19]), .SE(test_se), .CK(clk), 
        .RN(n8996), .Q(fft_d11[20]) );
  SDFFRXL fft_d11_reg_19_ ( .D(N940), .SI(fft_d11[18]), .SE(test_se), .CK(clk), 
        .RN(n9001), .Q(fft_d11[19]) );
  SDFFRXL fft_d11_reg_18_ ( .D(N939), .SI(fft_d11[17]), .SE(test_se), .CK(clk), 
        .RN(n9006), .Q(fft_d11[18]) );
  SDFFRXL fft_d11_reg_17_ ( .D(N938), .SI(fft_d11[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d11[17]) );
  SDFFRXL fft_d11_reg_16_ ( .D(N937), .SI(fft_d11[15]), .SE(test_se), .CK(clk), 
        .RN(n9017), .Q(fft_d11[16]) );
  SDFFRXL fft_d11_reg_15_ ( .D(N936), .SI(fft_d11[14]), .SE(test_se), .CK(clk), 
        .RN(n8980), .Q(fft_d11[15]) );
  SDFFRXL fft_d11_reg_14_ ( .D(N935), .SI(fft_d11[13]), .SE(test_se), .CK(clk), 
        .RN(n8975), .Q(fft_d11[14]) );
  SDFFRXL fft_d11_reg_13_ ( .D(N934), .SI(fft_d11[12]), .SE(test_se), .CK(clk), 
        .RN(n8970), .Q(fft_d11[13]) );
  SDFFRXL fft_d11_reg_12_ ( .D(N933), .SI(fft_d11[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d11[12]) );
  SDFFRXL fft_d11_reg_11_ ( .D(N932), .SI(fft_d11[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d11[11]) );
  SDFFRXL fft_d11_reg_10_ ( .D(N931), .SI(fft_d11[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d11[10]) );
  SDFFRXL fft_d11_reg_9_ ( .D(N930), .SI(fft_d11[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d11[9]) );
  SDFFRXL fft_d11_reg_8_ ( .D(N929), .SI(fft_d11[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d11[8]) );
  SDFFRXL fft_d11_reg_7_ ( .D(N928), .SI(fft_d11[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d11[7]) );
  SDFFRXL fft_d11_reg_6_ ( .D(N927), .SI(fft_d11[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d11[6]) );
  SDFFRXL fft_d11_reg_5_ ( .D(N926), .SI(fft_d11[4]), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(fft_d11[5]) );
  SDFFRXL fft_d11_reg_4_ ( .D(N925), .SI(fft_d11[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d11[4]) );
  SDFFRXL fft_d11_reg_3_ ( .D(N924), .SI(fft_d11[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d11[3]) );
  SDFFRXL fft_d11_reg_2_ ( .D(N923), .SI(fft_d11[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d11[2]) );
  SDFFRXL fft_d11_reg_1_ ( .D(N922), .SI(fft_d11[0]), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(fft_d11[1]) );
  SDFFRXL fft_d11_reg_0_ ( .D(N921), .SI(n10610), .SE(test_se), .CK(clk), .RN(
        n9014), .Q(fft_d11[0]) );
  SDFFRXL fft_d12_reg_31_ ( .D(N984), .SI(fft_d12[30]), .SE(test_se), .CK(clk), 
        .RN(n8984), .Q(fft_d12[31]) );
  SDFFRXL fft_d12_reg_30_ ( .D(N983), .SI(fft_d12[29]), .SE(test_se), .CK(clk), 
        .RN(n8979), .Q(fft_d12[30]) );
  SDFFRXL fft_d12_reg_29_ ( .D(N982), .SI(fft_d12[28]), .SE(test_se), .CK(clk), 
        .RN(n8974), .Q(fft_d12[29]) );
  SDFFRXL fft_d12_reg_28_ ( .D(N981), .SI(fft_d12[27]), .SE(test_se), .CK(clk), 
        .RN(n8969), .Q(fft_d12[28]) );
  SDFFRXL fft_d12_reg_27_ ( .D(N980), .SI(fft_d12[26]), .SE(test_se), .CK(clk), 
        .RN(n8964), .Q(fft_d12[27]) );
  SDFFRXL fft_d12_reg_26_ ( .D(N979), .SI(fft_d12[25]), .SE(test_se), .CK(clk), 
        .RN(n8959), .Q(fft_d12[26]) );
  SDFFRXL fft_d12_reg_25_ ( .D(N978), .SI(fft_d12[24]), .SE(test_se), .CK(clk), 
        .RN(n8954), .Q(fft_d12[25]) );
  SDFFRXL fft_d12_reg_24_ ( .D(N977), .SI(fft_d12[23]), .SE(test_se), .CK(clk), 
        .RN(n8949), .Q(fft_d12[24]) );
  SDFFRXL fft_d12_reg_23_ ( .D(N976), .SI(fft_d12[22]), .SE(test_se), .CK(clk), 
        .RN(n8944), .Q(fft_d12[23]) );
  SDFFRXL fft_d12_reg_22_ ( .D(N975), .SI(fft_d12[21]), .SE(test_se), .CK(clk), 
        .RN(n8939), .Q(fft_d12[22]) );
  SDFFRXL fft_d12_reg_21_ ( .D(N974), .SI(fft_d12[20]), .SE(test_se), .CK(clk), 
        .RN(n8992), .Q(fft_d12[21]) );
  SDFFRXL fft_d12_reg_20_ ( .D(N973), .SI(fft_d12[19]), .SE(test_se), .CK(clk), 
        .RN(n8997), .Q(fft_d12[20]) );
  SDFFRXL fft_d12_reg_19_ ( .D(N972), .SI(fft_d12[18]), .SE(test_se), .CK(clk), 
        .RN(n9002), .Q(fft_d12[19]) );
  SDFFRXL fft_d12_reg_18_ ( .D(N971), .SI(fft_d12[17]), .SE(test_se), .CK(clk), 
        .RN(n9007), .Q(fft_d12[18]) );
  SDFFRXL fft_d12_reg_17_ ( .D(N970), .SI(fft_d12[16]), .SE(test_se), .CK(clk), 
        .RN(n9012), .Q(fft_d12[17]) );
  SDFFRXL fft_d12_reg_16_ ( .D(N969), .SI(fft_d12[15]), .SE(test_se), .CK(clk), 
        .RN(n9018), .Q(fft_d12[16]) );
  SDFFRXL fft_d12_reg_15_ ( .D(N968), .SI(fft_d12[14]), .SE(test_se), .CK(clk), 
        .RN(n8981), .Q(fft_d12[15]) );
  SDFFRXL fft_d12_reg_14_ ( .D(N967), .SI(fft_d12[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d12[14]) );
  SDFFRXL fft_d12_reg_13_ ( .D(N966), .SI(fft_d12[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d12[13]) );
  SDFFRXL fft_d12_reg_12_ ( .D(N965), .SI(fft_d12[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d12[12]) );
  SDFFRXL fft_d12_reg_11_ ( .D(N964), .SI(fft_d12[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d12[11]) );
  SDFFRXL fft_d12_reg_10_ ( .D(N963), .SI(fft_d12[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d12[10]) );
  SDFFRXL fft_d12_reg_9_ ( .D(N962), .SI(fft_d12[8]), .SE(test_se), .CK(clk), 
        .RN(n8952), .Q(fft_d12[9]) );
  SDFFRXL fft_d12_reg_8_ ( .D(N961), .SI(fft_d12[7]), .SE(test_se), .CK(clk), 
        .RN(n8947), .Q(fft_d12[8]) );
  SDFFRXL fft_d12_reg_7_ ( .D(N960), .SI(fft_d12[6]), .SE(test_se), .CK(clk), 
        .RN(n8942), .Q(fft_d12[7]) );
  SDFFRXL fft_d12_reg_6_ ( .D(N959), .SI(fft_d12[5]), .SE(test_se), .CK(clk), 
        .RN(n8934), .Q(fft_d12[6]) );
  SDFFRXL fft_d12_reg_5_ ( .D(N958), .SI(fft_d12[4]), .SE(test_se), .CK(clk), 
        .RN(n8989), .Q(fft_d12[5]) );
  SDFFRXL fft_d12_reg_4_ ( .D(N957), .SI(fft_d12[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d12[4]) );
  SDFFRXL fft_d12_reg_3_ ( .D(N956), .SI(fft_d12[2]), .SE(test_se), .CK(clk), 
        .RN(n9000), .Q(fft_d12[3]) );
  SDFFRXL fft_d12_reg_2_ ( .D(N955), .SI(fft_d12[1]), .SE(test_se), .CK(clk), 
        .RN(n9005), .Q(fft_d12[2]) );
  SDFFRXL fft_d12_reg_1_ ( .D(N954), .SI(fft_d12[0]), .SE(test_se), .CK(clk), 
        .RN(n9010), .Q(fft_d12[1]) );
  SDFFRXL fft_d12_reg_0_ ( .D(N953), .SI(n10578), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d12[0]) );
  SDFFRXL fft_d13_reg_31_ ( .D(N1016), .SI(fft_d13[30]), .SE(test_se), .CK(clk), .RN(n8983), .Q(fft_d13[31]) );
  SDFFRXL fft_d13_reg_30_ ( .D(N1015), .SI(fft_d13[29]), .SE(test_se), .CK(clk), .RN(n8978), .Q(fft_d13[30]) );
  SDFFRXL fft_d13_reg_29_ ( .D(N1014), .SI(fft_d13[28]), .SE(test_se), .CK(clk), .RN(n8973), .Q(fft_d13[29]) );
  SDFFRXL fft_d13_reg_28_ ( .D(N1013), .SI(fft_d13[27]), .SE(test_se), .CK(clk), .RN(n8968), .Q(fft_d13[28]) );
  SDFFRXL fft_d13_reg_27_ ( .D(N1012), .SI(fft_d13[26]), .SE(test_se), .CK(clk), .RN(n8963), .Q(fft_d13[27]) );
  SDFFRXL fft_d13_reg_26_ ( .D(N1011), .SI(fft_d13[25]), .SE(test_se), .CK(clk), .RN(n8958), .Q(fft_d13[26]) );
  SDFFRXL fft_d13_reg_25_ ( .D(N1010), .SI(fft_d13[24]), .SE(test_se), .CK(clk), .RN(n8953), .Q(fft_d13[25]) );
  SDFFRXL fft_d13_reg_24_ ( .D(N1009), .SI(fft_d13[23]), .SE(test_se), .CK(clk), .RN(n8948), .Q(fft_d13[24]) );
  SDFFRXL fft_d13_reg_23_ ( .D(N1008), .SI(fft_d13[22]), .SE(test_se), .CK(clk), .RN(n8944), .Q(fft_d13[23]) );
  SDFFRXL fft_d13_reg_22_ ( .D(N1007), .SI(fft_d13[21]), .SE(test_se), .CK(clk), .RN(n8939), .Q(fft_d13[22]) );
  SDFFRXL fft_d13_reg_21_ ( .D(N1006), .SI(fft_d13[20]), .SE(test_se), .CK(clk), .RN(n8991), .Q(fft_d13[21]) );
  SDFFRXL fft_d13_reg_20_ ( .D(N1005), .SI(fft_d13[19]), .SE(test_se), .CK(clk), .RN(n8996), .Q(fft_d13[20]) );
  SDFFRXL fft_d13_reg_19_ ( .D(N1004), .SI(fft_d13[18]), .SE(test_se), .CK(clk), .RN(n9001), .Q(fft_d13[19]) );
  SDFFRXL fft_d13_reg_18_ ( .D(N1003), .SI(fft_d13[17]), .SE(test_se), .CK(clk), .RN(n9007), .Q(fft_d13[18]) );
  SDFFRXL fft_d13_reg_17_ ( .D(N1002), .SI(fft_d13[16]), .SE(test_se), .CK(clk), .RN(n9012), .Q(fft_d13[17]) );
  SDFFRXL fft_d13_reg_16_ ( .D(N1001), .SI(fft_d13[15]), .SE(test_se), .CK(clk), .RN(n9017), .Q(fft_d13[16]) );
  SDFFRXL fft_d13_reg_15_ ( .D(N1000), .SI(fft_d13[14]), .SE(test_se), .CK(clk), .RN(n8980), .Q(fft_d13[15]) );
  SDFFRXL fft_d13_reg_14_ ( .D(N999), .SI(fft_d13[13]), .SE(test_se), .CK(clk), 
        .RN(n8976), .Q(fft_d13[14]) );
  SDFFRXL fft_d13_reg_13_ ( .D(N998), .SI(fft_d13[12]), .SE(test_se), .CK(clk), 
        .RN(n8971), .Q(fft_d13[13]) );
  SDFFRXL fft_d13_reg_12_ ( .D(N997), .SI(fft_d13[11]), .SE(test_se), .CK(clk), 
        .RN(n8966), .Q(fft_d13[12]) );
  SDFFRXL fft_d13_reg_11_ ( .D(N996), .SI(fft_d13[10]), .SE(test_se), .CK(clk), 
        .RN(n8961), .Q(fft_d13[11]) );
  SDFFRXL fft_d13_reg_10_ ( .D(N995), .SI(fft_d13[9]), .SE(test_se), .CK(clk), 
        .RN(n8956), .Q(fft_d13[10]) );
  SDFFRXL fft_d13_reg_9_ ( .D(N994), .SI(fft_d13[8]), .SE(test_se), .CK(clk), 
        .RN(n8951), .Q(fft_d13[9]) );
  SDFFRXL fft_d13_reg_8_ ( .D(N993), .SI(fft_d13[7]), .SE(test_se), .CK(clk), 
        .RN(n8946), .Q(fft_d13[8]) );
  SDFFRXL fft_d13_reg_7_ ( .D(N992), .SI(fft_d13[6]), .SE(test_se), .CK(clk), 
        .RN(n8941), .Q(fft_d13[7]) );
  SDFFRXL fft_d13_reg_6_ ( .D(N991), .SI(fft_d13[5]), .SE(test_se), .CK(clk), 
        .RN(n8933), .Q(fft_d13[6]) );
  SDFFRXL fft_d13_reg_5_ ( .D(N990), .SI(fft_d13[4]), .SE(test_se), .CK(clk), 
        .RN(n8988), .Q(fft_d13[5]) );
  SDFFRXL fft_d13_reg_4_ ( .D(N989), .SI(fft_d13[3]), .SE(test_se), .CK(clk), 
        .RN(n8994), .Q(fft_d13[4]) );
  SDFFRXL fft_d13_reg_3_ ( .D(N988), .SI(fft_d13[2]), .SE(test_se), .CK(clk), 
        .RN(n8999), .Q(fft_d13[3]) );
  SDFFRXL fft_d13_reg_2_ ( .D(N987), .SI(fft_d13[1]), .SE(test_se), .CK(clk), 
        .RN(n9004), .Q(fft_d13[2]) );
  SDFFRXL fft_d13_reg_1_ ( .D(N986), .SI(fft_d13[0]), .SE(test_se), .CK(clk), 
        .RN(n9009), .Q(fft_d13[1]) );
  SDFFRXL fft_d13_reg_0_ ( .D(N985), .SI(n10546), .SE(test_se), .CK(clk), .RN(
        n9015), .Q(fft_d13[0]) );
  SDFFRXL done_reg ( .D(n6071), .SI(n11219), .SE(test_se), .CK(clk), .RN(n9127), .Q(done) );
  SDFFRXL freq_reg_3_ ( .D(N1233), .SI(freq[2]), .SE(test_se), .CK(clk), .RN(
        n8938), .Q(freq[3]) );
  SDFFRXL freq_reg_2_ ( .D(N1232), .SI(freq[1]), .SE(test_se), .CK(clk), .RN(
        n8938), .Q(freq[2]) );
  SDFFRXL freq_reg_1_ ( .D(N1231), .SI(freq[0]), .SE(test_se), .CK(clk), .RN(
        n8938), .Q(freq[1]) );
  SDFFRXL freq_reg_0_ ( .D(N1230), .SI(n11210), .SE(test_se), .CK(clk), .RN(
        n8938), .Q(freq[0]) );
  INVXL U8024 ( .A(n6078), .Y(n11211) );
  INVXL U8025 ( .A(n11211), .Y(n11212) );
  INVXL U8026 ( .A(n11211), .Y(n11213) );
  INVXL U8027 ( .A(n11223), .Y(n11214) );
  INVXL U8028 ( .A(n11214), .Y(n11215) );
  INVXL U8029 ( .A(n11214), .Y(n11216) );
  INVXL U8030 ( .A(d32[31]), .Y(n11217) );
  INVXL U8031 ( .A(n11217), .Y(n11218) );
  INVXL U8032 ( .A(n11217), .Y(n11219) );
  INVXL U8033 ( .A(n10471), .Y(n11220) );
  INVXL U8034 ( .A(n11220), .Y(n11221) );
  INVXL U8035 ( .A(n11220), .Y(n11222) );
  INVXL U8036 ( .A(n11220), .Y(n11223) );
  INVXL U8037 ( .A(n11220), .Y(n11224) );
endmodule

